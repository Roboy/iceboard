// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Sep  8 12:22:14 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, n624, 
        GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    
    wire n50736;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n26, n5;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n731, data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(352[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(360[15:20])
    
    wire pwm_setpoint_23__N_207, n62676, n12146, n12150, n37154, n10, 
        n260, n12186, n294, n298, n299, n300, n301, n302, n303, 
        n304, n305, n306, n307, n308, n309, n4930, n4929, n4928, 
        n4927, n4926, n4925, n4924, n4923, n4922, n4921, n4920, 
        n4919, n8, n7;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n42168;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    
    wire n29895;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n25568, GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, 
        GLC_N_400, dti_N_404, n29891, n29888, RX_N_2, n67210, n67204, 
        n67200, n67196, n69766, n1744, n1742;
    wire [31:0]motor_state_23__N_91;
    wire [32:0]encoder0_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        read_N_409, n62670, n1319, n68692, n68682, n68681, n15, 
        n13, n12, n11, n10_adj_5699, n9, n8_adj_5700, n4, n26_adj_5701, 
        n19, n17, n16, n15_adj_5702, n13_adj_5703, n1784, n1786, 
        n1788, n1790, n1792, n1794, n1796;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n1822, n1824;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [1:0]state;   // verilog/neopixel.v(16[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    
    wire n62664;
    wire [5:0]color_bit_N_502;
    
    wire n8_adj_5704, n4918, n4917, n4916, n4915, n4914, n4913, 
        n4912, n29885, n551, n62660, n29881, n4942, n4939, n70345, 
        n29878, n29875, n11_adj_5705, n9_adj_5706, n8_adj_5707, n7_adj_5708, 
        n6, n5_adj_5709, n4_adj_5710, n29872, n50735, n25573, n2, 
        n625, n623, n622, n621, n14, n15_adj_5711, n16_adj_5712, 
        n17_adj_5713, n18, n19_adj_5714, n20, n21, n22, n23, n24, 
        n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire n50734, n29869, n42981;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n19_adj_5715, n25_adj_5716, 
        n24_adj_5717, n17_adj_5718, n23_adj_5719, n22_adj_5720, n21_adj_5721, 
        n20_adj_5722, n2821, n50316, n29866, n2874, n22773, n62648, 
        n42331, n62644, n4911, n4910, n4909, n57733, n58988, n50299, 
        n29012, n57863, n57862, n57861, n57860, n57859, n57858, 
        n57864, n57857, n57856, n57855, n57854, n57853, n57852, 
        n28997, n57851, n57850, n57849, n57848, n57847, n57846, 
        n57845, n57844, n28988, n57843, n57842, n57841, n57840, 
        n57839, n57838, n57837, n57836, n57835, n57834, n57833, 
        n57832, n57831, n57830, n57829, n57828, n57827, n57826, 
        n57825, n57824, n57823, n57822, n57821, n57820, n57819, 
        n57735, n57818, n28960, n57817, n57816, n57815, n57814, 
        n57813, n57812, n57811, n57810, n57809, n57808, n57807, 
        n57806, n57805, n57804, n57736, n57737, n57738, n57739, 
        n57740, n28940, n57741, n57742, n57743, n57744, n57745, 
        n57746, n57747, n28932, n57748, n57749, n57750, n57751, 
        n57752, n57753, n57754, n28924, n57755, n57756, n57757, 
        n57758, n57759, n57760, n28917, n57761, n57762, n57763, 
        n28911, n28910, n57764, n57765, n57766, n57767, n57768, 
        n57769, n57770, n57771, n57772, n57773, n57774, n57775, 
        n57776, n57777, n57778, n57779, n28893, n57780, n57781, 
        n57782, n57783, n57784, n57785, n57786, n57787, n57788, 
        n57789, n57790, n57791, n57792, n57793, n57794, n57795, 
        n57796, n57797, n57798, n57799, n57800, n57801, n57802, 
        n57803, n57927, n62638, n28822, n23_adj_5723, n62636, n29863, 
        n62630, n25_adj_5724, n61029, n62628, n62620, n50986, n67956, 
        n50985, n62610, n68549, n62604, n69501, n50984, n50983, 
        n50982, n50981, n50980, n50979, n50978, n50977, n50976, 
        n50975, n68253, n50974, n62598, n50973, n50972, n14_adj_5725, 
        n50971, n10_adj_5726, n50715, n50714, n58929, n2076, n62592, 
        n62590, n62588, n58897, n62582, n67890, n61098, n70339, 
        n70333, n50713, n67976, n62568, n20_adj_5727, n50712, n66110, 
        n29860, n67884, n69078, n69279, n67151, n62562, n62556, 
        n62554, n62548, n62542, n50970, n29857, n62540, n50711, 
        n58821, n63902, n63659, n29854, n12184, n50969, n62536, 
        n67846, n62528, Kp_23__N_1301, n62524, n58801, n58799, n25555, 
        n58797, n58795, n62518, n58792, n62514, n69734, n29, n27, 
        n62506, n23_adj_5728, n62500, n10_adj_5729, n62494, n50968, 
        n12148, n50967, n29851, n32, n31, n30, n29_adj_5730, n28, 
        n27_adj_5731, n29848, n26_adj_5732, n25_adj_5733, n24_adj_5734, 
        n23_adj_5735, n22_adj_5736, n21_adj_5737, n20_adj_5738, n19_adj_5739, 
        n18_adj_5740, n62492, n17_adj_5741, n16_adj_5742, n15_adj_5743, 
        n14_adj_5744, n13_adj_5745, n12_adj_5746, \FRAME_MATCHER.i_31__N_2509 , 
        n11_adj_5747, n68618, n30779, n30778, n62486, n50710, n29844, 
        n29841, n29838, n29837, n29836, n29835, n29834, n29833, 
        n29832, n29831, n29830, n29829, n29828, n29827, n29826, 
        n29825, n62484, n29818, n29813, n29729, n29728, n29727, 
        n29726, n29725, n29724, n29723, n29722, n29721, n29720, 
        n29719, n29718, n29717, n29716, n29715, n29714, n29713, 
        n29712, n29709, n29708, n29707, n29706, n29703, n29702, 
        n29701, n29698, n29697, n29677, n29676, n29674, n29673, 
        n29672, n29671, n29669, n29666, n29664, n29657, n29656, 
        n29655, n29654, n50966, n50709, n50708, n10_adj_5748, n50707, 
        n29653, n29652, n29651, n29650, n29646, n29645, n29644, 
        n29641, n29640, n29639, n29637, n29630, n29625, n43043, 
        n29621, n29617, n29615, n29606, n43037, n29603, n43035, 
        n29600, n29596, n29595, n29592, n29591, n29590, n29584, 
        n43029, n29581, n29578, n43025, n29575, n29566, n29560, 
        n29559, n29558, n29557, n43019, n29541, n43013, n29538, 
        n42925, n43007, n43003, n43001, n29520, n42997, n29514, 
        n42995, n29511, n29508, n29505, n29502, n57169, n43039, 
        n43111, n43085, n43081, n29442, n6_adj_5749, n62468, n68619, 
        n67133, n9_adj_5750, n8_adj_5751, n7_adj_5752, n6_adj_5753, 
        n30_adj_5754, n68673, n23_adj_5755, n21_adj_5756, n19_adj_5757, 
        n17_adj_5758, n16_adj_5759, n15_adj_5760, n13_adj_5761, n11_adj_5762, 
        n10_adj_5763, n9_adj_5764, n8_adj_5765, n7_adj_5766, n6_adj_5767, 
        n4_adj_5768, n50706, n50965, n12_adj_5769, n62462, n30719, 
        n30718, n30717, n62456, n9_adj_5770, n62452, n30691, n30689, 
        n62448, n30687, n30686, n30680, n4_adj_5771, n4_adj_5772, 
        n62438, n67687, n62434, n11_adj_5773, n62428, n30568, n30561, 
        n30552, n70441, n6_adj_5774, n58046, n30452, n30445, n30441, 
        n30440, n5_adj_5775, n30436, n30429, n67123, n30425, n50705, 
        n135, n150, n156, n182, n187, n214, n219, n244, n405, 
        n406, n50704, n478, n500, n4_adj_5776;
    wire [23:0]duty_23__N_3602;
    
    wire n6_adj_5777, n3, n2_adj_5778;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3834, position_31__N_3837, n62402, 
        n30390, n8_adj_5779, n30389, n30388, n30387, n30386, n30385, 
        n30374, n30373;
    wire [1:0]a_new_adj_5988;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5989;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5782, b_prev_adj_5783, debounce_cnt_N_3834_adj_5784, 
        n30372, n30371, n30370, n30369, n30368, n30367, n30365, 
        position_31__N_3837_adj_5785, n30364, n62396, n8_adj_5786, n405_adj_5787, 
        n30363, n30362, n30361, n30360, n30359, n50703, n30358, 
        n21_adj_5788, n30357, n30356, n30355, n5_adj_5789;
    wire [7:0]data_adj_6002;   // verilog/eeprom.v(23[12:16])
    wire [7:0]state_7__N_3919;
    
    wire n70327, n70321, n62386, n70435, n8_adj_5790, n62384, n6619, 
        n11_adj_5791, n50702, n37050, n30294, n30293, n30292, n30291, 
        n30289, n4908, n4907, n30288;
    wire [15:0]data_adj_6010;   // verilog/tli4970.v(27[14:18])
    
    wire n25563, n62382, n30287, n30286, n30285, n19_adj_5800, n18_adj_5801, 
        n17_adj_5802, n4_adj_5803, n3_adj_5804, n2_adj_5805, n50315, 
        n62380, n15_adj_5806, n8_adj_5807, n30276, n15_adj_5808, n50701, 
        n6_adj_5809, n61122, n12152, n12154, n12156, n12158, n15_adj_5810, 
        state_7__N_4320, n22760, n16_adj_5811, n5_adj_5812, n62366, 
        r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n68617, n22841, n12160, n12162, n12164, n12166, n12168, 
        n12170, n12172, n12174, n62360;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n12176, n12178, n12180;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n15_adj_5813, n14_adj_5814, n13_adj_5815, n12_adj_5816, n51771, 
        n30187;
    wire [8:0]r_Clock_Count_adj_6024;   // verilog/uart_tx.v(33[16:29])
    
    wire n51770, n51769, n51768;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n11_adj_5825, n10_adj_5826, n9_adj_5827, n8_adj_5828, n7_adj_5829, 
        n6_adj_5830, n30169, n62350, n7_adj_5831;
    wire [7:0]state_adj_6035;   // verilog/i2c_controller.v(33[12:17])
    
    wire enable_slow_N_4214, n5_adj_5833;
    wire [7:0]state_7__N_4111;
    
    wire n51767, n6429, n62346;
    wire [7:0]state_7__N_4127;
    
    wire n30149, n62344, n51766, n62342, n57221, n57223, n51765, 
        n29423, n43071, n57225, n15_adj_5834, n62338, n59639, n29413, 
        n29410, n14_adj_5835, n51764, n62334, n62332, n7449, n7448, 
        n7447, n7446, n7445, n7444, n62330, n62328, n828, n829, 
        n830, n831, n832, n833, n834, n861, n896, n897, n898, 
        n899, n900, n901, n927, n928, n929, n930, n931, n932, 
        n933, n934, n935, n936, n937, n938, n939, n940, n941, 
        n942, n943, n944, n945, n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n960, n36515, 
        n995, n996, n997, n998, n999, n1000, n1001, n1026, n1027, 
        n1028, n1029, n1030, n1031, n1032, n1033, n62320, n1059, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
        n1132, n1133, n1158, n1193, n1194, n1195, n1196, n1197, 
        n1198, n1199, n1200, n1201, n1224_adj_5836, n1225_adj_5837, 
        n1226_adj_5838, n1227_adj_5839, n1228_adj_5840, n1229_adj_5841, 
        n1230_adj_5842, n1231_adj_5843, n1232_adj_5844, n1233_adj_5845, 
        n1257, n62312, n1292, n1293, n1294, n1295, n1296, n1297, 
        n1298, n1299, n1300, n1301, n59677, n1323, n1324, n1325, 
        n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, 
        n1356, n34, n1391, n1392, n1393, n1394, n1395, n1396, 
        n1397, n1398, n1399, n1400, n1401, n62308, n1422, n1423, 
        n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
        n1432, n1433, n1455, n51763, n51762, n51761, n51760, n1490, 
        n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
        n1499, n1500, n1501, n1521, n1522, n1523, n1524, n1525, 
        n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
        n1554, n51759, n1589, n1590, n1591, n1592, n1593, n1594, 
        n1595, n1596, n1597, n1598, n1599, n1600, n1601, n51758, 
        n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
        n1628, n1629, n1630, n1631, n1632, n1633, n62302, n1653, 
        n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
        n1696, n1697, n1698, n1699, n1700, n1701, n1719, n1720, 
        n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
        n1729, n1730, n1731, n1732, n1733, n1752, n51757, n478_adj_5846, 
        n1787, n1788_adj_5847, n1789, n1790_adj_5848, n1791, n1792_adj_5849, 
        n1793, n1794_adj_5850, n1795, n1796_adj_5851, n1797, n1798, 
        n1799, n1800, n1801, n1818, n1819, n1820, n1821, n1822_adj_5852, 
        n1823, n1824_adj_5853, n1825, n1826, n1827, n1828, n1829, 
        n1830, n1831, n1832, n1833, n18_adj_5854, n62294, n1851, 
        n50937, n62288, n1886, n1887, n1888, n1889, n1890, n1891, 
        n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
        n1900, n1901, n51756, n51755, n62286, n51754, n51753, 
        n51752, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
        n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
        n1932, n1933, n50298, n50936, n50935, n70357, n1950, n50934, 
        n51751, n50933, n51750, n51749, n50932, n50931, n51294, 
        n51748, n51747, n51293, n51292, n51746, n51291, n1985, 
        n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
        n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
        n50930, n62280, n2016, n2017, n2018, n2019, n2020, n2021, 
        n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
        n2030, n2031, n2032, n2033, n62278, n7_adj_5855, n2049, 
        n50929, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
        n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
        n2099, n2100, n2101, n2115, n2116, n2117, n2118, n2119, 
        n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
        n2128, n2129, n2130, n2131, n2132, n2133, n2148, n51290, 
        n50928, n50927, n51745, n50926, n50925, n51289, n51288, 
        n51287, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
        n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
        n2198, n2199, n2200, n2201, n50924, n50923, n51744, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n51743, n51742, n62272, n2247, n51286, 
        n51741, n51285, n51284, n2282, n2283, n2284, n2285, n2286, 
        n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
        n2295, n2296, n2297, n2298, n2299, n2300, n2301, n70423, 
        n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
        n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
        n2329, n2330, n2331, n2332, n2333, n2346, n2381, n2382, 
        n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
        n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
        n2399, n2400, n2401, n2412, n2413, n2414, n2415, n2416, 
        n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
        n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
        n2433, n2445, n51283, n2480, n2481, n2482, n2483, n2484, 
        n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
        n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
        n2501, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
        n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, 
        n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
        n2544, n51282, n67527, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
        n2600, n2601, n2610, n2611, n2612, n2613, n2614, n2615, 
        n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2643, n51281, n51280, n62256, n2677, n2678, 
        n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
        n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
        n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2709, 
        n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
        n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
        n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
        n2742, n50922, n67525, n2776, n2777, n2778, n2779, n2780, 
        n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
        n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
        n2797, n2798, n2799, n2800, n2801, n51279, n2808, n2809, 
        n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
        n2818, n2819, n2820, n2821_adj_5856, n2822, n2823, n2824, 
        n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
        n2833, n2841, n51278, n2876, n2877, n2878, n2879, n2880, 
        n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
        n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
        n2897, n2898, n2899, n2900, n2901, n2907, n2908, n2909, 
        n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
        n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
        n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
        n2940, n62250, n51277, n51276, n70042, n405_adj_5857, n2975, 
        n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
        n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
        n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
        n3000, n3001, n3006, n3007, n3008, n3009, n3010, n3011, 
        n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
        n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
        n3028, n3029, n3030, n3031, n3032, n3033, n3039, n3074, 
        n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
        n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, 
        n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
        n3099, n3100, n3101, n3105, n3106, n3107, n3108, n3109, 
        n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
        n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
        n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
        n3138, n67519, n3173, n3174, n3175, n3176, n3177, n3178, 
        n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
        n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
        n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3204, 
        n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
        n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, 
        n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
        n3229, n3230, n3231, n3232, n3233, n69467, n3237, n3271, 
        n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
        n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, 
        n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, 
        n3296, n3298, n3301, n50921, n51275, n58169, n50920, n50919, 
        n51274, n62244, n50918, n50917, n51273, n7_adj_5858, n62236, 
        n67509, n62232, n50688, n24_adj_5859, n51272, n62226, n62224, 
        n62, n51271, n25457, n50687, n51270, n62222, n62220, n50686, 
        n62218, n51269, n51268, n51267, n69704, n62212, n27924, 
        n27922, n62210, n40525, n62204, n62198, n27845, n51266, 
        n43047, n51265, n51264, n60931, n27799, n25532, n50685, 
        n27779, n51263, n61008, n51262, n51261, n51260, n62188, 
        n27735, n62182, n62180, n27722, n70417, n70025, n41, n69461, 
        n70007, n62174, n27704, n62172, n62160, n332, n51259, 
        n51258, n51257, n51256, n51255, n68672, n259, n51254, 
        n50684, n25666, n62154, n51253, n51252, n59761, n8_adj_5860, 
        n27648, n7_adj_5861, n62148, n51251, n70411, n18_adj_5862, 
        n51250, n21_adj_5863, n50683, n61041, n20_adj_5864, n19_adj_5865, 
        n62142, n67027, n62136, n186, n62132, n62128, n43051, 
        n25579, n27624, n69991, n69278, n62118, n51249, n37407, 
        n113, n62112, n56, n62_adj_5866, n51248, n51247, n51246, 
        n51245, n50682, n62106, n51244, n41_adj_5867, n51243, n62100, 
        n50898, n62098, n17_adj_5868, n50897, n51242, n51241, n50896, 
        n51240, n62092, n62090, n51239, n51238, n50681, n62088, 
        n50895, n5_adj_5869, n51237, n50680, n51236, n50894, n50297, 
        n67265, n51235, n51234, n51233, n60683, n58793, n54403, 
        n51232, n50679, n62074, n53323, n62068, n62062, n70252, 
        n62058, n51231, n51230, n50678, n51229, n50677, n26405, 
        n62046, n26306, n62040, n68749, n26235, n62036, n50676, 
        n50893, n51228, n51227, n50892, n51226, n50675, n50891, 
        n51225, n51224, n50890, n62030, n62028, n50889, n4_adj_5870, 
        n6_adj_5871, n8_adj_5872, n9_adj_5873, n4_adj_5874, n6_adj_5875, 
        n8_adj_5876, n9_adj_5877, n11_adj_5878, n13_adj_5879, n15_adj_5880, 
        n51223, n51222, n20935, n50888, n69976, n50314, n51221, 
        n50887, n51220, n50886, n51219, n51218, n51217, n38, n39, 
        n40, n41_adj_5881, n42, n43, n44, n45, n29404, n29403, 
        n29401, n51216, n50885, n50884, n50313, n50674, n50673, 
        n50883, n50882, n50672, n51215, n51214, n50671, n51213, 
        n50881, n50670, n50669, n51212, n51211, n50880, n11573, 
        n69300, n66980, n11571, n51210, n50879, n51209, n51208, 
        n51207, n51206, n69654, n70405, n29059, n57900, n57899, 
        n57898, n57897, n57896, n57895, n57894, n57893, n57892, 
        n57891, n57890, n57889, n57888, n57887, n57886, n57885, 
        n57884, n57883, n57882, n57881, n29037, n57880, n29035, 
        n29034, n57879, n29032, n57878, n29030, n58405, n57877, 
        n57876, n57875, n57874, n57873, n57872, n57871, n57870, 
        n57869, n63531, n58010, n58011, n28365, n28363, n28361, 
        n28358, n28355, n28352, n28338, n28804, n28310, n28308, 
        n28304, n28300, n53943, n51205, n51204, n51203, n50668, 
        n50312, n51202, n51201, n51200, n50667, n51199, n50666, 
        n51198, n50665, n51197, n66471, n51196, n51195, n51194, 
        n42234, n50664, n50663, n50662, n51193, n50661, n51192, 
        n50660, n50296, n51191, n51190, n51189, n51188, n51187, 
        n51186, n51185, n51184, n51183, n68423, n51182, n51181, 
        n51180, n51179, n51178, n51177, n29397, n51176, n20158, 
        n51175, n20112, n51174, n51173, n29394, n25819, n20159, 
        n50854, n51172, n51171, n50659, n42953, n51170, n29391, 
        n51169, n50658, n25460, n51168, n50853, n51167, n29388, 
        n29385, n43103, n51166, n50852, n50657, n57235, n57237, 
        n43101, n43099, n43095, n43093, n51165, n51164, n66452, 
        n68415, n51163, n51162, n51161, n51160, n50851, n50850, 
        n29901, n29898, n57868, n50849, n51159, n51158, n50848, 
        n51157, n50847, n51156, n51155, n51154, n50846, n50845, 
        n50656, n51153, n50844, n50655, n50843, n50654, n50653, 
        n50842, n51152, n50841, n50840, n51151, n51150, n51149, 
        n51148, n50652, n50839, n50651, n50650, n50838, n50649, 
        n50648, n51147, n60799, n50647, n51146, n50646, n50645, 
        n51145, n50644, n50643, n51144, n51143, n50837, n50642, 
        n51142, n51141, n50836, n51140, n50641, n50640, n14_adj_5882, 
        n50639, n51139, n50638, n51138, n51137, n50637, n10_adj_5883, 
        n51136, n2_adj_5884, n3_adj_5885, n4_adj_5886, n5_adj_5887, 
        n6_adj_5888, n7_adj_5889, n8_adj_5890, n9_adj_5891, n10_adj_5892, 
        n11_adj_5893, n12_adj_5894, n13_adj_5895, n14_adj_5896, n15_adj_5897, 
        n16_adj_5898, n17_adj_5899, n18_adj_5900, n19_adj_5901, n20_adj_5902, 
        n21_adj_5903, n22_adj_5904, n23_adj_5905, n24_adj_5906, n25_adj_5907, 
        n26_adj_5908, n27_adj_5909, n28_adj_5910, n29_adj_5911, n30_adj_5912, 
        n31_adj_5913, n32_adj_5914, n51135, n51134, n51133, n50636, 
        n51132, n50635, n51131, n51130, n50819, n51129, n50634, 
        n50818, n50633, n51128, n50817, n51127, n50816, n50632, 
        n51126, n51125, n50631, n50630, n51124, n50815, n50629, 
        n50628, n50627, n50814, n51123, n50626, n51122, n50625, 
        n51121, n50624, n50623, n69962, n50622, n51120, n50621, 
        n51119, n50620, n51118, n51117, n50619, n50813, n50618, 
        n50812, n50617, n50616, n51116, n51115, n50431, n50615, 
        n50811, n50810, n50614, n66446, n50430, n50001, n51114, 
        n51113, n66444, n59736, n50809, n50613, n50311, n50808, 
        n50612, n51112, n50611, n50807, n50806, n51111, n51110, 
        n48949, n50610, n50609, n50429, n50608, n50428, n51109, 
        n51108, n50607, n50805, n51543, n50804, n51107, n50606, 
        n51106, n50605, n50427, n50426, n50604, n66441, n51542, 
        n50803, n50603, n50310, n50425, n51541, n51540, n50802, 
        n50602, n50309, n51539, n51538, n51537, n50601, n4_adj_5915, 
        n50600, n50599, n50424, n50598, n50597, n50423, n50422, 
        n50295, n50596, n50421, n6_adj_5916, n50595, n50594, n42355, 
        n50420, n50419, n42880, n50418, n50417, n50416, n50415, 
        n50414, n50308, n50307, n50413, n51083, n51082, n50412, 
        n68443, n114, n50411, n51081, n50294, n51080, n51079, 
        n50410, n50409, n51078, n51077, n51076, n51075, n51074, 
        n41_adj_5917, n51073, n4_adj_5918, n51072, n51071, n50306, 
        n50305, n51070, n51069, n51068, n51067, n50560, n51066, 
        n51065, n50559, n50558, n51064, n50780, n50779, n51063, 
        n50557, n51062, n50778, n50556, n50777, n51061, n50555, 
        n50554, n51060, n50204, n50776, n50553, n50775, n50774, 
        n50773, n50552, n50293, n50292, n50551, n50322, n50550, 
        n50549, n50548, n42285, n50547, n50772, n50771, n50321, 
        n50304, n50770, n50546, n50769, n50303, n50768, n50545, 
        n50302, n50767, n42275, n50766, n50544, n50765, n50543, 
        n50542, n50301, n50320, n50541, n50540, n50764, n50539, 
        n50538, n50537, n50536, n50300, n50535, n50534, n50533, 
        n50532, n50319, n50318, n50317, n13_adj_5919, n15_adj_5920, 
        n110, n17_adj_5921, n19_adj_5922, n23_adj_5923, n29_adj_5924, 
        n31_adj_5925, n33, n61, n50531, n50530, n50529, n50528, 
        n50527, n50526, n50525, n51029, n51028, n51027, n20194, 
        n20897, n51026, n70399, n51025, n20185, n50749, n51024, 
        n51023, n50748, n51022, n57867, n61826, n63899, n51021, 
        n61820, n68671, n57866, n61814, n51020, n29017, n29016, 
        n29015, n51019, n61810, n51018, n51017, n50747, n12144, 
        n25961, n25771, n50746, n51016, n50745, n50744, n51015, 
        n51014, n57865, n51013, n50743, n50742, n50741, n51012, 
        n52894, n51011, n29013, n50740, n50739, n50738, n61804, 
        n25452, n68691, n50737, n61798, n51010, n70393, n61794, 
        n51009, n20113, n51008, n69620, n25544, n59833, n61788, 
        n52805, n60917, n61782, n26111, n51007, n61778, n70387, 
        n61772, n25566, n69892, n61766, n25705, n69661, n25676, 
        n61762, n57734, n69870, n70381, n69587, n68988, n61756, 
        n61750, n61746, n61740, n66396, n61734, n61730, n66389, 
        n66388, n61724, n61718, n61714, n4_adj_5926, n61708, n61702, 
        n62758, n63308, n17_adj_5927, n25_adj_5928, n56399, n5_adj_5929, 
        n24_adj_5930, n59785, n56483, n62752, n63312, n69845, n4_adj_5931, 
        n6_adj_5932, n58099, n58075, n4_adj_5933, n61049, n58366, 
        n56711, n58520, n58498, n58561, n58556, n22_adj_5934, n31_adj_5935, 
        n6_adj_5936, n58651, n58009, n58711, n63316, n59647, n58766, 
        n60713, n59714, n58008, n66302, n60784, n62698, n68056, 
        n61478, n62692, n61472, n4_adj_5937, n62684, n63547, n61043, 
        n59636, n62680, n59730, n57117, n59634, n57155, n70375, 
        n57159, n57163, n57167, n8_adj_5938, n57179, n57183, n57187, 
        n57191, n66280, n57195, n69555, n57199, n57203, n57207, 
        n57211, n57215, n57219, n57229, n57233, n69821, n58570, 
        n63903, n63900, n7_adj_5939, n70369, n69223, n61392, n59655, 
        n70569, n63665, n63663, n63662, n61190, n69222, n69152, 
        n69224, n70351, n63533, n57383, n69079, n61336, n10_adj_5940, 
        n69371, n4_adj_5941, n69045, n69534, n70363, n69797, n59716, 
        n69044, n68912, n68860, n69062, n69064, n7_adj_5942;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 encoder0_position_30__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n27624), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i29112_3_lut (.I0(n952), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n43039));
    defparam i29112_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut (.I0(n2722), .I1(n2724), .I2(n2728), .I3(GND_net), 
            .O(n62058));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i2_3_lut (.I0(encoder0_position[1]), .I1(n31), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i21_3_lut (.I0(encoder0_position[20]), .I1(n12_adj_5746), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n937));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4127[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n51176), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_25_lut (.I0(n69797), .I1(n2511), 
            .I2(VCC_net), .I3(n51029), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .timer({timer}), .GND_net(GND_net), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n29644(n29644), .n27799(n27799), .\bit_ctr[4] (bit_ctr[4]), 
            .n30294(n30294), .n30293(n30293), .n30292(n30292), .n30291(n30291), 
            .n30289(n30289), .n30288(n30288), .n30287(n30287), .n30286(n30286), 
            .n30285(n30285), .n30276(n30276), .n30187(n30187), .\bit_ctr[1] (bit_ctr[1]), 
            .n56711(n56711), .state({state}), .neopxl_color({neopxl_color}), 
            .\bit_ctr[0] (bit_ctr[0]), .NEOPXL_c(NEOPXL_c), .n110(n110), 
            .LED_c(LED_c), .n42981(n42981), .n52805(n52805), .n66110(n66110), 
            .\color_bit_N_502[1] (color_bit_N_502[1]), .n31(n31_adj_5935)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 encoder0_position_30__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n2720), .I1(n62058), .I2(n2726), .I3(n2725), 
            .O(n62062));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n11573_bdd_4_lut (.I0(n11573), .I1(current[15]), .I2(duty[22]), 
            .I3(n11571), .O(n70441));
    defparam n11573_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70441_bdd_4_lut (.I0(n70441), .I1(duty[19]), .I2(n4911), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[19]));
    defparam n70441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n2729), .I1(n43039), .I2(n2730), .I3(n2731), 
            .O(n59716));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11573_bdd_4_lut_54657 (.I0(n11573), .I1(current[15]), .I2(duty[21]), 
            .I3(n11571), .O(n70435));
    defparam n11573_bdd_4_lut_54657.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n50629));
    SB_LUT4 i53775_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69501));
    defparam i53775_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n3122), .I1(n3126), .I2(n3128), .I3(n3123), 
            .O(n62088));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1787 (.I0(n3119), .I1(n3120), .I2(n3125), .I3(GND_net), 
            .O(n62090));
    defparam i1_3_lut_adj_1787.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n51028), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n3121), .I1(n62088), .I2(n3124), .I3(n3127), 
            .O(n62092));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n59716), .I1(n2717), .I2(n2718), .I3(n62062), 
            .O(n62068));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_766_11_lut (.I0(n69976), .I1(n1125), 
            .I2(VCC_net), .I3(n50628), .O(n1224_adj_5836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i29184_4_lut (.I0(n956), .I1(n3131), .I2(n3132), .I3(n3133), 
            .O(n43111));
    defparam i29184_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n3117), .I1(n3118), .I2(n62092), .I3(n62090), 
            .O(n62098));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n3129), .I1(n62098), .I2(n43111), .I3(n3130), 
            .O(n62100));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n3114), .I1(n3115), .I2(n62100), .I3(n3116), 
            .O(n62106));
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n62106), 
            .O(n62112));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n62112), 
            .O(n62118));
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i53778_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n62118), 
            .O(n3138));
    defparam i53778_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5908));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n2712), .I1(n2710), .I2(n2719), .I3(n2721), 
            .O(n60917));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i3_3_lut (.I0(encoder0_position[2]), .I1(n30), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n2713), .I1(n2715), .I2(n2716), .I3(n62068), 
            .O(n62074));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53894_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69620));
    defparam i53894_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n3023), .I1(n3018), .I2(n3026), .I3(n3020), 
            .O(n62630));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1798 (.I0(n3021), .I1(n3019), .I2(n3027), .I3(GND_net), 
            .O(n62628));
    defparam i1_3_lut_adj_1798.LUT_INIT = 16'hfefe;
    SB_LUT4 i29120_4_lut (.I0(n955), .I1(n3031), .I2(n3032), .I3(n3033), 
            .O(n43047));
    defparam i29120_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n2709), .I1(n2714), .I2(n2727), .I3(n2723), 
            .O(n62272));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n3016), .I1(n62628), .I2(n3017), .I3(n62630), 
            .O(n62636));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'hfffe;
    SB_LUT4 i54011_4_lut (.I0(n2711), .I1(n62272), .I2(n62074), .I3(n60917), 
            .O(n2742));
    defparam i54011_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1801 (.I0(n3029), .I1(n62636), .I2(n43047), .I3(n3030), 
            .O(n62638));
    defparam i1_4_lut_adj_1801.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1802 (.I0(n3022), .I1(n3025), .I2(n3028), .I3(n3024), 
            .O(n62692));
    defparam i1_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n3010), .I1(n3011), .I2(n3014), .I3(n62638), 
            .O(n62644));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n3012), .I1(n3013), .I2(n3015), .I3(n62692), 
            .O(n62698));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n3008), .I1(n62698), .I2(n62644), .I3(n3009), 
            .O(n62648));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i53897_3_lut (.I0(n3007), .I1(n3006), .I2(n62648), .I3(GND_net), 
            .O(n3039));
    defparam i53897_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 encoder0_position_30__I_0_i1180_3_lut (.I0(n1729), .I1(n1796_adj_5851), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5907));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15635_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n22773), .I3(GND_net), .O(n29666));   // verilog/coms.v(130[12] 305[6])
    defparam i15635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15638_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n22773), .I3(GND_net), .O(n29669));   // verilog/coms.v(130[12] 305[6])
    defparam i15638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5906));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15640_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n22773), .I3(GND_net), .O(n29671));   // verilog/coms.v(130[12] 305[6])
    defparam i15640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15641_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3834), 
            .I3(GND_net), .O(n29672));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15642_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n22773), .I3(GND_net), .O(n29673));   // verilog/coms.v(130[12] 305[6])
    defparam i15642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15643_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n22773), .I3(GND_net), .O(n29674));   // verilog/coms.v(130[12] 305[6])
    defparam i15643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5905));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5904));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15645_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n22773), .I3(GND_net), .O(n29676));   // verilog/coms.v(130[12] 305[6])
    defparam i15645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5903));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n70435_bdd_4_lut (.I0(n70435), .I1(duty[18]), .I2(n4912), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[18]));
    defparam n70435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53861_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69587));
    defparam i53861_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(n2927), .I1(n2922), .I2(GND_net), .I3(GND_net), 
            .O(n62128));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n2926), .I1(n2921), .I2(n2925), .I3(n2928), 
            .O(n62132));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(n2923), .I1(n2920), .I2(n62128), .I3(n2924), 
            .O(n62136));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'hfffe;
    SB_LUT4 i29116_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n43043));
    defparam i29116_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n2918), .I1(n2919), .I2(n62136), .I3(n62132), 
            .O(n62142));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut (.I0(n58711), .I1(\data_out_frame[11] [0]), .I2(n58099), 
            .I3(n25676), .O(n14_adj_5725));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_out_frame[13] [2]), .I1(n14_adj_5725), .I2(n10_adj_5726), 
            .I3(\data_out_frame[11] [1]), .O(n25705));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(n2929), .I1(n43043), .I2(n2930), .I3(n2931), 
            .O(n59730));
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n2916), .I1(n59730), .I2(n2917), .I3(n62142), 
            .O(n62148));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n62148), 
            .O(n62154));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n62154), 
            .O(n62160));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 i53864_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n62160), 
            .O(n2940));
    defparam i53864_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5902));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15646_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n22773), .I3(GND_net), .O(n29677));   // verilog/coms.v(130[12] 305[6])
    defparam i15646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53928_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69654));
    defparam i53928_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1813 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58711));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1813.LUT_INIT = 16'h6666;
    SB_LUT4 i54008_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69734));
    defparam i54008_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i54040_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69766));
    defparam i54040_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15666_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n22773), .I3(GND_net), .O(n29697));   // verilog/coms.v(130[12] 305[6])
    defparam i15666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15670_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n22760), .I3(GND_net), .O(n29701));   // verilog/coms.v(130[12] 305[6])
    defparam i15670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35324_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[14]));
    defparam i35324_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1814 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1814.LUT_INIT = 16'h6666;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5927));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i15675_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3834), 
            .I3(GND_net), .O(n29706));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1972_22 (.CI(n51176), .I0(n2914), 
            .I1(VCC_net), .CO(n51177));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54071_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69797));
    defparam i54071_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n51175), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53935_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69661));
    defparam i53935_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5712));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53978_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69704));
    defparam i53978_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5711));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53808_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69534));
    defparam i53808_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1815 (.I0(n37154), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_1815.LUT_INIT = 16'h8888;
    SB_LUT4 i15677_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n22760), .I3(GND_net), .O(n29708));   // verilog/coms.v(130[12] 305[6])
    defparam i15677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_24 (.CI(n51028), .I0(n2512), 
            .I1(VCC_net), .CO(n51029));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54144_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69870));
    defparam i54144_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15681_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n22760), .I3(GND_net), .O(n29712));   // verilog/coms.v(130[12] 305[6])
    defparam i15681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54119_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69845));
    defparam i54119_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5901));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54095_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69821));
    defparam i54095_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1816 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58046));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1816.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1817 (.I0(\data_out_frame[5] [1]), .I1(n25666), 
            .I2(\data_out_frame[11] [7]), .I3(n58498), .O(n15_adj_5834));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1817.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5834), .I1(\data_out_frame[9] [5]), .I2(n14_adj_5835), 
            .I3(n58046), .O(n52894));   // verilog/coms.v(100[12:26])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15682_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n22760), .I3(GND_net), .O(n29713));   // verilog/coms.v(130[12] 305[6])
    defparam i15682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15683_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n22760), .I3(GND_net), .O(n29714));   // verilog/coms.v(130[12] 305[6])
    defparam i15683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1818 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58498));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1818.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53645_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69371));
    defparam i53645_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53829_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69555));
    defparam i53829_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1819 (.I0(n37050), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_5866));
    defparam i1_2_lut_adj_1819.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23183_3_lut (.I0(n214), .I1(IntegralLimit[18]), .I2(n156), 
            .I3(GND_net), .O(n37154));
    defparam i23183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_4306_i14_3_lut (.I0(encoder0_position[13]), .I1(n19_adj_5739), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n51027), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_21 (.CI(n51175), .I0(n2915), 
            .I1(VCC_net), .CO(n51176));
    SB_CARRY encoder0_position_30__I_0_add_1704_23 (.CI(n51027), .I0(n2513), 
            .I1(VCC_net), .CO(n51028));
    SB_LUT4 encoder0_position_30__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n50627), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n51026), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_10 (.CI(n50627), .I0(n1126), 
            .I1(VCC_net), .CO(n50628));
    SB_LUT4 mux_1587_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n12148));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5813));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_3_lut (.I0(n135), .I1(n187), .I2(n182), .I3(GND_net), 
            .O(n9_adj_5770));
    defparam i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(n9_adj_5770), .I1(IntegralLimit[20]), .I2(n156), 
            .I3(GND_net), .O(n37050));
    defparam i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1704_22 (.CI(n51026), .I0(n2514), 
            .I1(VCC_net), .CO(n51027));
    SB_LUT4 encoder0_position_30__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n51174), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n50626), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_9 (.CI(n50626), .I0(n1127), 
            .I1(VCC_net), .CO(n50627));
    SB_LUT4 encoder0_position_30__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n50625), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_766_8 (.CI(n50625), .I0(n1128), 
            .I1(VCC_net), .CO(n50626));
    SB_LUT4 i15366_3_lut (.I0(b_prev_adj_5783), .I1(b_new_adj_5989[1]), 
            .I2(debounce_cnt_N_3834_adj_5784), .I3(GND_net), .O(n29397));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821_adj_5856));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n11573_bdd_4_lut_54652 (.I0(n11573), .I1(current[15]), .I2(duty[20]), 
            .I3(n11571), .O(n70423));
    defparam n11573_bdd_4_lut_54652.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n51025), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n70423_bdd_4_lut (.I0(n70423), .I1(duty[17]), .I2(n4913), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[17]));
    defparam n70423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n50624), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15684_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n22760), .I3(GND_net), .O(n29715));   // verilog/coms.v(130[12] 305[6])
    defparam i15684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15685_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n22760), .I3(GND_net), .O(n29716));   // verilog/coms.v(130[12] 305[6])
    defparam i15685_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n2821_adj_5856), .I1(n2825), .I2(n2828), 
            .I3(n2824), .O(n62588));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_766_7 (.CI(n50624), .I0(n1129), 
            .I1(GND_net), .CO(n50625));
    SB_LUT4 encoder0_position_30__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n50623), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_6 (.CI(n50623), .I0(n1130), 
            .I1(GND_net), .CO(n50624));
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 n11573_bdd_4_lut_54643 (.I0(n11573), .I1(current[15]), .I2(duty[19]), 
            .I3(n11571), .O(n70417));
    defparam n11573_bdd_4_lut_54643.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5900));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n50622), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15370_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n22773), .I3(GND_net), .O(n29401));   // verilog/coms.v(130[12] 305[6])
    defparam i15370_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1704_21 (.CI(n51025), .I0(n2515), 
            .I1(VCC_net), .CO(n51026));
    SB_LUT4 i15686_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n22760), .I3(GND_net), .O(n29717));   // verilog/coms.v(130[12] 305[6])
    defparam i15686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15687_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n22760), .I3(GND_net), .O(n29718));   // verilog/coms.v(130[12] 305[6])
    defparam i15687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15688_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n22760), .I3(GND_net), .O(n29719));   // verilog/coms.v(130[12] 305[6])
    defparam i15688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16649_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n30680));   // verilog/coms.v(130[12] 305[6])
    defparam i16649_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15372_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n22773), .I3(GND_net), .O(n29403));   // verilog/coms.v(130[12] 305[6])
    defparam i15372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15689_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n22760), .I3(GND_net), .O(n29720));   // verilog/coms.v(130[12] 305[6])
    defparam i15689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54166_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69892));
    defparam i54166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1369_20_lut (.I0(n69821), .I1(n2016), 
            .I2(VCC_net), .I3(n50819), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1972_20 (.CI(n51174), .I0(n2916), 
            .I1(VCC_net), .CO(n51175));
    SB_LUT4 encoder0_position_30__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n51024), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n50818), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_19 (.CI(n50818), .I0(n2017), 
            .I1(VCC_net), .CO(n50819));
    SB_LUT4 encoder0_position_30__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n50817), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n51173), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_20 (.CI(n51024), .I0(n2516), 
            .I1(VCC_net), .CO(n51025));
    SB_LUT4 mux_4306_i11_3_lut (.I0(encoder0_position[10]), .I1(n22_adj_5736), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5899));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_30__I_0_add_766_5 (.CI(n50622), .I0(n1131), 
            .I1(VCC_net), .CO(n50623));
    SB_LUT4 i54299_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70025));
    defparam i54299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n50621), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n51023), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_19 (.CI(n51173), .I0(n2917), 
            .I1(VCC_net), .CO(n51174));
    SB_CARRY encoder0_position_30__I_0_add_1369_18 (.CI(n50817), .I0(n2018), 
            .I1(VCC_net), .CO(n50818));
    SB_LUT4 encoder0_position_30__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n50816), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_17 (.CI(n50816), .I0(n2019), 
            .I1(VCC_net), .CO(n50817));
    SB_LUT4 i15690_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n22760), .I3(GND_net), .O(n29721));   // verilog/coms.v(130[12] 305[6])
    defparam i15690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15691_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n22760), .I3(GND_net), .O(n29722));   // verilog/coms.v(130[12] 305[6])
    defparam i15691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_19 (.CI(n51023), .I0(n2517), 
            .I1(VCC_net), .CO(n51024));
    SB_LUT4 encoder0_position_30__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n51172), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1972_18 (.CI(n51172), .I0(n2918), 
            .I1(VCC_net), .CO(n51173));
    SB_LUT4 i15692_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n22760), .I3(GND_net), .O(n29723));   // verilog/coms.v(130[12] 305[6])
    defparam i15692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15693_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n22760), .I3(GND_net), .O(n29724));   // verilog/coms.v(130[12] 305[6])
    defparam i15693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54316_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70042));
    defparam i54316_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n50815), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n51022), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15694_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n22760), .I3(GND_net), .O(n29725));   // verilog/coms.v(130[12] 305[6])
    defparam i15694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15695_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n22760), .I3(GND_net), .O(n29726));   // verilog/coms.v(130[12] 305[6])
    defparam i15695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54281_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70007));
    defparam i54281_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1369_16 (.CI(n50815), .I0(n2020), 
            .I1(VCC_net), .CO(n50816));
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n51171), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15696_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n22760), .I3(GND_net), .O(n29727));   // verilog/coms.v(130[12] 305[6])
    defparam i15696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n70417_bdd_4_lut (.I0(n70417), .I1(duty[16]), .I2(n4914), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[16]));
    defparam n70417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5898));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1972_17 (.CI(n51171), .I0(n2919), 
            .I1(VCC_net), .CO(n51172));
    SB_LUT4 encoder0_position_30__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n50814), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_4 (.CI(n50621), .I0(n1132), 
            .I1(GND_net), .CO(n50622));
    SB_LUT4 encoder0_position_30__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n50620), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_18 (.CI(n51022), .I0(n2518), 
            .I1(VCC_net), .CO(n51023));
    SB_LUT4 encoder0_position_30__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n51170), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_16 (.CI(n51170), .I0(n2920), 
            .I1(VCC_net), .CO(n51171));
    SB_LUT4 encoder0_position_30__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n51021), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_3 (.CI(n50620), .I0(n1133), 
            .I1(VCC_net), .CO(n50621));
    SB_LUT4 encoder0_position_30__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n51169), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_15 (.CI(n50814), .I0(n2021), 
            .I1(VCC_net), .CO(n50815));
    SB_CARRY encoder0_position_30__I_0_add_1972_15 (.CI(n51169), .I0(n2921), 
            .I1(VCC_net), .CO(n51170));
    SB_LUT4 encoder0_position_30__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n50813), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_14 (.CI(n50813), .I0(n2022), 
            .I1(VCC_net), .CO(n50814));
    SB_LUT4 encoder0_position_30__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_17 (.CI(n51021), .I0(n2519), 
            .I1(VCC_net), .CO(n51022));
    SB_LUT4 encoder0_position_30__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n51020), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_16 (.CI(n51020), .I0(n2520), 
            .I1(VCC_net), .CO(n51021));
    SB_LUT4 encoder0_position_30__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n51019), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n50812), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_13 (.CI(n50812), .I0(n2023), 
            .I1(VCC_net), .CO(n50813));
    SB_LUT4 encoder0_position_30__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n51168), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_15 (.CI(n51019), .I0(n2521), 
            .I1(VCC_net), .CO(n51020));
    SB_LUT4 encoder0_position_30__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n50811), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n51018), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_12 (.CI(n50811), .I0(n2024), 
            .I1(VCC_net), .CO(n50812));
    SB_CARRY encoder0_position_30__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n50620));
    SB_LUT4 encoder0_position_30__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n50810), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n50619), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_14 (.CI(n51168), .I0(n2922), 
            .I1(VCC_net), .CO(n51169));
    SB_LUT4 encoder0_position_30__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n51167), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_14 (.CI(n51018), .I0(n2522), 
            .I1(VCC_net), .CO(n51019));
    SB_LUT4 encoder0_position_30__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n50618), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_9 (.CI(n50618), .I0(n1027), 
            .I1(VCC_net), .CO(n50619));
    SB_CARRY encoder0_position_30__I_0_add_1369_11 (.CI(n50810), .I0(n2025), 
            .I1(VCC_net), .CO(n50811));
    SB_LUT4 encoder0_position_30__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n50809), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_13 (.CI(n51167), .I0(n2923), 
            .I1(VCC_net), .CO(n51168));
    SB_LUT4 encoder0_position_30__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n51017), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27614_3_lut (.I0(n478), .I1(PWMLimit[4]), .I2(n406), .I3(GND_net), 
            .O(n7_adj_5855));
    defparam i27614_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1704_13 (.CI(n51017), .I0(n2523), 
            .I1(VCC_net), .CO(n51018));
    SB_CARRY encoder0_position_30__I_0_add_1369_10 (.CI(n50809), .I0(n2026), 
            .I1(VCC_net), .CO(n50810));
    SB_LUT4 encoder0_position_30__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n51016), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n50617), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_12 (.CI(n51016), .I0(n2524), 
            .I1(VCC_net), .CO(n51017));
    SB_CARRY encoder0_position_30__I_0_add_699_8 (.CI(n50617), .I0(n1028), 
            .I1(VCC_net), .CO(n50618));
    SB_LUT4 encoder0_position_30__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n50808), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_9 (.CI(n50808), .I0(n2027), 
            .I1(VCC_net), .CO(n50809));
    SB_LUT4 i27615_4_lut (.I0(setpoint[4]), .I1(n7_adj_5855), .I2(n15_adj_5808), 
            .I3(n405), .O(duty_23__N_3602[4]));
    defparam i27615_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 encoder0_position_30__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n51015), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_11 (.CI(n51015), .I0(n2525), 
            .I1(VCC_net), .CO(n51016));
    SB_LUT4 encoder0_position_30__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n50807), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_8 (.CI(n50807), .I0(n2028), 
            .I1(VCC_net), .CO(n50808));
    SB_LUT4 encoder0_position_30__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n50806), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_7 (.CI(n50806), .I0(n2029), 
            .I1(GND_net), .CO(n50807));
    SB_LUT4 encoder0_position_30__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n51014), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_10 (.CI(n51014), .I0(n2526), 
            .I1(VCC_net), .CO(n51015));
    SB_LUT4 encoder0_position_30__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n50805), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n50616), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_6 (.CI(n50805), .I0(n2030), 
            .I1(GND_net), .CO(n50806));
    SB_CARRY encoder0_position_30__I_0_add_699_7 (.CI(n50616), .I0(n1029), 
            .I1(GND_net), .CO(n50617));
    SB_LUT4 encoder0_position_30__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n50615), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_6 (.CI(n50615), .I0(n1030), 
            .I1(GND_net), .CO(n50616));
    SB_LUT4 encoder0_position_30__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n51013), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n50804), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n50614), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_5 (.CI(n50804), .I0(n2031), 
            .I1(VCC_net), .CO(n50805));
    SB_LUT4 encoder0_position_30__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n50803), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_5 (.CI(n50614), .I0(n1031), 
            .I1(VCC_net), .CO(n50615));
    SB_CARRY encoder0_position_30__I_0_add_1369_4 (.CI(n50803), .I0(n2032), 
            .I1(GND_net), .CO(n50804));
    SB_LUT4 encoder0_position_30__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n50613), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_4 (.CI(n50613), .I0(n1032), 
            .I1(GND_net), .CO(n50614));
    SB_LUT4 dti_counter_1938_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n51543), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n50612), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_3 (.CI(n50612), .I0(n1033), 
            .I1(VCC_net), .CO(n50613));
    SB_LUT4 dti_counter_1938_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n51542), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n50802), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1938_add_4_8 (.CI(n51542), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n51543));
    SB_LUT4 encoder0_position_30__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n51166), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_3 (.CI(n50802), .I0(n2033), 
            .I1(VCC_net), .CO(n50803));
    SB_LUT4 dti_counter_1938_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n51541), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_12 (.CI(n51166), .I0(n2924), 
            .I1(VCC_net), .CO(n51167));
    SB_CARRY encoder0_position_30__I_0_add_1704_9 (.CI(n51013), .I0(n2527), 
            .I1(VCC_net), .CO(n51014));
    SB_LUT4 encoder0_position_30__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54265_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69991));
    defparam i54265_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1821 (.I0(n2819), .I1(n2826), .I2(GND_net), .I3(GND_net), 
            .O(n62582));
    defparam i1_2_lut_adj_1821.LUT_INIT = 16'heeee;
    SB_CARRY dti_counter_1938_add_4_7 (.CI(n51541), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n51542));
    SB_LUT4 encoder0_position_30__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n51012), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_8 (.CI(n51012), .I0(n2528), 
            .I1(VCC_net), .CO(n51013));
    SB_LUT4 i15697_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n22760), .I3(GND_net), .O(n29728));   // verilog/coms.v(130[12] 305[6])
    defparam i15697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n51165), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_11 (.CI(n51165), .I0(n2925), 
            .I1(VCC_net), .CO(n51166));
    SB_CARRY encoder0_position_30__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n50802));
    SB_LUT4 encoder0_position_30__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n51011), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_7 (.CI(n51011), .I0(n2529), 
            .I1(GND_net), .CO(n51012));
    SB_LUT4 encoder0_position_30__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n51010), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n51164), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1938_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n51540), .O(n41_adj_5881)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1822 (.I0(n62588), .I1(n2820), .I2(n2823), .I3(GND_net), 
            .O(n62590));
    defparam i1_3_lut_adj_1822.LUT_INIT = 16'hfefe;
    SB_CARRY dti_counter_1938_add_4_6 (.CI(n51540), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n51541));
    SB_CARRY encoder0_position_30__I_0_add_1972_10 (.CI(n51164), .I0(n2926), 
            .I1(VCC_net), .CO(n51165));
    SB_CARRY encoder0_position_30__I_0_add_1704_6 (.CI(n51010), .I0(n2530), 
            .I1(GND_net), .CO(n51011));
    SB_LUT4 n11573_bdd_4_lut_54638 (.I0(n11573), .I1(current[15]), .I2(duty[18]), 
            .I3(n11571), .O(n70411));
    defparam n11573_bdd_4_lut_54638.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n51009), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1938_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n51539), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_5 (.CI(n51009), .I0(n2531), 
            .I1(VCC_net), .CO(n51010));
    SB_CARRY encoder0_position_30__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n50612));
    SB_LUT4 encoder0_position_30__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n50611), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n50610), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n51163), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1938_add_4_5 (.CI(n51539), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n51540));
    SB_CARRY encoder0_position_30__I_0_add_632_8 (.CI(n50610), .I0(n928), 
            .I1(VCC_net), .CO(n50611));
    SB_LUT4 n70411_bdd_4_lut (.I0(n70411), .I1(duty[15]), .I2(n4915), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[15]));
    defparam n70411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i27649_4_lut (.I0(setpoint[7]), .I1(n500), .I2(n15_adj_5808), 
            .I3(n405), .O(duty_23__N_3602[7]));
    defparam i27649_4_lut.LUT_INIT = 16'hca0a;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n50609), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_9 (.CI(n51163), .I0(n2927), 
            .I1(VCC_net), .CO(n51164));
    SB_LUT4 encoder0_position_30__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n51008), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n2818), .I1(n2822), .I2(n62582), .I3(n2827), 
            .O(n62592));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 dti_counter_1938_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n51538), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_4 (.CI(n51008), .I0(n2532), 
            .I1(GND_net), .CO(n51009));
    SB_LUT4 encoder0_position_30__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n51162), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n51007), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54250_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69976));
    defparam i54250_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_632_7 (.CI(n50609), .I0(n929), 
            .I1(GND_net), .CO(n50610));
    SB_LUT4 encoder0_position_30__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n50608), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_6 (.CI(n50608), .I0(n930), 
            .I1(GND_net), .CO(n50609));
    SB_CARRY encoder0_position_30__I_0_add_1704_3 (.CI(n51007), .I0(n2533), 
            .I1(VCC_net), .CO(n51008));
    SB_LUT4 encoder0_position_30__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n51007));
    SB_LUT4 i8753_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n20897));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i8753_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_30__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n50607), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_5 (.CI(n50607), .I0(n931), 
            .I1(VCC_net), .CO(n50608));
    SB_LUT4 encoder0_position_30__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n50606), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_8 (.CI(n51162), .I0(n2928), 
            .I1(VCC_net), .CO(n51163));
    SB_CARRY add_151_14 (.CI(n50303), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n50304));
    SB_LUT4 encoder0_position_30__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n51161), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7341_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i7341_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n11573_bdd_4_lut_54633 (.I0(n11573), .I1(current[15]), .I2(duty[17]), 
            .I3(n11571), .O(n70405));
    defparam n11573_bdd_4_lut_54633.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_632_4 (.CI(n50606), .I0(n932), 
            .I1(GND_net), .CO(n50607));
    SB_LUT4 i43156_3_lut (.I0(n4_adj_5937), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n58821));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i43156_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i15698_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n58010), 
            .I3(GND_net), .O(n29729));   // verilog/coms.v(130[12] 305[6])
    defparam i15698_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1972_7 (.CI(n51161), .I0(n2929), 
            .I1(GND_net), .CO(n51162));
    SB_LUT4 encoder0_position_30__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n50605), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n51160), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_6 (.CI(n51160), .I0(n2930), 
            .I1(GND_net), .CO(n51161));
    SB_LUT4 encoder0_position_30__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n51159), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_5 (.CI(n51159), .I0(n2931), 
            .I1(VCC_net), .CO(n51160));
    SB_CARRY encoder0_position_30__I_0_add_632_3 (.CI(n50605), .I0(n933), 
            .I1(VCC_net), .CO(n50606));
    SB_LUT4 encoder0_position_30__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n50605));
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n50294), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n50302), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n50604), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_151_13 (.CI(n50302), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n50303));
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5897));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27735), 
            .D(n1238), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27735), 
            .D(n1237), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i54236_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69962));
    defparam i54236_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n50603), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27735), 
            .D(n1236), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5896));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n51158), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_7 (.CI(n50603), .I0(n829), 
            .I1(GND_net), .CO(n50604));
    SB_CARRY encoder0_position_30__I_0_add_1972_4 (.CI(n51158), .I0(n2932), 
            .I1(GND_net), .CO(n51159));
    SB_CARRY dti_counter_1938_add_4_4 (.CI(n51538), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n51539));
    SB_LUT4 encoder0_position_30__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n51157), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n50602), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n70405_bdd_4_lut (.I0(n70405), .I1(duty[14]), .I2(n4916), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[14]));
    defparam n70405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_565_6 (.CI(n50602), .I0(n830), 
            .I1(GND_net), .CO(n50603));
    SB_CARRY encoder0_position_30__I_0_add_1972_3 (.CI(n51157), .I0(n2933), 
            .I1(VCC_net), .CO(n51158));
    SB_LUT4 encoder0_position_30__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n50601), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_5 (.CI(n50601), .I0(n831), 
            .I1(VCC_net), .CO(n50602));
    SB_LUT4 encoder0_position_30__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n50600), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_565_4 (.CI(n50600), .I0(n832), 
            .I1(GND_net), .CO(n50601));
    SB_LUT4 dti_counter_1938_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n51537), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n50599), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n51157));
    SB_CARRY encoder0_position_30__I_0_add_565_3 (.CI(n50599), .I0(n833), 
            .I1(VCC_net), .CO(n50600));
    SB_LUT4 encoder0_position_30__I_0_add_1905_28_lut (.I0(n69654), .I1(n2808), 
            .I2(VCC_net), .I3(n51156), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n51155), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_27 (.CI(n51155), .I0(n2809), 
            .I1(VCC_net), .CO(n51156));
    SB_LUT4 encoder0_position_30__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n50599));
    SB_LUT4 encoder0_position_30__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n51154), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2457_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n50598), 
            .O(n7444)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2457_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2457_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n50597), 
            .O(n7445)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2457_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_26 (.CI(n51154), .I0(n2810), 
            .I1(VCC_net), .CO(n51155));
    SB_LUT4 encoder0_position_30__I_0_add_1302_19_lut (.I0(n69371), .I1(n1917), 
            .I2(VCC_net), .I3(n50780), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n50779), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_18 (.CI(n50779), .I0(n1918), 
            .I1(VCC_net), .CO(n50780));
    SB_CARRY add_2457_6 (.CI(n50597), .I0(n622), .I1(GND_net), .CO(n50598));
    SB_LUT4 encoder0_position_30__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n50778), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2457_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n50596), 
            .O(n7446)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2457_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2457_5 (.CI(n50596), .I0(n623), .I1(VCC_net), .CO(n50597));
    SB_CARRY dti_counter_1938_add_4_3 (.CI(n51537), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n51538));
    SB_CARRY encoder0_position_30__I_0_add_1302_17 (.CI(n50778), .I0(n1919), 
            .I1(VCC_net), .CO(n50779));
    SB_LUT4 encoder0_position_30__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n50777), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2457_4_lut (.I0(GND_net), .I1(n405_adj_5787), .I2(GND_net), 
            .I3(n50595), .O(n7447)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2457_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n51153), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2457_4 (.CI(n50595), .I0(n405_adj_5787), .I1(GND_net), 
            .CO(n50596));
    SB_LUT4 add_2457_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n50594), 
            .O(n7448)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2457_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_25 (.CI(n51153), .I0(n2811), 
            .I1(VCC_net), .CO(n51154));
    SB_CARRY encoder0_position_30__I_0_add_1302_16 (.CI(n50777), .I0(n1920), 
            .I1(VCC_net), .CO(n50778));
    SB_LUT4 encoder0_position_30__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n50776), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_15 (.CI(n50776), .I0(n1921), 
            .I1(VCC_net), .CO(n50777));
    SB_LUT4 encoder0_position_30__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n50775), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2457_3 (.CI(n50594), .I0(n625), .I1(VCC_net), .CO(n50595));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5895));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1302_14 (.CI(n50775), .I0(n1922), 
            .I1(VCC_net), .CO(n50776));
    SB_LUT4 encoder0_position_30__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n51152), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_24 (.CI(n51152), .I0(n2812), 
            .I1(VCC_net), .CO(n51153));
    SB_LUT4 add_2457_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7449)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2457_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n50774), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1938_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1938_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_13 (.CI(n50774), .I0(n1923), 
            .I1(VCC_net), .CO(n50775));
    SB_LUT4 encoder0_position_30__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n50773), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n51151), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1302_12 (.CI(n50773), .I0(n1924), 
            .I1(VCC_net), .CO(n50774));
    SB_CARRY encoder0_position_30__I_0_add_1905_23 (.CI(n51151), .I0(n2813), 
            .I1(VCC_net), .CO(n51152));
    SB_LUT4 encoder0_position_30__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n50772), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n51150), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_11 (.CI(n50772), .I0(n1925), 
            .I1(VCC_net), .CO(n50773));
    SB_LUT4 encoder0_position_30__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n50771), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_22 (.CI(n51150), .I0(n2814), 
            .I1(VCC_net), .CO(n51151));
    SB_CARRY encoder0_position_30__I_0_add_1302_10 (.CI(n50771), .I0(n1926), 
            .I1(VCC_net), .CO(n50772));
    SB_LUT4 encoder0_position_30__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n50770), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_9 (.CI(n50770), .I0(n1927), 
            .I1(VCC_net), .CO(n50771));
    SB_CARRY add_2457_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n50594));
    SB_LUT4 encoder0_position_30__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n50769), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_8 (.CI(n50769), .I0(n1928), 
            .I1(VCC_net), .CO(n50770));
    SB_LUT4 encoder0_position_30__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n50768), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4306_i15_3_lut (.I0(encoder0_position[14]), .I1(n18_adj_5740), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1302_7 (.CI(n50768), .I0(n1929), 
            .I1(GND_net), .CO(n50769));
    SB_LUT4 encoder0_position_30__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n50767), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_6 (.CI(n50767), .I0(n1930), 
            .I1(GND_net), .CO(n50768));
    SB_LUT4 encoder0_position_30__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n50766), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_5 (.CI(n50766), .I0(n1931), 
            .I1(VCC_net), .CO(n50767));
    SB_CARRY dti_counter_1938_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n51537));
    SB_LUT4 encoder0_position_30__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n50765), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n51149), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_24_lut (.I0(n69704), .I1(n2412), 
            .I2(VCC_net), .I3(n50986), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1302_4 (.CI(n50765), .I0(n1932), 
            .I1(GND_net), .CO(n50766));
    SB_CARRY encoder0_position_30__I_0_add_1905_21 (.CI(n51149), .I0(n2815), 
            .I1(VCC_net), .CO(n51150));
    SB_LUT4 encoder0_position_30__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n50764), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1302_3 (.CI(n50764), .I0(n1933), 
            .I1(VCC_net), .CO(n50765));
    SB_LUT4 encoder0_position_30__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n50985), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_23 (.CI(n50985), .I0(n2413), 
            .I1(VCC_net), .CO(n50986));
    SB_LUT4 encoder0_position_30__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n50764));
    SB_LUT4 encoder0_position_30__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29027_3_lut (.I0(n953), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n42953));
    defparam i29027_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61043), .O(n61472));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61472), .O(n61478));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n50984), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n51148), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_22 (.CI(n50984), .I0(n2414), 
            .I1(VCC_net), .CO(n50985));
    SB_LUT4 encoder0_position_30__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n50983), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_21 (.CI(n50983), .I0(n2415), 
            .I1(VCC_net), .CO(n50984));
    SB_LUT4 encoder0_position_30__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1905_20 (.CI(n51148), .I0(n2816), 
            .I1(VCC_net), .CO(n51149));
    SB_LUT4 encoder0_position_30__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n50982), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n51147), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1905_19 (.CI(n51147), .I0(n2817), 
            .I1(VCC_net), .CO(n51148));
    SB_CARRY encoder0_position_30__I_0_add_1637_20 (.CI(n50982), .I0(n2416), 
            .I1(VCC_net), .CO(n50983));
    SB_LUT4 encoder0_position_30__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n50981), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n51146), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_19 (.CI(n50981), .I0(n2417), 
            .I1(VCC_net), .CO(n50982));
    SB_LUT4 i15678_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n58010), 
            .I3(GND_net), .O(n29709));   // verilog/coms.v(130[12] 305[6])
    defparam i15678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29154_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n43081));
    defparam i29154_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5894));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29256_4_lut (.I0(n829), .I1(n828), .I2(n43081), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i29256_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i43130_3_lut (.I0(n4_adj_5776), .I1(n7446), .I2(n58792), .I3(GND_net), 
            .O(n58795));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n50980), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i43131_3_lut (.I0(encoder0_position[28]), .I1(n58795), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29158_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n43085));
    defparam i29158_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_30__I_0_add_1905_18 (.CI(n51146), .I0(n2818), 
            .I1(VCC_net), .CO(n51147));
    SB_LUT4 encoder0_position_30__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n51145), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_18 (.CI(n50980), .I0(n2418), 
            .I1(VCC_net), .CO(n50981));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5893));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1905_17 (.CI(n51145), .I0(n2819), 
            .I1(VCC_net), .CO(n51146));
    SB_LUT4 encoder0_position_30__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n50979), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n51144), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_16 (.CI(n51144), .I0(n2820), 
            .I1(VCC_net), .CO(n51145));
    SB_CARRY encoder0_position_30__I_0_add_1637_17 (.CI(n50979), .I0(n2419), 
            .I1(VCC_net), .CO(n50980));
    SB_LUT4 encoder0_position_30__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821_adj_5856), 
            .I2(VCC_net), .I3(n51143), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n50978), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1826 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n62320));
    defparam i1_2_lut_adj_1826.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_1637_16 (.CI(n50978), .I0(n2420), 
            .I1(VCC_net), .CO(n50979));
    SB_LUT4 encoder0_position_30__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n50977), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_15 (.CI(n51143), .I0(n2821_adj_5856), 
            .I1(VCC_net), .CO(n51144));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5892));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n927), .I1(n62320), .I2(n928), .I3(n43085), 
            .O(n960));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_30__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n51142), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_14 (.CI(n51142), .I0(n2822), 
            .I1(VCC_net), .CO(n51143));
    SB_LUT4 encoder0_position_30__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n51141), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1637_15 (.CI(n50977), .I0(n2421), 
            .I1(VCC_net), .CO(n50978));
    SB_LUT4 n11573_bdd_4_lut_54628 (.I0(n11573), .I1(current[15]), .I2(duty[16]), 
            .I3(n11571), .O(n70399));
    defparam n11573_bdd_4_lut_54628.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n50976), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5891));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1905_13 (.CI(n51141), .I0(n2823), 
            .I1(VCC_net), .CO(n51142));
    SB_LUT4 encoder0_position_30__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n51140), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_14 (.CI(n50976), .I0(n2422), 
            .I1(VCC_net), .CO(n50977));
    SB_LUT4 encoder0_position_30__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n50975), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_12 (.CI(n51140), .I0(n2824), 
            .I1(VCC_net), .CO(n51141));
    SB_CARRY encoder0_position_30__I_0_add_1637_13 (.CI(n50975), .I0(n2423), 
            .I1(VCC_net), .CO(n50976));
    SB_LUT4 i29068_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n42995));
    defparam i29068_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5884), .I3(n51771), .O(n2_adj_5778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n50974), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_12 (.CI(n50974), .I0(n2424), 
            .I1(VCC_net), .CO(n50975));
    SB_LUT4 encoder0_position_30__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n51139), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n50973), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_18_lut (.I0(n69555), .I1(n1818), 
            .I2(VCC_net), .I3(n50749), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1637_11 (.CI(n50973), .I0(n2425), 
            .I1(VCC_net), .CO(n50974));
    SB_LUT4 encoder0_position_30__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n50748), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5885), .I3(n51770), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_32 (.CI(n51770), 
            .I0(GND_net), .I1(n3_adj_5885), .CO(n51771));
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_30__I_0_add_1235_17 (.CI(n50748), .I0(n1819), 
            .I1(VCC_net), .CO(n50749));
    SB_LUT4 n70399_bdd_4_lut (.I0(n70399), .I1(duty[13]), .I2(n4917), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[13]));
    defparam n70399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n2816), .I1(n2817), .I2(n62592), .I3(n62590), 
            .O(n62598));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 n11573_bdd_4_lut_54623 (.I0(n11573), .I1(current[15]), .I2(duty[15]), 
            .I3(n11571), .O(n70393));
    defparam n11573_bdd_4_lut_54623.LUT_INIT = 16'he4aa;
    SB_LUT4 n70393_bdd_4_lut (.I0(n70393), .I1(duty[12]), .I2(n4918), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[12]));
    defparam n70393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n2829), .I1(n42953), .I2(n2830), .I3(n2831), 
            .O(n59761));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'ha080;
    SB_LUT4 n11573_bdd_4_lut_54618 (.I0(n11573), .I1(current[11]), .I2(duty[14]), 
            .I3(n11571), .O(n70387));
    defparam n11573_bdd_4_lut_54618.LUT_INIT = 16'he4aa;
    SB_LUT4 n70387_bdd_4_lut (.I0(n70387), .I1(duty[11]), .I2(n4919), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[11]));
    defparam n70387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n2814), .I1(n2815), .I2(n59761), .I3(n62598), 
            .O(n62604));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'hfffe;
    SB_LUT4 n11573_bdd_4_lut_54613 (.I0(n11573), .I1(current[10]), .I2(duty[13]), 
            .I3(n11571), .O(n70381));
    defparam n11573_bdd_4_lut_54613.LUT_INIT = 16'he4aa;
    SB_LUT4 n70381_bdd_4_lut (.I0(n70381), .I1(duty[10]), .I2(n4920), 
            .I3(n11571), .O(pwm_setpoint_23__N_3[10]));
    defparam n70381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n62604), 
            .O(n62610));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    SB_LUT4 n11573_bdd_4_lut_54608 (.I0(n11573), .I1(current[9]), .I2(duty[12]), 
            .I3(n11571), .O(n70375));
    defparam n11573_bdd_4_lut_54608.LUT_INIT = 16'he4aa;
    SB_LUT4 n70375_bdd_4_lut (.I0(n70375), .I1(duty[9]), .I2(n4921), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n70375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i53931_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n62610), 
            .O(n2841));
    defparam i53931_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n11573_bdd_4_lut_54603 (.I0(n11573), .I1(current[8]), .I2(duty[11]), 
            .I3(n11571), .O(n70369));
    defparam n11573_bdd_4_lut_54603.LUT_INIT = 16'he4aa;
    SB_LUT4 n70369_bdd_4_lut (.I0(n70369), .I1(duty[8]), .I2(n4922), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n70369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11573_bdd_4_lut_54598 (.I0(n11573), .I1(current[7]), .I2(duty[10]), 
            .I3(n11571), .O(n70363));
    defparam n11573_bdd_4_lut_54598.LUT_INIT = 16'he4aa;
    SB_LUT4 n70363_bdd_4_lut (.I0(n70363), .I1(duty[7]), .I2(n4923), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n70363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11573_bdd_4_lut_54593 (.I0(n11573), .I1(current[6]), .I2(duty[9]), 
            .I3(n11571), .O(n70357));
    defparam n11573_bdd_4_lut_54593.LUT_INIT = 16'he4aa;
    SB_LUT4 n70357_bdd_4_lut (.I0(n70357), .I1(duty[6]), .I2(n4924), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n70357_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11573_bdd_4_lut_54588 (.I0(n11573), .I1(current[5]), .I2(duty[8]), 
            .I3(n11571), .O(n70351));
    defparam n11573_bdd_4_lut_54588.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1905_11 (.CI(n51139), .I0(n2825), 
            .I1(VCC_net), .CO(n51140));
    SB_LUT4 i15572_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n58009), 
            .I3(GND_net), .O(n29603));   // verilog/coms.v(130[12] 305[6])
    defparam i15572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5886), .I3(n51769), .O(n4_adj_5776)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5890));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n50972), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5889));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5888));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_31 (.CI(n51769), 
            .I0(GND_net), .I1(n4_adj_5886), .CO(n51770));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5887), .I3(n51768), .O(n5_adj_5775)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n50747), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n1029), .I1(n42995), .I2(n1030), .I3(n1031), 
            .O(n59639));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_30 (.CI(n51768), 
            .I0(GND_net), .I1(n5_adj_5887), .CO(n51769));
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27735), 
            .D(n1235), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5888), .I3(n51767), .O(n6_adj_5753)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54239_4_lut (.I0(n1026), .I1(n59639), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i54239_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29074_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n43001));
    defparam i29074_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1833 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n62236));
    defparam i1_3_lut_adj_1833.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1834 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n62328));
    defparam i1_2_lut_adj_1834.LUT_INIT = 16'h8888;
    SB_LUT4 i54253_4_lut (.I0(n62328), .I1(n1125), .I2(n62236), .I3(n43001), 
            .O(n1158));
    defparam i54253_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_30__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29076_3_lut (.I0(n937), .I1(n1232_adj_5844), .I2(n1233_adj_5845), 
            .I3(GND_net), .O(n43003));
    defparam i29076_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1835 (.I0(n1226_adj_5838), .I1(n1227_adj_5839), 
            .I2(n1228_adj_5840), .I3(GND_net), .O(n62350));
    defparam i1_3_lut_adj_1835.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n1229_adj_5841), .I1(n43003), .I2(n1230_adj_5842), 
            .I3(n1231_adj_5843), .O(n59636));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'ha080;
    SB_LUT4 i54268_4_lut (.I0(n1225_adj_5837), .I1(n1224_adj_5836), .I2(n59636), 
            .I3(n62350), .O(n1257));
    defparam i54268_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226_adj_5838));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29070_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n42997));
    defparam i29070_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n62198));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(n1329), .I1(n42997), .I2(n1330), .I3(n1331), 
            .O(n59634));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'ha080;
    SB_LUT4 i54284_4_lut (.I0(n59634), .I1(n1323), .I2(n1324), .I3(n62198), 
            .O(n1356));
    defparam i54284_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i837_3_lut (.I0(n1226_adj_5838), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29080_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n43007));
    defparam i29080_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1839 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n62360));
    defparam i1_2_lut_adj_1839.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(n1429), .I1(n43007), .I2(n1430), .I3(n1431), 
            .O(n59647));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1841 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n62360), 
            .O(n62366));
    defparam i1_4_lut_adj_1841.LUT_INIT = 16'hfffe;
    SB_LUT4 n70351_bdd_4_lut (.I0(n70351), .I1(duty[5]), .I2(n4925), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n70351_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1842 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5941));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'h7bde;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_29 (.CI(n51767), 
            .I0(GND_net), .I1(n6_adj_5888), .CO(n51768));
    SB_LUT4 encoder0_position_30__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n51138), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5887));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5889), .I3(n51766), .O(n7_adj_5752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_16 (.CI(n50747), .I0(n1820), 
            .I1(VCC_net), .CO(n50748));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_28 (.CI(n51766), 
            .I0(GND_net), .I1(n7_adj_5889), .CO(n51767));
    SB_LUT4 encoder0_position_30__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n50746), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_10 (.CI(n50972), .I0(n2426), 
            .I1(VCC_net), .CO(n50973));
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27735), 
            .D(n1234), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27735), 
            .D(n1233), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27735), 
            .D(n1232), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27735), 
            .D(n1231), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_CARRY encoder0_position_30__I_0_add_1235_15 (.CI(n50746), .I0(n1821), 
            .I1(VCC_net), .CO(n50747));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5890), .I3(n51765), .O(n8_adj_5751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n50971), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822_adj_5852), 
            .I2(VCC_net), .I3(n50745), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_10 (.CI(n51138), .I0(n2826), 
            .I1(VCC_net), .CO(n51139));
    SB_LUT4 encoder0_position_30__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n51137), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_14 (.CI(n50745), .I0(n1822_adj_5852), 
            .I1(VCC_net), .CO(n50746));
    SB_CARRY encoder0_position_30__I_0_add_1905_9 (.CI(n51137), .I0(n2827), 
            .I1(VCC_net), .CO(n51138));
    SB_LUT4 encoder0_position_30__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n50744), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_9 (.CI(n50971), .I0(n2427), 
            .I1(VCC_net), .CO(n50972));
    SB_CARRY encoder0_position_30__I_0_add_1235_13 (.CI(n50744), .I0(n1823), 
            .I1(VCC_net), .CO(n50745));
    SB_LUT4 encoder0_position_30__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n50970), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5886));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n51136), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_8 (.CI(n51136), .I0(n2828), 
            .I1(VCC_net), .CO(n51137));
    SB_LUT4 encoder0_position_30__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824_adj_5853), 
            .I2(VCC_net), .I3(n50743), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_12 (.CI(n50743), .I0(n1824_adj_5853), 
            .I1(VCC_net), .CO(n50744));
    SB_CARRY encoder0_position_30__I_0_add_1637_8 (.CI(n50970), .I0(n2428), 
            .I1(VCC_net), .CO(n50971));
    SB_LUT4 encoder0_position_30__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n51135), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_7 (.CI(n51135), .I0(n2829), 
            .I1(GND_net), .CO(n51136));
    SB_LUT4 encoder0_position_30__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n50742), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_27 (.CI(n51765), 
            .I0(GND_net), .I1(n8_adj_5890), .CO(n51766));
    SB_CARRY encoder0_position_30__I_0_add_1235_11 (.CI(n50742), .I0(n1825), 
            .I1(VCC_net), .CO(n50743));
    SB_LUT4 encoder0_position_30__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n50969), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5885));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5891), .I3(n51764), .O(n9_adj_5750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_26 (.CI(n51764), 
            .I0(GND_net), .I1(n9_adj_5891), .CO(n51765));
    SB_LUT4 encoder0_position_30__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n50741), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n51134), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_7 (.CI(n50969), .I0(n2429), 
            .I1(GND_net), .CO(n50970));
    SB_CARRY encoder0_position_30__I_0_add_1235_10 (.CI(n50741), .I0(n1826), 
            .I1(VCC_net), .CO(n50742));
    SB_LUT4 encoder0_position_30__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n50968), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n50740), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_9 (.CI(n50740), .I0(n1827), 
            .I1(VCC_net), .CO(n50741));
    SB_CARRY encoder0_position_30__I_0_add_1637_6 (.CI(n50968), .I0(n2430), 
            .I1(GND_net), .CO(n50969));
    SB_LUT4 encoder0_position_30__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n50739), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_6 (.CI(n51134), .I0(n2830), 
            .I1(GND_net), .CO(n51135));
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27735), 
            .D(n1230), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n51133), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11573_bdd_4_lut_54583 (.I0(n11573), .I1(current[4]), .I2(duty[7]), 
            .I3(n11571), .O(n70345));
    defparam n11573_bdd_4_lut_54583.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5892), .I3(n51763), .O(n10_adj_5748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n50967), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_8 (.CI(n50739), .I0(n1828), 
            .I1(VCC_net), .CO(n50740));
    SB_CARRY encoder0_position_30__I_0_add_1637_5 (.CI(n50967), .I0(n2431), 
            .I1(VCC_net), .CO(n50968));
    SB_LUT4 encoder0_position_30__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n50966), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n50738), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_5 (.CI(n51133), .I0(n2831), 
            .I1(VCC_net), .CO(n51134));
    SB_CARRY encoder0_position_30__I_0_add_1637_4 (.CI(n50966), .I0(n2432), 
            .I1(GND_net), .CO(n50967));
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_25 (.CI(n51763), 
            .I0(GND_net), .I1(n10_adj_5892), .CO(n51764));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5893), .I3(n51762), .O(n11_adj_5747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_7 (.CI(n50738), .I0(n1829), 
            .I1(GND_net), .CO(n50739));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5884));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_24 (.CI(n51762), 
            .I0(GND_net), .I1(n11_adj_5893), .CO(n51763));
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n50965), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n51132), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5894), .I3(n51761), .O(n12_adj_5746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54319_4_lut (.I0(n1423), .I1(n1422), .I2(n62366), .I3(n59647), 
            .O(n1455));
    defparam i54319_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n70345_bdd_4_lut (.I0(n70345), .I1(duty[4]), .I2(n4926), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n70345_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_23 (.CI(n51761), 
            .I0(GND_net), .I1(n12_adj_5894), .CO(n51762));
    SB_CARRY encoder0_position_30__I_0_add_1905_4 (.CI(n51132), .I0(n2832), 
            .I1(GND_net), .CO(n51133));
    SB_CARRY encoder0_position_30__I_0_add_1637_3 (.CI(n50965), .I0(n2433), 
            .I1(VCC_net), .CO(n50966));
    SB_LUT4 encoder0_position_30__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n50965));
    SB_LUT4 encoder0_position_30__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n50737), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_6 (.CI(n50737), .I0(n1830), 
            .I1(GND_net), .CO(n50738));
    SB_LUT4 encoder0_position_30__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n50736), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_5 (.CI(n50736), .I0(n1831), 
            .I1(VCC_net), .CO(n50737));
    SB_LUT4 encoder0_position_30__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n50735), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_4 (.CI(n50735), .I0(n1832), 
            .I1(GND_net), .CO(n50736));
    SB_LUT4 encoder0_position_30__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n50734), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1235_3 (.CI(n50734), .I0(n1833), 
            .I1(VCC_net), .CO(n50735));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5895), .I3(n51760), .O(n13_adj_5745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n51131), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_3 (.CI(n51131), .I0(n2833), 
            .I1(VCC_net), .CO(n51132));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_22 (.CI(n51760), 
            .I0(GND_net), .I1(n13_adj_5895), .CO(n51761));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5896), .I3(n51759), .O(n14_adj_5744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1843 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n62204));
    defparam i1_2_lut_adj_1843.LUT_INIT = 16'heeee;
    SB_LUT4 i29086_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n43013));
    defparam i29086_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i22928_3_lut (.I0(n219), .I1(IntegralLimit[13]), .I2(n156), 
            .I3(GND_net), .O(n244));
    defparam i22928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1844 (.I0(n244), .I1(Ki[0]), .I2(GND_net), .I3(GND_net), 
            .O(n41_adj_5867));
    defparam i1_2_lut_adj_1844.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_25_lut (.I0(n69962), .I1(n2_adj_5884), .I2(n1059), 
            .I3(n51294), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 n11573_bdd_4_lut_54578 (.I0(n11573), .I1(current[3]), .I2(duty[6]), 
            .I3(n11571), .O(n70339));
    defparam n11573_bdd_4_lut_54578.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_21 (.CI(n51759), 
            .I0(GND_net), .I1(n14_adj_5896), .CO(n51760));
    SB_CARRY encoder0_position_30__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n50734));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5897), .I3(n51758), .O(n15_adj_5743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5883));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i6_4_lut_adj_1845 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5882));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n58821));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i7_4_lut_adj_1846 (.I0(dti_counter[0]), .I1(n14_adj_5882), .I2(n10_adj_5883), 
            .I3(dti_counter[3]), .O(n22841));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n51131));
    SB_LUT4 add_2507_24_lut (.I0(n69976), .I1(n2_adj_5884), .I2(n1158), 
            .I3(n51293), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15672_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n58009), 
            .I3(GND_net), .O(n29703));   // verilog/coms.v(130[12] 305[6])
    defparam i15672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_27_lut (.I0(GND_net), .I1(n2709), 
            .I2(VCC_net), .I3(n51130), .O(n2776)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n51129), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n50322), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1847 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n62204), 
            .O(n62210));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY add_2507_24 (.CI(n51293), .I0(n2_adj_5884), .I1(n1158), .CO(n51294));
    SB_CARRY encoder0_position_30__I_0_add_1838_26 (.CI(n51129), .I0(n2710), 
            .I1(VCC_net), .CO(n51130));
    SB_LUT4 i1_4_lut_adj_1848 (.I0(n1529), .I1(n62210), .I2(n43013), .I3(n1530), 
            .O(n62212));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'heccc;
    SB_LUT4 add_2507_23_lut (.I0(n69991), .I1(n2_adj_5884), .I2(n1257), 
            .I3(n51292), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n50301), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n51128), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_25 (.CI(n51128), .I0(n2711), 
            .I1(VCC_net), .CO(n51129));
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n50321), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_23 (.CI(n51292), .I0(n2_adj_5884), .I1(n1257), .CO(n51293));
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n51127), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i54302_4_lut (.I0(n1522), .I1(n1521), .I2(n62212), .I3(n1523), 
            .O(n1554));
    defparam i54302_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_20 (.CI(n51758), 
            .I0(GND_net), .I1(n15_adj_5897), .CO(n51759));
    SB_LUT4 i54226_2_lut (.I0(n22841), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i54226_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5898), .I3(n51757), .O(n16_adj_5742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n70339_bdd_4_lut (.I0(n70339), .I1(duty[3]), .I2(n4927), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n70339_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_1838_24 (.CI(n51127), .I0(n2712), 
            .I1(VCC_net), .CO(n51128));
    SB_LUT4 encoder0_position_30__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n51126), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_22_lut (.I0(n70007), .I1(n2_adj_5884), .I2(n1356), 
            .I3(n51291), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_22_lut.LUT_INIT = 16'h8BB8;
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1838_23 (.CI(n51126), .I0(n2713), 
            .I1(VCC_net), .CO(n51127));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_19 (.CI(n51757), 
            .I0(GND_net), .I1(n16_adj_5898), .CO(n51758));
    SB_CARRY add_2507_22 (.CI(n51291), .I0(n2_adj_5884), .I1(n1356), .CO(n51292));
    SB_LUT4 encoder0_position_30__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n51125), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_21_lut (.I0(n70042), .I1(n2_adj_5884), .I2(n1455), 
            .I3(n51290), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_21 (.CI(n51290), .I0(n2_adj_5884), .I1(n1455), .CO(n51291));
    SB_CARRY encoder0_position_30__I_0_add_1838_22 (.CI(n51125), .I0(n2714), 
            .I1(VCC_net), .CO(n51126));
    SB_LUT4 encoder0_position_30__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28999_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n42925));
    defparam i28999_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(n1629), .I1(n42925), .I2(n1630), .I3(n1631), 
            .O(n59655));
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'ha080;
    SB_LUT4 add_2507_20_lut (.I0(n70025), .I1(n2_adj_5884), .I2(n1554), 
            .I3(n51289), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5899), .I3(n51756), .O(n17_adj_5741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_20 (.CI(n51289), .I0(n2_adj_5884), .I1(n1554), .CO(n51290));
    SB_LUT4 add_2507_19_lut (.I0(n69892), .I1(n2_adj_5884), .I2(n1653), 
            .I3(n51288), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1850 (.I0(n1623), .I1(n59655), .I2(n1625), .I3(n1628), 
            .O(n62396));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(n1624), .I1(n1622), .I2(n1626), .I3(n1627), 
            .O(n61049));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_18 (.CI(n51756), 
            .I0(GND_net), .I1(n17_adj_5899), .CO(n51757));
    SB_LUT4 encoder0_position_30__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n51124), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5900), .I3(n51755), .O(n18_adj_5740)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_19 (.CI(n51288), .I0(n2_adj_5884), .I1(n1653), .CO(n51289));
    SB_LUT4 add_2507_18_lut (.I0(n69661), .I1(n2_adj_5884), .I2(n1752), 
            .I3(n51287), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1838_21 (.CI(n51124), .I0(n2715), 
            .I1(VCC_net), .CO(n51125));
    SB_CARRY add_2507_18 (.CI(n51287), .I0(n2_adj_5884), .I1(n1752), .CO(n51288));
    SB_LUT4 encoder0_position_30__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n51123), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54169_4_lut (.I0(n61049), .I1(n1620), .I2(n1621), .I3(n62396), 
            .O(n1653));
    defparam i54169_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_2507_17_lut (.I0(n69555), .I1(n2_adj_5884), .I2(n1851), 
            .I3(n51286), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_17 (.CI(n51286), .I0(n2_adj_5884), .I1(n1851), .CO(n51287));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_17 (.CI(n51755), 
            .I0(GND_net), .I1(n18_adj_5900), .CO(n51756));
    SB_LUT4 add_2507_16_lut (.I0(n69371), .I1(n2_adj_5884), .I2(n1950), 
            .I3(n51285), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n50560), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_20 (.CI(n51123), .I0(n2716), 
            .I1(VCC_net), .CO(n51124));
    SB_LUT4 n11573_bdd_4_lut_54573 (.I0(n11573), .I1(current[2]), .I2(duty[5]), 
            .I3(n11571), .O(n70333));
    defparam n11573_bdd_4_lut_54573.LUT_INIT = 16'he4aa;
    SB_CARRY add_2507_16 (.CI(n51285), .I0(n2_adj_5884), .I1(n1950), .CO(n51286));
    SB_LUT4 add_2507_15_lut (.I0(n69821), .I1(n2_adj_5884), .I2(n2049), 
            .I3(n51284), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n51122), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5901), .I3(n51754), .O(n19_adj_5739)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n50559), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_15 (.CI(n51284), .I0(n2_adj_5884), .I1(n2049), .CO(n51285));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_16 (.CI(n51754), 
            .I0(GND_net), .I1(n19_adj_5901), .CO(n51755));
    SB_LUT4 add_2507_14_lut (.I0(n69845), .I1(n2_adj_5884), .I2(n2148), 
            .I3(n51283), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_14 (.CI(n51283), .I0(n2_adj_5884), .I1(n2148), .CO(n51284));
    SB_CARRY unary_minus_16_add_3_14 (.CI(n50559), .I0(GND_net), .I1(n2), 
            .CO(n50560));
    SB_CARRY encoder0_position_30__I_0_add_1838_19 (.CI(n51122), .I0(n2717), 
            .I1(VCC_net), .CO(n51123));
    SB_LUT4 add_2507_13_lut (.I0(n69870), .I1(n2_adj_5884), .I2(n2247), 
            .I3(n51282), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n50558), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_13 (.CI(n51282), .I0(n2_adj_5884), .I1(n2247), .CO(n51283));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n50558), .I0(GND_net), .I1(n14), 
            .CO(n50559));
    SB_LUT4 add_2507_12_lut (.I0(n69534), .I1(n2_adj_5884), .I2(n2346), 
            .I3(n51281), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_12 (.CI(n51281), .I0(n2_adj_5884), .I1(n2346), .CO(n51282));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5711), 
            .I3(n50557), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n50557), .I0(GND_net), .I1(n15_adj_5711), 
            .CO(n50558));
    SB_LUT4 encoder0_position_30__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n51121), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_11_lut (.I0(n69704), .I1(n2_adj_5884), .I2(n2445), 
            .I3(n51280), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1838_18 (.CI(n51121), .I0(n2718), 
            .I1(VCC_net), .CO(n51122));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5712), 
            .I3(n50556), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n50556), .I0(GND_net), .I1(n16_adj_5712), 
            .CO(n50557));
    SB_LUT4 encoder0_position_30__I_0_add_1168_17_lut (.I0(n69661), .I1(n1719), 
            .I2(VCC_net), .I3(n50715), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2507_11 (.CI(n51280), .I0(n2_adj_5884), .I1(n2445), .CO(n51281));
    SB_LUT4 encoder0_position_30__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n50714), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_10_lut (.I0(n69797), .I1(n2_adj_5884), .I2(n2544), 
            .I3(n51279), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1168_16 (.CI(n50714), .I0(n1720), 
            .I1(VCC_net), .CO(n50715));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5713), 
            .I3(n50555), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_5 (.CI(n50294), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n50295));
    SB_LUT4 encoder0_position_30__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n50713), .O(n1788_adj_5847)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n50555), .I0(GND_net), .I1(n17_adj_5713), 
            .CO(n50556));
    SB_CARRY encoder0_position_30__I_0_add_1168_15 (.CI(n50713), .I0(n1721), 
            .I1(VCC_net), .CO(n50714));
    SB_LUT4 encoder0_position_30__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n50712), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_10 (.CI(n51279), .I0(n2_adj_5884), .I1(n2544), .CO(n51280));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n50554), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_12 (.CI(n50301), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n50302));
    SB_LUT4 i28132_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n22773), .I3(GND_net), .O(n29423));
    defparam i28132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15569_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n58929), 
            .I3(GND_net), .O(n29600));   // verilog/coms.v(130[12] 305[6])
    defparam i15569_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1168_14 (.CI(n50712), .I0(n1722), 
            .I1(VCC_net), .CO(n50713));
    SB_LUT4 encoder0_position_30__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n51120), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n50554), .I0(GND_net), .I1(n18), 
            .CO(n50555));
    SB_LUT4 encoder0_position_30__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n50711), .O(n1790_adj_5848)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_13 (.CI(n50711), .I0(n1723), 
            .I1(VCC_net), .CO(n50712));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5714), 
            .I3(n50553), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n50553), .I0(GND_net), .I1(n19_adj_5714), 
            .CO(n50554));
    SB_LUT4 encoder0_position_30__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1852 (.I0(n1728), .I1(n1726), .I2(n1727), .I3(GND_net), 
            .O(n62302));
    defparam i1_3_lut_adj_1852.LUT_INIT = 16'hfefe;
    SB_LUT4 i29092_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n43019));
    defparam i29092_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n50710), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_17 (.CI(n51120), .I0(n2719), 
            .I1(VCC_net), .CO(n51121));
    SB_LUT4 add_2507_9_lut (.I0(n69766), .I1(n2_adj_5884), .I2(n2643), 
            .I3(n51278), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_151_32 (.CI(n50321), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n50322));
    SB_CARRY encoder0_position_30__I_0_add_1168_12 (.CI(n50710), .I0(n1724), 
            .I1(VCC_net), .CO(n50711));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n50320), .O(n1210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n50320), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n50321));
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n1723), .I1(n1724), .I2(n62302), .I3(n1725), 
            .O(n62308));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1854 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n62402));
    defparam i1_2_lut_adj_1854.LUT_INIT = 16'h8888;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n50709), .O(n1792_adj_5849)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5814));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15561_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n58929), 
            .I3(GND_net), .O(n29592));   // verilog/coms.v(130[12] 305[6])
    defparam i15561_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2507_9 (.CI(n51278), .I0(n2_adj_5884), .I1(n2643), .CO(n51279));
    SB_LUT4 add_2507_8_lut (.I0(n69734), .I1(n2_adj_5884), .I2(n2742), 
            .I3(n51277), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_8 (.CI(n51277), .I0(n2_adj_5884), .I1(n2742), .CO(n51278));
    SB_LUT4 encoder0_position_30__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n51119), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_16 (.CI(n51119), .I0(n2720), 
            .I1(VCC_net), .CO(n51120));
    SB_LUT4 encoder0_position_30__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n51118), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_11 (.CI(n50709), .I0(n1725), 
            .I1(VCC_net), .CO(n50710));
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n50300), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1587_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n12146));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5815));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1855 (.I0(n62402), .I1(n1722), .I2(n62308), .I3(n43019), 
            .O(n62312));
    defparam i1_4_lut_adj_1855.LUT_INIT = 16'hfefc;
    SB_LUT4 encoder0_position_30__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n50708), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_7_lut (.I0(n69654), .I1(n2_adj_5884), .I2(n2841), 
            .I3(n51276), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_7 (.CI(n51276), .I0(n2_adj_5884), .I1(n2841), .CO(n51277));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5902), .I3(n51753), .O(n20_adj_5738)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_10 (.CI(n50708), .I0(n1726), 
            .I1(VCC_net), .CO(n50709));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_15 (.CI(n51753), 
            .I0(GND_net), .I1(n20_adj_5902), .CO(n51754));
    SB_LUT4 add_2507_6_lut (.I0(n69587), .I1(n2_adj_5884), .I2(n2940), 
            .I3(n51275), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n50707), .O(n1794_adj_5850)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5903), .I3(n51752), .O(n21_adj_5737)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_6 (.CI(n51275), .I0(n2_adj_5884), .I1(n2940), .CO(n51276));
    SB_CARRY encoder0_position_30__I_0_add_1168_9 (.CI(n50707), .I0(n1727), 
            .I1(VCC_net), .CO(n50708));
    SB_LUT4 i53954_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n62312), 
            .O(n1752));
    defparam i53954_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_14 (.CI(n51752), 
            .I0(GND_net), .I1(n21_adj_5903), .CO(n51753));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5904), .I3(n51751), .O(n22_adj_5736)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_13 (.CI(n51751), 
            .I0(GND_net), .I1(n22_adj_5904), .CO(n51752));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5905), .I3(n51750), .O(n23_adj_5735)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_12 (.CI(n51750), 
            .I0(GND_net), .I1(n23_adj_5905), .CO(n51751));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20), 
            .I3(n50552), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_15 (.CI(n51118), .I0(n2721), 
            .I1(VCC_net), .CO(n51119));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5906), .I3(n51749), .O(n24_adj_5734)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n50706), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n50552), .I0(GND_net), .I1(n20), 
            .CO(n50553));
    SB_LUT4 mux_1587_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n12144));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i18_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(n17_adj_5868));
    defparam i18_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_11 (.CI(n51749), 
            .I0(GND_net), .I1(n24_adj_5906), .CO(n51750));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5907), .I3(n51748), .O(n25_adj_5733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_8 (.CI(n50706), .I0(n1728), 
            .I1(VCC_net), .CO(n50707));
    SB_LUT4 encoder0_position_30__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n50705), .O(n1796_adj_5851)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_5_lut (.I0(n69620), .I1(n2_adj_5884), .I2(n3039), 
            .I3(n51274), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_10 (.CI(n51748), 
            .I0(GND_net), .I1(n25_adj_5907), .CO(n51749));
    SB_CARRY add_2507_5 (.CI(n51274), .I0(n2_adj_5884), .I1(n3039), .CO(n51275));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21), 
            .I3(n50551), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n50551), .I0(GND_net), .I1(n21), 
            .CO(n50552));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n50319), .O(n1211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n51117), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5908), .I3(n51747), .O(n26_adj_5732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_4_lut (.I0(n69501), .I1(n2_adj_5884), .I2(n3138), 
            .I3(n51273), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_9 (.CI(n51747), 
            .I0(GND_net), .I1(n26_adj_5908), .CO(n51748));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5909), .I3(n51746), .O(n27_adj_5731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_8 (.CI(n51746), 
            .I0(GND_net), .I1(n27_adj_5909), .CO(n51747));
    SB_CARRY add_2507_4 (.CI(n51273), .I0(n2_adj_5884), .I1(n3138), .CO(n51274));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22), 
            .I3(n50550), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n50550), .I0(GND_net), .I1(n22), 
            .CO(n50551));
    SB_CARRY add_151_30 (.CI(n50319), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n50320));
    SB_CARRY encoder0_position_30__I_0_add_1838_14 (.CI(n51117), .I0(n2722), 
            .I1(VCC_net), .CO(n51118));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5910), .I3(n51745), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2507_3_lut (.I0(n69461), .I1(n2_adj_5884), .I2(n3237), 
            .I3(n51272), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2507_3 (.CI(n51272), .I0(n2_adj_5884), .I1(n3237), .CO(n51273));
    SB_CARRY encoder0_position_30__I_0_add_1168_7 (.CI(n50705), .I0(n1729), 
            .I1(GND_net), .CO(n50706));
    SB_LUT4 i15553_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n58929), 
            .I3(GND_net), .O(n29584));   // verilog/coms.v(130[12] 305[6])
    defparam i15553_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n50293), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n50318), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_7 (.CI(n51745), 
            .I0(GND_net), .I1(n28_adj_5910), .CO(n51746));
    SB_LUT4 add_2507_2_lut (.I0(n69467), .I1(n2_adj_5884), .I2(n43071), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2507_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n51116), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n50704), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23), 
            .I3(n50549), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_6 (.CI(n50704), .I0(n1730), 
            .I1(GND_net), .CO(n50705));
    SB_CARRY add_151_11 (.CI(n50300), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n50301));
    SB_LUT4 encoder0_position_30__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n50703), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5911), .I3(n51744), .O(n29_adj_5730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2507_2 (.CI(VCC_net), .I0(n2_adj_5884), .I1(n43071), 
            .CO(n51272));
    SB_CARRY unary_minus_16_add_3_4 (.CI(n50549), .I0(GND_net), .I1(n23), 
            .CO(n50550));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n50548), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_5 (.CI(n50703), .I0(n1731), 
            .I1(VCC_net), .CO(n50704));
    SB_CARRY unary_minus_16_add_3_3 (.CI(n50548), .I0(GND_net), .I1(n24), 
            .CO(n50549));
    SB_LUT4 i15550_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n58929), 
            .I3(GND_net), .O(n29581));   // verilog/coms.v(130[12] 305[6])
    defparam i15550_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15547_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n58929), 
            .I3(GND_net), .O(n29578));   // verilog/coms.v(130[12] 305[6])
    defparam i15547_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_33_lut (.I0(GND_net), .I1(n3204), 
            .I2(VCC_net), .I3(n51271), .O(n3271)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n50702), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_4 (.CI(n50702), .I0(n1732), 
            .I1(GND_net), .CO(n50703));
    SB_LUT4 encoder0_position_30__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n50701), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n51270), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_32 (.CI(n51270), .I0(n3205), 
            .I1(VCC_net), .CO(n51271));
    SB_LUT4 encoder0_position_30__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n51269), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15544_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n58929), 
            .I3(GND_net), .O(n29575));   // verilog/coms.v(130[12] 305[6])
    defparam i15544_3_lut.LUT_INIT = 16'hacac;
    SB_DFF read_197 (.Q(state_7__N_3919[0]), .C(clk16MHz), .D(n61190));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_CARRY encoder0_position_30__I_0_add_1168_3 (.CI(n50701), .I0(n1733), 
            .I1(VCC_net), .CO(n50702));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n42880), .I1(GND_net), .I2(n25), 
            .I3(VCC_net), .O(n66280)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_31 (.CI(n51269), .I0(n3206), 
            .I1(VCC_net), .CO(n51270));
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n50548));
    SB_CARRY add_151_29 (.CI(n50318), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n50319));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5805), .I3(n50547), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5804), .I3(n50546), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n51268), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_13 (.CI(n51116), .I0(n2723), 
            .I1(VCC_net), .CO(n51117));
    SB_LUT4 encoder0_position_30__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n50317), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_6 (.CI(n51744), 
            .I0(GND_net), .I1(n29_adj_5911), .CO(n51745));
    SB_CARRY encoder0_position_30__I_0_add_2173_30 (.CI(n51268), .I0(n3207), 
            .I1(VCC_net), .CO(n51269));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n50546), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5804), .CO(n50547));
    SB_LUT4 encoder0_position_30__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n50701));
    SB_LUT4 encoder0_position_30__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n51267), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5803), .I3(n50545), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n51115), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_151_28 (.CI(n50317), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n50318));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5912), .I3(n51743), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_12 (.CI(n51115), .I0(n2724), 
            .I1(VCC_net), .CO(n51116));
    SB_LUT4 encoder0_position_30__I_0_add_1570_23_lut (.I0(n69534), .I1(n2313), 
            .I2(VCC_net), .I3(n50937), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_5 (.CI(n51743), 
            .I0(GND_net), .I1(n30_adj_5912), .CO(n51744));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5913), .I3(n51742), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27735), 
            .D(n1229), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_4 (.CI(n51742), 
            .I0(GND_net), .I1(n31_adj_5913), .CO(n51743));
    SB_CARRY encoder0_position_30__I_0_add_2173_29 (.CI(n51267), .I0(n3208), 
            .I1(VCC_net), .CO(n51268));
    SB_LUT4 encoder0_position_30__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n51266), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n70333_bdd_4_lut (.I0(n70333), .I1(duty[2]), .I2(n4928), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n70333_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5914), .I3(n51741), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_3 (.CI(n51741), 
            .I0(GND_net), .I1(n32_adj_5914), .CO(n51742));
    SB_CARRY encoder0_position_30__I_0_add_2173_28 (.CI(n51266), .I0(n3209), 
            .I1(VCC_net), .CO(n51267));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n50545), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5803), .CO(n50546));
    SB_LUT4 encoder0_position_30__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n51265), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_27 (.CI(n51265), .I0(n3210), 
            .I1(VCC_net), .CO(n51266));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n51741));
    SB_LUT4 encoder0_position_30__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n51114), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n51264), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1856 (.I0(n1826), .I1(n1827), .I2(n1825), .I3(n1828), 
            .O(n62428));
    defparam i1_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 n11573_bdd_4_lut_54568 (.I0(n11573), .I1(current[1]), .I2(duty[4]), 
            .I3(n11571), .O(n70327));
    defparam n11573_bdd_4_lut_54568.LUT_INIT = 16'he4aa;
    SB_LUT4 n70327_bdd_4_lut (.I0(n70327), .I1(duty[1]), .I2(n4929), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n70327_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15860_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n58897), 
            .I3(GND_net), .O(n29891));   // verilog/coms.v(130[12] 305[6])
    defparam i15860_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_11 (.CI(n51114), .I0(n2725), 
            .I1(VCC_net), .CO(n51115));
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n50936), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48176_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63902));
    defparam i48176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48177_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63903));
    defparam i48177_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2173_26 (.CI(n51264), .I0(n3211), 
            .I1(VCC_net), .CO(n51265));
    SB_LUT4 encoder0_position_30__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n51263), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n50316), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n51113), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_25 (.CI(n51263), .I0(n3212), 
            .I1(VCC_net), .CO(n51264));
    SB_CARRY encoder0_position_30__I_0_add_1570_22 (.CI(n50936), .I0(n2314), 
            .I1(VCC_net), .CO(n50937));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5833), .I3(n50544), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n51262), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48174_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63900));
    defparam i48174_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2173_24 (.CI(n51262), .I0(n3213), 
            .I1(VCC_net), .CO(n51263));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n50544), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5833), .CO(n50545));
    SB_LUT4 i48173_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63899));
    defparam i48173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5830), .I3(n50543), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29102_4_lut (.I0(n943), .I1(n1831), .I2(n1832), .I3(n1833), 
            .O(n43029));
    defparam i29102_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n51261), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_23 (.CI(n51261), .I0(n3214), 
            .I1(VCC_net), .CO(n51262));
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n1822_adj_5852), .I1(n1823), .I2(n1824_adj_5853), 
            .I3(n62428), .O(n62434));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1858 (.I0(n1829), .I1(n1830), .I2(GND_net), .I3(GND_net), 
            .O(n62536));
    defparam i1_2_lut_adj_1858.LUT_INIT = 16'h8888;
    SB_LUT4 n11573_bdd_4_lut_54563 (.I0(n11573), .I1(current[0]), .I2(duty[3]), 
            .I3(n11571), .O(n70321));
    defparam n11573_bdd_4_lut_54563.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(n1821), .I1(n62536), .I2(n62434), .I3(n43029), 
            .O(n62438));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_30__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n51260), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n50935), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_21 (.CI(n50935), .I0(n2315), 
            .I1(VCC_net), .CO(n50936));
    SB_LUT4 i53832_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n62438), 
            .O(n1851));
    defparam i53832_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1172_3_lut (.I0(n1721), .I1(n1788_adj_5847), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n50934), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_22 (.CI(n51260), .I0(n3215), 
            .I1(VCC_net), .CO(n51261));
    SB_LUT4 LessThan_1089_i15_2_lut (.I0(r_Clock_Count_adj_6024[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5880));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1089_i9_2_lut (.I0(r_Clock_Count_adj_6024[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5877));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_151_27 (.CI(n50316), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n50317));
    SB_LUT4 LessThan_1089_i13_2_lut (.I0(r_Clock_Count_adj_6024[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5879));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1089_i11_2_lut (.I0(r_Clock_Count_adj_6024[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5878));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n50543), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5830), .CO(n50544));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5829), .I3(n50542), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n50542), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5829), .CO(n50543));
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n50315), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n51259), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_1089_i4_4_lut (.I0(r_Clock_Count_adj_6024[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_6024[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5874));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52891_3_lut (.I0(n4_adj_5874), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5878), 
            .I3(GND_net), .O(n68617));   // verilog/uart_tx.v(117[17:57])
    defparam i52891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52892_3_lut (.I0(n68617), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5879), 
            .I3(GND_net), .O(n68618));   // verilog/uart_tx.v(117[17:57])
    defparam i52892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52330_4_lut (.I0(n13_adj_5879), .I1(n11_adj_5878), .I2(n9_adj_5877), 
            .I3(n67204), .O(n68056));
    defparam i52330_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1089_i8_3_lut (.I0(n6_adj_5875), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5877), .I3(GND_net), .O(n8_adj_5876));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51961_3_lut (.I0(n68618), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5880), 
            .I3(GND_net), .O(n67687));   // verilog/uart_tx.v(117[17:57])
    defparam i51961_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27735), 
            .D(n1228), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27735), 
            .D(n1227), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i52893_4_lut (.I0(n67687), .I1(n8_adj_5876), .I2(n15_adj_5880), 
            .I3(n68056), .O(n68619));   // verilog/uart_tx.v(117[17:57])
    defparam i52893_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY encoder0_position_30__I_0_add_2173_21 (.CI(n51259), .I0(n3216), 
            .I1(VCC_net), .CO(n51260));
    SB_LUT4 i52894_3_lut (.I0(n68619), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_6024[8]), 
            .I3(GND_net), .O(n4942));   // verilog/uart_tx.v(117[17:57])
    defparam i52894_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1860 (.I0(n23_adj_5728), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n4942), .I3(GND_net), .O(n61392));
    defparam i1_3_lut_adj_1860.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n61392), .O(r_SM_Main_2__N_3536[1]));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1838_10 (.CI(n51113), .I0(n2726), 
            .I1(VCC_net), .CO(n51114));
    SB_CARRY encoder0_position_30__I_0_add_1570_20 (.CI(n50934), .I0(n2316), 
            .I1(VCC_net), .CO(n50935));
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27735), 
            .D(n1226), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27735), 
            .D(n1225), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27735), 
            .D(n1224), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27735), 
            .D(n1223), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27735), 
            .D(n1222), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27735), 
            .D(n1221), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27735), 
            .D(n1220), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27735), 
            .D(n1219), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27735), 
            .D(n1218), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27735), 
            .D(n1217), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27735), 
            .D(n1216), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27735), 
            .D(n1215), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27735), 
            .D(n1214), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27735), 
            .D(n1213), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27735), 
            .D(n1212), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27735), 
            .D(n1211), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27735), 
            .D(n1210), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27735), 
            .D(n1209), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27735), 
            .D(n1208), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR dti_counter_1938__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n27779), 
            .D(n44), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1938__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n27779), 
            .D(n43), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1938__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n27779), 
            .D(n42), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1938__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n27779), 
            .D(n41_adj_5881), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1938__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n27779), 
            .D(n40), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1938__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n27779), 
            .D(n39), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1938__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n27779), 
            .D(n38), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n50933), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n51258), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_20 (.CI(n51258), .I0(n3217), 
            .I1(VCC_net), .CO(n51259));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5828), .I3(n50541), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15782_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n58010), 
            .I3(GND_net), .O(n29813));   // verilog/coms.v(130[12] 305[6])
    defparam i15782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n51257), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_19 (.CI(n50933), .I0(n2317), 
            .I1(VCC_net), .CO(n50934));
    SB_CARRY encoder0_position_30__I_0_add_2173_19 (.CI(n51257), .I0(n3218), 
            .I1(VCC_net), .CO(n51258));
    SB_CARRY add_151_26 (.CI(n50315), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n50316));
    SB_LUT4 encoder0_position_30__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n51256), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n51112), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_18 (.CI(n51256), .I0(n3219), 
            .I1(VCC_net), .CO(n51257));
    SB_LUT4 i15626_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n58009), 
            .I3(GND_net), .O(n29657));   // verilog/coms.v(130[12] 305[6])
    defparam i15626_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_9 (.CI(n51112), .I0(n2727), 
            .I1(VCC_net), .CO(n51113));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n50541), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5828), .CO(n50542));
    SB_LUT4 encoder0_position_30__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n51111), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15610_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n58009), 
            .I3(GND_net), .O(n29641));   // verilog/coms.v(130[12] 305[6])
    defparam i15610_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n50932), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1086_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5873));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1086_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1086_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5870));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1086_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_1086_i8_3_lut (.I0(n6_adj_5871), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5873), .I3(GND_net), .O(n8_adj_5872));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1086_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53318_4_lut (.I0(n8_adj_5872), .I1(n4_adj_5870), .I2(n9_adj_5873), 
            .I3(n67210), .O(n69044));   // verilog/uart_rx.v(119[17:57])
    defparam i53318_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53319_3_lut (.I0(n69044), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n69045));   // verilog/uart_rx.v(119[17:57])
    defparam i53319_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n51255), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_18 (.CI(n50932), .I0(n2318), 
            .I1(VCC_net), .CO(n50933));
    SB_CARRY encoder0_position_30__I_0_add_2173_17 (.CI(n51255), .I0(n3220), 
            .I1(VCC_net), .CO(n51256));
    SB_LUT4 i53186_3_lut (.I0(n69045), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n68912));   // verilog/uart_rx.v(119[17:57])
    defparam i53186_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51959_3_lut (.I0(n68912), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4939));   // verilog/uart_rx.v(119[17:57])
    defparam i51959_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n23_adj_5728), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n4939), .I3(o_Rx_DV_N_3488[8]), .O(n61336));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n61336), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1838_8 (.CI(n51111), .I0(n2728), 
            .I1(VCC_net), .CO(n51112));
    SB_LUT4 encoder0_position_30__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n51254), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_16 (.CI(n51254), .I0(n3221), 
            .I1(VCC_net), .CO(n51255));
    SB_LUT4 encoder0_position_30__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n51110), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dti_counter_1938__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n27779), 
            .D(n45), .R(n29059));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_add_1101_16_lut (.I0(n69892), .I1(n1620), 
            .I2(VCC_net), .I3(n50688), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n51253), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n50931), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_15 (.CI(n51253), .I0(n3222), 
            .I1(VCC_net), .CO(n51254));
    SB_LUT4 i15787_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n58010), 
            .I3(GND_net), .O(n29818));   // verilog/coms.v(130[12] 305[6])
    defparam i15787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut (.I0(ID[0]), .I1(ID[6]), .I2(ID[2]), .I3(ID[4]), 
            .O(n61122));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(ID[5]), .I1(n61122), .I2(ID[3]), .I3(GND_net), 
            .O(n8_adj_5860));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_adj_1864 (.I0(ID[1]), .I1(ID[7]), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_5861));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i2_2_lut_adj_1864.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n51252), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28248_4_lut (.I0(n7_adj_5861), .I1(baudrate[0]), .I2(n8_adj_5860), 
            .I3(n25566), .O(n42168));
    defparam i28248_4_lut.LUT_INIT = 16'hc8fa;
    SB_CARRY encoder0_position_30__I_0_add_2173_14 (.CI(n51252), .I0(n3223), 
            .I1(VCC_net), .CO(n51253));
    SB_LUT4 encoder0_position_30__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n51251), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_17 (.CI(n50931), .I0(n2319), 
            .I1(VCC_net), .CO(n50932));
    SB_LUT4 i1_2_lut_adj_1865 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5933));
    defparam i1_2_lut_adj_1865.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_5933), .I2(delay_counter[10]), 
            .I3(n25452), .O(n59833));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1866 (.I0(n59833), .I1(n25457), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n60784));
    defparam i2_4_lut_adj_1866.LUT_INIT = 16'hffec;
    SB_LUT4 encoder0_position_30__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n50930), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n50687), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_13 (.CI(n51251), .I0(n3224), 
            .I1(VCC_net), .CO(n51252));
    SB_CARRY encoder0_position_30__I_0_add_1838_7 (.CI(n51110), .I0(n2729), 
            .I1(GND_net), .CO(n51111));
    SB_LUT4 encoder0_position_30__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n51109), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_3_lut_adj_1867 (.I0(delay_counter[20]), .I1(delay_counter[21]), 
            .I2(delay_counter[23]), .I3(GND_net), .O(n8));
    defparam i3_3_lut_adj_1867.LUT_INIT = 16'h8080;
    SB_CARRY encoder0_position_30__I_0_add_1570_16 (.CI(n50930), .I0(n2320), 
            .I1(VCC_net), .CO(n50931));
    SB_CARRY encoder0_position_30__I_0_add_1101_15 (.CI(n50687), .I0(n1621), 
            .I1(VCC_net), .CO(n50688));
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n56399));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n50929), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n50686), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_14 (.CI(n50686), .I0(n1622), 
            .I1(VCC_net), .CO(n50687));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5827), .I3(n50540), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n50685), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30425));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n51250), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_12 (.CI(n51250), .I0(n3225), 
            .I1(VCC_net), .CO(n51251));
    SB_CARRY encoder0_position_30__I_0_add_1570_15 (.CI(n50929), .I0(n2321), 
            .I1(VCC_net), .CO(n50930));
    SB_LUT4 i2_4_lut_adj_1868 (.I0(delay_counter[22]), .I1(n60784), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7));
    defparam i2_4_lut_adj_1868.LUT_INIT = 16'ha8a0;
    SB_CARRY encoder0_position_30__I_0_add_1101_13 (.CI(n50685), .I0(n1623), 
            .I1(VCC_net), .CO(n50686));
    SB_LUT4 encoder0_position_30__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n50684), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n50540), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5827), .CO(n50541));
    SB_LUT4 encoder0_position_30__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n51249), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_11 (.CI(n51249), .I0(n3226), 
            .I1(VCC_net), .CO(n51250));
    SB_CARRY encoder0_position_30__I_0_add_1838_6 (.CI(n51109), .I0(n2730), 
            .I1(GND_net), .CO(n51110));
    SB_CARRY encoder0_position_30__I_0_add_1101_12 (.CI(n50684), .I0(n1624), 
            .I1(VCC_net), .CO(n50685));
    SB_LUT4 encoder0_position_30__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n50683), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n70321_bdd_4_lut (.I0(n70321), .I1(duty[0]), .I2(n4930), .I3(n11571), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n70321_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n50928), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5826), .I3(n50539), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n51248), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_10 (.CI(n51248), .I0(n3227), 
            .I1(VCC_net), .CO(n51249));
    SB_CARRY encoder0_position_30__I_0_add_1101_11 (.CI(n50683), .I0(n1625), 
            .I1(VCC_net), .CO(n50684));
    SB_LUT4 i28451_4_lut (.I0(n7), .I1(delay_counter[31]), .I2(n25460), 
            .I3(n8), .O(n1319));   // verilog/TinyFPGA_B.v(380[14:38])
    defparam i28451_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_3_lut (.I0(delay_counter[17]), .I1(delay_counter[16]), .I2(delay_counter[15]), 
            .I3(GND_net), .O(n25457));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5769));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1869 (.I0(delay_counter[28]), .I1(n12_adj_5769), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n25460));
    defparam i6_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n50539), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5826), .CO(n50540));
    SB_CARRY encoder0_position_30__I_0_add_1570_14 (.CI(n50928), .I0(n2322), 
            .I1(VCC_net), .CO(n50929));
    SB_LUT4 encoder0_position_30__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n51247), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_3_lut_adj_1870 (.I0(delay_counter[0]), .I1(delay_counter[4]), 
            .I2(delay_counter[8]), .I3(GND_net), .O(n8_adj_5786));
    defparam i3_3_lut_adj_1870.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n50682), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1871 (.I0(delay_counter[5]), .I1(delay_counter[6]), 
            .I2(delay_counter[1]), .I3(delay_counter[2]), .O(n60799));
    defparam i3_4_lut_adj_1871.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1872 (.I0(n60799), .I1(delay_counter[7]), .I2(n8_adj_5786), 
            .I3(delay_counter[3]), .O(n25452));
    defparam i8_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n50927), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4888_4_lut (.I0(n25452), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5859));
    defparam i4888_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1873 (.I0(n24_adj_5859), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n60713));
    defparam i2_4_lut_adj_1873.LUT_INIT = 16'hc800;
    SB_LUT4 i1_4_lut_adj_1874 (.I0(delay_counter[22]), .I1(delay_counter[21]), 
            .I2(n25460), .I3(delay_counter[23]), .O(n4_adj_5931));
    defparam i1_4_lut_adj_1874.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1101_10 (.CI(n50682), .I0(n1626), 
            .I1(VCC_net), .CO(n50683));
    SB_LUT4 encoder0_position_30__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n50681), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5825), .I3(n50538), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_9 (.CI(n51247), .I0(n3228), 
            .I1(VCC_net), .CO(n51248));
    SB_LUT4 encoder0_position_30__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n51246), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_9 (.CI(n50681), .I0(n1627), 
            .I1(VCC_net), .CO(n50682));
    SB_LUT4 encoder0_position_30__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n51108), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_8 (.CI(n51246), .I0(n3229), 
            .I1(GND_net), .CO(n51247));
    SB_LUT4 encoder0_position_30__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n51245), .O(n66396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1838_5 (.CI(n51108), .I0(n2731), 
            .I1(VCC_net), .CO(n51109));
    SB_CARRY encoder0_position_30__I_0_add_1570_13 (.CI(n50927), .I0(n2323), 
            .I1(VCC_net), .CO(n50928));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n50538), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5825), .CO(n50539));
    SB_LUT4 encoder0_position_30__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n50926), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_7 (.CI(n51245), .I0(n3230), 
            .I1(GND_net), .CO(n51246));
    SB_LUT4 encoder0_position_30__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n50680), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n51107), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1875 (.I0(n60713), .I1(delay_counter[18]), .I2(n25457), 
            .I3(GND_net), .O(n61098));
    defparam i2_3_lut_adj_1875.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1876 (.I0(n61098), .I1(n4_adj_5931), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n62));
    defparam i2_4_lut_adj_1876.LUT_INIT = 16'heccc;
    SB_LUT4 i28450_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(366[12:35])
    defparam i28450_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY encoder0_position_30__I_0_add_1101_8 (.CI(n50680), .I0(n1628), 
            .I1(VCC_net), .CO(n50681));
    SB_LUT4 encoder0_position_30__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n50679), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_7 (.CI(n50679), .I0(n1629), 
            .I1(GND_net), .CO(n50680));
    SB_CARRY encoder0_position_30__I_0_add_1570_12 (.CI(n50926), .I0(n2324), 
            .I1(VCC_net), .CO(n50927));
    SB_LUT4 i586_2_lut (.I0(n1319), .I1(n42168), .I2(GND_net), .I3(GND_net), 
            .O(n2821));   // verilog/TinyFPGA_B.v(384[18] 386[12])
    defparam i586_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n50925), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n51244), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_4 (.CI(n51107), .I0(n2732), 
            .I1(GND_net), .CO(n51108));
    SB_CARRY encoder0_position_30__I_0_add_1570_11 (.CI(n50925), .I0(n2325), 
            .I1(VCC_net), .CO(n50926));
    SB_LUT4 encoder0_position_30__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n50924), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_10 (.CI(n50924), .I0(n2326), 
            .I1(VCC_net), .CO(n50925));
    SB_LUT4 encoder0_position_30__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n50678), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16521_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n30552));   // verilog/coms.v(130[12] 305[6])
    defparam i16521_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_2173_6 (.CI(n51244), .I0(n3231), 
            .I1(VCC_net), .CO(n51245));
    SB_LUT4 i47830_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n63547));
    defparam i47830_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54333_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6619), .I2(n63547), 
            .I3(n25_adj_5928), .O(n17_adj_5927));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i54333_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5816), .I3(n50537), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n51106), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_6 (.CI(n50678), .I0(n1630), 
            .I1(GND_net), .CO(n50679));
    SB_LUT4 encoder0_position_30__I_0_add_2173_5_lut (.I0(n6_adj_5749), .I1(n3232), 
            .I2(GND_net), .I3(n51243), .O(n66389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_5_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 encoder0_position_30__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n50923), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_3 (.CI(n51106), .I0(n2733), 
            .I1(VCC_net), .CO(n51107));
    SB_CARRY encoder0_position_30__I_0_add_1570_9 (.CI(n50923), .I0(n2327), 
            .I1(VCC_net), .CO(n50924));
    SB_CARRY encoder0_position_30__I_0_add_2173_5 (.CI(n51243), .I0(n3232), 
            .I1(GND_net), .CO(n51244));
    SB_LUT4 encoder0_position_30__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n50922), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_8 (.CI(n50922), .I0(n2328), 
            .I1(VCC_net), .CO(n50923));
    SB_LUT4 encoder0_position_30__I_0_add_2173_4_lut (.I0(n3301), .I1(n3233), 
            .I2(VCC_net), .I3(n51242), .O(n6_adj_5749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n51106));
    SB_CARRY encoder0_position_30__I_0_add_2173_4 (.CI(n51242), .I0(n3233), 
            .I1(VCC_net), .CO(n51243));
    SB_LUT4 encoder0_position_30__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n50677), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n50921), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_7 (.CI(n50921), .I0(n2329), 
            .I1(GND_net), .CO(n50922));
    SB_CARRY encoder0_position_30__I_0_add_1101_5 (.CI(n50677), .I0(n1631), 
            .I1(VCC_net), .CO(n50678));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n50537), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5816), .CO(n50538));
    SB_LUT4 encoder0_position_30__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n50676), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n50431), .O(n4907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_4 (.CI(n50676), .I0(n1632), 
            .I1(GND_net), .CO(n50677));
    SB_LUT4 encoder0_position_30__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n50920), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n51241), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_3 (.CI(n51241), .I0(n957), 
            .I1(GND_net), .CO(n51242));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n50314), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15535_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n7_adj_5939), 
            .I3(GND_net), .O(n29566));   // verilog/coms.v(130[12] 305[6])
    defparam i15535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n50675), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n51241));
    SB_CARRY encoder0_position_30__I_0_add_1101_3 (.CI(n50675), .I0(n1633), 
            .I1(VCC_net), .CO(n50676));
    SB_CARRY encoder0_position_30__I_0_add_1570_6 (.CI(n50920), .I0(n2330), 
            .I1(GND_net), .CO(n50921));
    SB_LUT4 encoder0_position_30__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n50919), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_5 (.CI(n50919), .I0(n2331), 
            .I1(VCC_net), .CO(n50920));
    SB_LUT4 add_1100_24_lut (.I0(GND_net), .I1(GND_net), .I2(n12144), 
            .I3(n50430), .O(n4908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n50918), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_31_lut (.I0(n69501), .I1(n3105), 
            .I2(VCC_net), .I3(n51240), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1570_4 (.CI(n50918), .I0(n2332), 
            .I1(GND_net), .CO(n50919));
    SB_LUT4 encoder0_position_30__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n50917), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n50675));
    SB_CARRY add_151_25 (.CI(n50314), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n50315));
    SB_CARRY add_1100_24 (.CI(n50430), .I0(GND_net), .I1(n12144), .CO(n50431));
    SB_LUT4 encoder0_position_30__I_0_add_1034_15_lut (.I0(n70025), .I1(n1521), 
            .I2(VCC_net), .I3(n50674), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5815), .I3(n50536), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n50536), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5815), .CO(n50537));
    SB_LUT4 add_1100_23_lut (.I0(GND_net), .I1(GND_net), .I2(n12146), 
            .I3(n50429), .O(n4909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n50673), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5816));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15529_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n7_adj_5939), 
            .I3(GND_net), .O(n29560));   // verilog/coms.v(130[12] 305[6])
    defparam i15529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1877 (.I0(n1927), .I1(n1926), .I2(n1925), .I3(n1928), 
            .O(n62244));
    defparam i1_4_lut_adj_1877.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5814), .I3(n50535), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_3 (.CI(n50917), .I0(n2333), 
            .I1(VCC_net), .CO(n50918));
    SB_LUT4 encoder0_position_30__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n51239), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n50917));
    SB_LUT4 mux_4306_i27_3_lut (.I0(encoder0_position[26]), .I1(n6_adj_5753), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_4306_i28_3_lut (.I0(encoder0_position[27]), .I1(n5_adj_5775), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n405_adj_5787));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29110_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n43037));
    defparam i29110_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15510_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n7_adj_5939), 
            .I3(GND_net), .O(n29541));   // verilog/coms.v(130[12] 305[6])
    defparam i15510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i29_3_lut (.I0(encoder0_position[28]), .I1(n4_adj_5776), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15507_3_lut (.I0(\data_in_frame[2] [0]), .I1(rx_data[0]), .I2(n7_adj_5939), 
            .I3(GND_net), .O(n29538));   // verilog/coms.v(130[12] 305[6])
    defparam i15507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1878 (.I0(n1922), .I1(n1923), .I2(n62244), .I3(n1924), 
            .O(n62250));
    defparam i1_4_lut_adj_1878.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_2106_30 (.CI(n51239), .I0(n3106), 
            .I1(VCC_net), .CO(n51240));
    SB_LUT4 i1_4_lut_adj_1879 (.I0(n1929), .I1(n43037), .I2(n1930), .I3(n1931), 
            .O(n59677));
    defparam i1_4_lut_adj_1879.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1880 (.I0(n1920), .I1(n59677), .I2(n1921), .I3(n62250), 
            .O(n62256));
    defparam i1_4_lut_adj_1880.LUT_INIT = 16'hfffe;
    SB_LUT4 i53648_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n62256), 
            .O(n1950));
    defparam i53648_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1881 (.I0(n2027), .I1(n2024), .I2(GND_net), .I3(GND_net), 
            .O(n62452));
    defparam i1_2_lut_adj_1881.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1882 (.I0(n2025), .I1(n62452), .I2(n2026), .I3(n2028), 
            .O(n62456));
    defparam i1_4_lut_adj_1882.LUT_INIT = 16'hfffe;
    SB_LUT4 i29108_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n43035));
    defparam i29108_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_4306_i30_3_lut (.I0(encoder0_position[29]), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5996_2_lut (.I0(n2_adj_5778), .I1(encoder0_position[30]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i5996_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15489_3_lut (.I0(\data_in_frame[22] [7]), .I1(rx_data[7]), 
            .I2(n28352), .I3(GND_net), .O(n29520));   // verilog/coms.v(130[12] 305[6])
    defparam i15489_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1883 (.I0(n2021), .I1(n2022), .I2(n62456), .I3(n2023), 
            .O(n62462));
    defparam i1_4_lut_adj_1883.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1884 (.I0(n2029), .I1(n43035), .I2(n2030), .I3(n2031), 
            .O(n59714));
    defparam i1_4_lut_adj_1884.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1885 (.I0(n2019), .I1(n2020), .I2(n59714), .I3(n62462), 
            .O(n62468));
    defparam i1_4_lut_adj_1885.LUT_INIT = 16'hfffe;
    SB_LUT4 i54098_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n62468), 
            .O(n2049));
    defparam i54098_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n51238), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_29 (.CI(n51238), .I0(n3107), 
            .I1(VCC_net), .CO(n51239));
    SB_LUT4 i1_3_lut_adj_1886 (.I0(n2125), .I1(n2124), .I2(n2128), .I3(GND_net), 
            .O(n62278));
    defparam i1_3_lut_adj_1886.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1887 (.I0(n2123), .I1(n2127), .I2(n2126), .I3(GND_net), 
            .O(n62280));
    defparam i1_3_lut_adj_1887.LUT_INIT = 16'hfefe;
    SB_LUT4 i29176_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n43103));
    defparam i29176_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1888 (.I0(n2121), .I1(n2122), .I2(n62280), .I3(n62278), 
            .O(n62286));
    defparam i1_4_lut_adj_1888.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n2129), .I1(n62286), .I2(n43103), .I3(n2130), 
            .O(n62288));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1890 (.I0(n2118), .I1(n2119), .I2(n62288), .I3(n2120), 
            .O(n62294));
    defparam i1_4_lut_adj_1890.LUT_INIT = 16'hfffe;
    SB_LUT4 i15794_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[1]), .I2(n5_adj_5812), 
            .I3(n25563), .O(n29825));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15794_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54122_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n62294), 
            .O(n2148));
    defparam i54122_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15795_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[2]), .I2(n5_adj_5789), 
            .I3(n25563), .O(n29826));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15795_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1891 (.I0(n2226), .I1(n2223), .I2(n2227), .I3(n2225), 
            .O(n62484));
    defparam i1_4_lut_adj_1891.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1892 (.I0(n62484), .I1(n2224), .I2(n2228), .I3(GND_net), 
            .O(n62486));
    defparam i1_3_lut_adj_1892.LUT_INIT = 16'hfefe;
    SB_LUT4 i15796_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[3]), .I2(n6_adj_5809), 
            .I3(n25555), .O(n29827));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15796_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15797_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[4]), .I2(n6_adj_5777), 
            .I3(n25544), .O(n29828));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15797_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15798_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[5]), .I2(n6_adj_5777), 
            .I3(n25579), .O(n29829));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15798_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29174_4_lut (.I0(n947), .I1(n2231), .I2(n2232), .I3(n2233), 
            .O(n43101));
    defparam i29174_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15799_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[6]), .I2(n6_adj_5777), 
            .I3(n25573), .O(n29830));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15799_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1893 (.I0(n2220), .I1(n2221), .I2(n62486), .I3(n2222), 
            .O(n62492));
    defparam i1_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 i15800_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[7]), .I2(n6_adj_5777), 
            .I3(n25555), .O(n29831));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15800_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15483_3_lut (.I0(\data_in_frame[22] [5]), .I1(rx_data[5]), 
            .I2(n28352), .I3(GND_net), .O(n29514));   // verilog/coms.v(130[12] 305[6])
    defparam i15483_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15801_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[8]), .I2(n6_adj_5774), 
            .I3(n25544), .O(n29832));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15801_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1894 (.I0(n2229), .I1(n62492), .I2(n43101), .I3(n2230), 
            .O(n62494));
    defparam i1_4_lut_adj_1894.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1895 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n62494), 
            .O(n62500));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 i15802_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[9]), .I2(n6_adj_5774), 
            .I3(n25579), .O(n29833));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15802_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_1086_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5871));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1086_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i54147_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n62500), 
            .O(n2247));
    defparam i54147_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51484_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n67210));   // verilog/uart_rx.v(119[17:57])
    defparam i51484_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i15803_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[10]), .I2(n6_adj_5774), 
            .I3(n25573), .O(n29834));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15803_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15804_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[11]), .I2(n6_adj_5774), 
            .I3(n25555), .O(n29835));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15804_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15480_3_lut (.I0(\data_in_frame[22] [4]), .I1(rx_data[4]), 
            .I2(n28352), .I3(GND_net), .O(n29511));   // verilog/coms.v(130[12] 305[6])
    defparam i15480_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n51237), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4306_i4_3_lut (.I0(encoder0_position[3]), .I1(n29_adj_5730), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15805_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[12]), .I2(n42331), 
            .I3(n25544), .O(n29836));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15805_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15477_3_lut (.I0(\data_in_frame[22] [3]), .I1(rx_data[3]), 
            .I2(n28352), .I3(GND_net), .O(n29508));   // verilog/coms.v(130[12] 305[6])
    defparam i15477_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2106_28 (.CI(n51237), .I0(n3108), 
            .I1(VCC_net), .CO(n51238));
    SB_LUT4 i15474_3_lut (.I0(\data_in_frame[22] [2]), .I1(rx_data[2]), 
            .I2(n28352), .I3(GND_net), .O(n29505));   // verilog/coms.v(130[12] 305[6])
    defparam i15474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51478_3_lut_4_lut (.I0(r_Clock_Count_adj_6024[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_6024[2]), .O(n67204));   // verilog/uart_tx.v(117[17:57])
    defparam i51478_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i15806_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[15]), .I2(n42331), 
            .I3(n25555), .O(n29837));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15806_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15807_3_lut (.I0(\data_in_frame[0] [1]), .I1(rx_data[1]), .I2(n58008), 
            .I3(GND_net), .O(n29838));   // verilog/coms.v(130[12] 305[6])
    defparam i15807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15810_3_lut (.I0(\data_in_frame[0] [2]), .I1(rx_data[2]), .I2(n58008), 
            .I3(GND_net), .O(n29841));   // verilog/coms.v(130[12] 305[6])
    defparam i15810_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1089_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_6024[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5875));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1089_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i15471_3_lut (.I0(\data_in_frame[22] [1]), .I1(rx_data[1]), 
            .I2(n28352), .I3(GND_net), .O(n29502));   // verilog/coms.v(130[12] 305[6])
    defparam i15471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n51236), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15813_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n58008), 
            .I3(GND_net), .O(n29844));   // verilog/coms.v(130[12] 305[6])
    defparam i15813_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2106_27 (.CI(n51236), .I0(n3109), 
            .I1(VCC_net), .CO(n51237));
    SB_LUT4 i15590_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n58009), 
            .I3(GND_net), .O(n29621));   // verilog/coms.v(130[12] 305[6])
    defparam i15590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15817_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n58010), 
            .I3(GND_net), .O(n29848));   // verilog/coms.v(130[12] 305[6])
    defparam i15817_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15820_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n58010), 
            .I3(GND_net), .O(n29851));   // verilog/coms.v(130[12] 305[6])
    defparam i15820_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15823_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n58010), 
            .I3(GND_net), .O(n29854));   // verilog/coms.v(130[12] 305[6])
    defparam i15823_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15826_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n58010), 
            .I3(GND_net), .O(n29857));   // verilog/coms.v(130[12] 305[6])
    defparam i15826_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15829_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n58011), 
            .I3(GND_net), .O(n29860));   // verilog/coms.v(130[12] 305[6])
    defparam i15829_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15832_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n58011), 
            .I3(GND_net), .O(n29863));   // verilog/coms.v(130[12] 305[6])
    defparam i15832_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15835_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n58011), 
            .I3(GND_net), .O(n29866));   // verilog/coms.v(130[12] 305[6])
    defparam i15835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50944_4_lut (.I0(bit_ctr[0]), .I1(n66110), .I2(n52805), .I3(color_bit_N_502[1]), 
            .O(n66446));   // verilog/neopixel.v(34[12] 116[6])
    defparam i50944_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i15838_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n58011), 
            .I3(GND_net), .O(n29869));   // verilog/coms.v(130[12] 305[6])
    defparam i15838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n51235), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15841_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n58011), 
            .I3(GND_net), .O(n29872));   // verilog/coms.v(130[12] 305[6])
    defparam i15841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_2106_26 (.CI(n51235), .I0(n3110), 
            .I1(VCC_net), .CO(n51236));
    SB_LUT4 i1_4_lut_adj_1896 (.I0(n2324), .I1(n2323), .I2(n2327), .I3(n2325), 
            .O(n62028));
    defparam i1_4_lut_adj_1896.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1897 (.I0(n2322), .I1(n2328), .I2(n2326), .I3(GND_net), 
            .O(n62030));
    defparam i1_3_lut_adj_1897.LUT_INIT = 16'hfefe;
    SB_LUT4 i15844_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n58011), 
            .I3(GND_net), .O(n29875));   // verilog/coms.v(130[12] 305[6])
    defparam i15844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15847_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n58011), 
            .I3(GND_net), .O(n29878));   // verilog/coms.v(130[12] 305[6])
    defparam i15847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29172_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n43099));
    defparam i29172_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i26_4_lut (.I0(n110), .I1(n66446), .I2(state[1]), .I3(n4_adj_5926), 
            .O(n56711));   // verilog/neopixel.v(34[12] 116[6])
    defparam i26_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 encoder0_position_30__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15850_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n58011), 
            .I3(GND_net), .O(n29881));   // verilog/coms.v(130[12] 305[6])
    defparam i15850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n57742));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i15854_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n58897), 
            .I3(GND_net), .O(n29885));   // verilog/coms.v(130[12] 305[6])
    defparam i15854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n57743));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n50535), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5814), .CO(n50536));
    SB_LUT4 encoder0_position_30__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n51234), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_14 (.CI(n50673), .I0(n1522), 
            .I1(VCC_net), .CO(n50674));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n57744));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n57745));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n57746));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n57747));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n28932));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n57748));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n50672), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_23 (.CI(n50429), .I0(GND_net), .I1(n12146), .CO(n50430));
    SB_LUT4 i1_4_lut_adj_1905 (.I0(n2320), .I1(n2321), .I2(n62030), .I3(n62028), 
            .O(n62036));
    defparam i1_4_lut_adj_1905.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[21] [5]), .I1(n28300), .I2(n28355), 
            .I3(rx_data[5]), .O(n57155));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5825));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n57749));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1907 (.I0(\data_in_frame[21] [4]), .I1(n28300), 
            .I2(n28355), .I3(rx_data[4]), .O(n57159));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1907.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_30__I_0_add_2106_25 (.CI(n51234), .I0(n3111), 
            .I1(VCC_net), .CO(n51235));
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n56483));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n57750));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i14791_4_lut (.I0(n27735), .I1(n1319), .I2(n66302), .I3(n42285), 
            .O(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i14791_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1909 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n62506));
    defparam i1_2_lut_adj_1909.LUT_INIT = 16'h8888;
    SB_LUT4 i16512_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2874));   // verilog/coms.v(130[12] 305[6])
    defparam i16512_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n57751));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n57752));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1912 (.I0(\data_in_frame[21] [3]), .I1(n28300), 
            .I2(n28355), .I3(rx_data[3]), .O(n57163));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1912.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n51233), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1913 (.I0(\data_in_frame[21] [2]), .I1(n28300), 
            .I2(n28355), .I3(rx_data[2]), .O(n57167));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1913.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n57753));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n57754));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n28924));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1917 (.I0(\data_in_frame[21] [1]), .I1(n28300), 
            .I2(n28355), .I3(rx_data[1]), .O(n57169));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1917.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n57755));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n57756));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n57757));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1921 (.I0(n62506), .I1(n2319), .I2(n62036), .I3(n43099), 
            .O(n62040));
    defparam i1_4_lut_adj_1921.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1922 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n62040), 
            .O(n62046));
    defparam i1_4_lut_adj_1922.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1923 (.I0(n5_adj_5929), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n62448));
    defparam i1_3_lut_adj_1923.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5813), .I3(n50534), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n57758));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n57759));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h2300;
    SB_LUT4 add_1100_22_lut (.I0(GND_net), .I1(GND_net), .I2(n12148), 
            .I3(n50428), .O(n4910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n57760));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1927 (.I0(n8_adj_5779), .I1(n40525), .I2(GND_net), 
            .I3(GND_net), .O(n28300));
    defparam i1_2_lut_adj_1927.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12_4_lut_adj_1928 (.I0(\data_in_frame[21] [0]), .I1(n28300), 
            .I2(n28355), .I3(rx_data[0]), .O(n57117));
    defparam i12_4_lut_adj_1928.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_i500_4_lut (.I0(n2_adj_5778), .I1(n7444), 
            .I2(n62448), .I3(encoder0_position[30]), .O(n828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_CARRY add_1100_22 (.CI(n50428), .I0(GND_net), .I1(n12148), .CO(n50429));
    SB_LUT4 i12_4_lut_adj_1929 (.I0(\data_in_frame[17] [7]), .I1(n28308), 
            .I2(n28363), .I3(rx_data[7]), .O(n57187));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1929.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n66280), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5755));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16138_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n28363), .I3(GND_net), .O(n30169));   // verilog/coms.v(130[12] 305[6])
    defparam i16138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5766));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5764));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51316_2_lut (.I0(n70252), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n66452));
    defparam i51316_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n50534), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5813), .CO(n50535));
    SB_LUT4 i12_4_lut_adj_1930 (.I0(\data_in_frame[17] [5]), .I1(n28308), 
            .I2(n28363), .I3(rx_data[5]), .O(n57191));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1930.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_30__I_0_add_2106_24 (.CI(n51233), .I0(n3112), 
            .I1(VCC_net), .CO(n51234));
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5758));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1034_13 (.CI(n50672), .I0(n1523), 
            .I1(VCC_net), .CO(n50673));
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5757));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5756));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n51232), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1931 (.I0(\data_in_frame[17] [4]), .I1(n28308), 
            .I2(n28363), .I3(rx_data[4]), .O(n57195));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1931.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_adj_1932 (.I0(n8_adj_5704), .I1(n40525), .I2(GND_net), 
            .I3(GND_net), .O(n28308));
    defparam i1_2_lut_adj_1932.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_30__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1933 (.I0(\data_in_frame[17] [3]), .I1(n28308), 
            .I2(n28363), .I3(rx_data[3]), .O(n57199));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1933.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5762));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5761));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5760));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27735), 
            .D(n1239), .R(n28822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5702));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5703));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n28917));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n41_adj_5917));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n57761));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 i16118_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n28363), .I3(GND_net), .O(n30149));   // verilog/coms.v(130[12] 305[6])
    defparam i16118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5706));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1937 (.I0(\data_in_frame[16] [7]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[7]), .O(n57203));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1937.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_30__I_0_add_2106_23 (.CI(n51232), .I0(n3113), 
            .I1(VCC_net), .CO(n51233));
    SB_LUT4 i12_4_lut_adj_1938 (.I0(\data_in_frame[16] [6]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[6]), .O(n57207));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1938.LUT_INIT = 16'h3a0a;
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n27648), .D(GHC_N_391), 
            .R(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n27648), .D(GHB_N_377), 
            .R(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n27648), .D(GHA_N_355), 
            .R(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5942), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i12_4_lut_adj_1939 (.I0(\data_in_frame[16] [5]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[5]), .O(n57211));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1939.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n57762));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1941 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n57763));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1941.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5705));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1942 (.I0(\data_in_frame[16] [4]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[4]), .O(n57215));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1942.LUT_INIT = 16'h3a0a;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[25]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[24]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n27648), .D(GLA_N_372), 
            .R(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n27648), .D(GLB_N_386), 
            .R(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n27648), .D(GLC_N_400), 
            .R(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n25_adj_5724));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5708));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    GND i1 (.Y(GND_net));
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n50313), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n50671), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5811), .I3(n50533), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n50313), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n50314));
    SB_LUT4 add_1100_21_lut (.I0(GND_net), .I1(GND_net), .I2(n12150), 
            .I3(n50427), .O(n4911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n50533), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5811), .CO(n50534));
    SB_LUT4 encoder0_position_30__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n51231), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_12 (.CI(n50671), .I0(n1524), 
            .I1(VCC_net), .CO(n50672));
    SB_CARRY encoder0_position_30__I_0_add_2106_22 (.CI(n51231), .I0(n3114), 
            .I1(VCC_net), .CO(n51232));
    SB_CARRY add_1100_21 (.CI(n50427), .I0(GND_net), .I1(n12150), .CO(n50428));
    SB_LUT4 encoder0_position_30__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n51230), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n50670), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_20_lut (.I0(GND_net), .I1(GND_net), .I2(n12152), 
            .I3(n50426), .O(n4912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_21 (.CI(n51230), .I0(n3115), 
            .I1(VCC_net), .CO(n51231));
    SB_LUT4 encoder0_position_30__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n51229), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_11 (.CI(n50670), .I0(n1525), 
            .I1(VCC_net), .CO(n50671));
    SB_CARRY add_1100_20 (.CI(n50426), .I0(GND_net), .I1(n12152), .CO(n50427));
    SB_LUT4 add_1100_19_lut (.I0(GND_net), .I1(GND_net), .I2(n12154), 
            .I3(n50425), .O(n4913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_22_lut (.I0(n69870), .I1(n2214), 
            .I2(VCC_net), .I3(n50898), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n50897), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_21 (.CI(n50897), .I0(n2215), 
            .I1(VCC_net), .CO(n50898));
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5709));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n50669), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_20 (.CI(n51229), .I0(n3116), 
            .I1(VCC_net), .CO(n51230));
    SB_LUT4 encoder0_position_30__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n50896), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5802), .I3(n50532), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n51228), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_19 (.CI(n51228), .I0(n3117), 
            .I1(VCC_net), .CO(n51229));
    SB_CARRY add_1100_19 (.CI(n50425), .I0(GND_net), .I1(n12154), .CO(n50426));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n50312), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n50299), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_10 (.CI(n50669), .I0(n1526), 
            .I1(VCC_net), .CO(n50670));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n50532), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5802), .CO(n50533));
    SB_CARRY encoder0_position_30__I_0_add_1503_20 (.CI(n50896), .I0(n2216), 
            .I1(VCC_net), .CO(n50897));
    SB_LUT4 add_1100_18_lut (.I0(GND_net), .I1(GND_net), .I2(n12156), 
            .I3(n50424), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n50668), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n50895), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_18 (.CI(n50424), .I0(GND_net), .I1(n12156), .CO(n50425));
    SB_LUT4 add_1100_17_lut (.I0(GND_net), .I1(GND_net), .I2(n12158), 
            .I3(n50423), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5801), .I3(n50531), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_19 (.CI(n50895), .I0(n2217), 
            .I1(VCC_net), .CO(n50896));
    SB_LUT4 i51425_4_lut (.I0(n11_adj_5705), .I1(n9_adj_5706), .I2(n7_adj_5708), 
            .I3(n5_adj_5709), .O(n67151));
    defparam i51425_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n28911));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_CARRY add_151_23 (.CI(n50312), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n50313));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n50531), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5801), .CO(n50532));
    SB_LUT4 encoder0_position_30__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n51227), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n50894), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_9 (.CI(n50668), .I0(n1527), 
            .I1(VCC_net), .CO(n50669));
    SB_CARRY encoder0_position_30__I_0_add_1503_18 (.CI(n50894), .I0(n2218), 
            .I1(VCC_net), .CO(n50895));
    SB_CARRY add_1100_17 (.CI(n50423), .I0(GND_net), .I1(n12158), .CO(n50424));
    SB_LUT4 encoder0_position_30__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n50667), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n50893), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_18 (.CI(n51227), .I0(n3118), 
            .I1(VCC_net), .CO(n51228));
    SB_LUT4 add_1100_16_lut (.I0(GND_net), .I1(GND_net), .I2(n12160), 
            .I3(n50422), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5800), .I3(n50530), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_17 (.CI(n50893), .I0(n2219), 
            .I1(VCC_net), .CO(n50894));
    SB_CARRY encoder0_position_30__I_0_add_1034_8 (.CI(n50667), .I0(n1528), 
            .I1(VCC_net), .CO(n50668));
    SB_LUT4 encoder0_position_30__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n50892), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n50530), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5800), .CO(n50531));
    SB_LUT4 encoder0_position_30__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n51226), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_16 (.CI(n50892), .I0(n2220), 
            .I1(VCC_net), .CO(n50893));
    SB_CARRY add_1100_16 (.CI(n50422), .I0(GND_net), .I1(n12160), .CO(n50423));
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n50311), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n50666), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_7 (.CI(n50666), .I0(n1529), 
            .I1(GND_net), .CO(n50667));
    SB_LUT4 encoder0_position_30__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n50891), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_15 (.CI(n50891), .I0(n2221), 
            .I1(VCC_net), .CO(n50892));
    SB_CARRY add_151_22 (.CI(n50311), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n50312));
    SB_LUT4 add_1100_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12162), 
            .I3(n50421), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_15 (.CI(n50421), .I0(GND_net), .I1(n12162), .CO(n50422));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5722), .I3(n50529), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n50890), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_17 (.CI(n51226), .I0(n3119), 
            .I1(VCC_net), .CO(n51227));
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i15575_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n58009), 
            .I3(GND_net), .O(n29606));   // verilog/coms.v(130[12] 305[6])
    defparam i15575_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n50529), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5722), .CO(n50530));
    SB_LUT4 add_1100_14_lut (.I0(GND_net), .I1(GND_net), .I2(n12164), 
            .I3(n50420), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_14 (.CI(n50890), .I0(n2222), 
            .I1(VCC_net), .CO(n50891));
    SB_LUT4 encoder0_position_30__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n51225), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_10 (.CI(n50299), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n50300));
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n50298), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n50665), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n50889), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_13 (.CI(n50889), .I0(n2223), 
            .I1(VCC_net), .CO(n50890));
    SB_CARRY encoder0_position_30__I_0_add_2106_16 (.CI(n51225), .I0(n3120), 
            .I1(VCC_net), .CO(n51226));
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n50310), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_6 (.CI(n50665), .I0(n1530), 
            .I1(GND_net), .CO(n50666));
    SB_CARRY add_1100_14 (.CI(n50420), .I0(GND_net), .I1(n12164), .CO(n50421));
    SB_LUT4 add_1100_13_lut (.I0(GND_net), .I1(GND_net), .I2(n12166), 
            .I3(n50419), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_13 (.CI(n50419), .I0(GND_net), .I1(n12166), .CO(n50420));
    SB_LUT4 encoder0_position_30__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n50888), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_12 (.CI(n50888), .I0(n2224), 
            .I1(VCC_net), .CO(n50889));
    SB_LUT4 encoder0_position_30__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n51224), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n50887), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_4 (.CI(n50293), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n50294));
    SB_CARRY encoder0_position_30__I_0_add_1503_11 (.CI(n50887), .I0(n2225), 
            .I1(VCC_net), .CO(n50888));
    SB_CARRY encoder0_position_30__I_0_add_2106_15 (.CI(n51224), .I0(n3121), 
            .I1(VCC_net), .CO(n51225));
    SB_LUT4 encoder0_position_30__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n50664), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n51223), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_14 (.CI(n51223), .I0(n3122), 
            .I1(VCC_net), .CO(n51224));
    SB_LUT4 encoder0_position_30__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n50886), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n51222), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_12_lut (.I0(GND_net), .I1(GND_net), .I2(n12168), 
            .I3(n50418), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_13 (.CI(n51222), .I0(n3123), 
            .I1(VCC_net), .CO(n51223));
    SB_CARRY encoder0_position_30__I_0_add_1503_10 (.CI(n50886), .I0(n2226), 
            .I1(VCC_net), .CO(n50887));
    SB_LUT4 encoder0_position_30__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n50885), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_9 (.CI(n50885), .I0(n2227), 
            .I1(VCC_net), .CO(n50886));
    SB_LUT4 encoder0_position_30__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n51221), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n50884), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_26_lut (.I0(GND_net), .I1(n2610), 
            .I2(VCC_net), .I3(n51083), .O(n2677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_12 (.CI(n50418), .I0(GND_net), .I1(n12168), .CO(n50419));
    SB_LUT4 encoder0_position_30__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n51082), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_8 (.CI(n50884), .I0(n2228), 
            .I1(VCC_net), .CO(n50885));
    SB_CARRY encoder0_position_30__I_0_add_2106_12 (.CI(n51221), .I0(n3124), 
            .I1(VCC_net), .CO(n51222));
    SB_LUT4 encoder0_position_30__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n50883), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_7 (.CI(n50883), .I0(n2229), 
            .I1(GND_net), .CO(n50884));
    SB_LUT4 add_1100_11_lut (.I0(GND_net), .I1(GND_net), .I2(n12170), 
            .I3(n50417), .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_5 (.CI(n50664), .I0(n1531), 
            .I1(VCC_net), .CO(n50665));
    SB_CARRY add_1100_11 (.CI(n50417), .I0(GND_net), .I1(n12170), .CO(n50418));
    SB_CARRY add_151_9 (.CI(n50298), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n50299));
    SB_LUT4 encoder0_position_30__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n50663), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_21 (.CI(n50310), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n50311));
    SB_CARRY encoder0_position_30__I_0_add_1771_25 (.CI(n51082), .I0(n2611), 
            .I1(VCC_net), .CO(n51083));
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n50309), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n50882), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_4 (.CI(n50663), .I0(n1532), 
            .I1(GND_net), .CO(n50664));
    SB_CARRY encoder0_position_30__I_0_add_1503_6 (.CI(n50882), .I0(n2230), 
            .I1(GND_net), .CO(n50883));
    SB_LUT4 encoder0_position_30__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n51081), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n50881), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_10_lut (.I0(GND_net), .I1(GND_net), .I2(n12172), 
            .I3(n50416), .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_10 (.CI(n50416), .I0(GND_net), .I1(n12172), .CO(n50417));
    SB_CARRY add_151_20 (.CI(n50309), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n50310));
    SB_LUT4 encoder0_position_30__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n50662), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_9_lut (.I0(GND_net), .I1(GND_net), .I2(n12174), .I3(n50415), 
            .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_3 (.CI(n50662), .I0(n1533), 
            .I1(VCC_net), .CO(n50663));
    SB_LUT4 encoder0_position_30__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_5 (.CI(n50881), .I0(n2231), 
            .I1(VCC_net), .CO(n50882));
    SB_LUT4 encoder0_position_30__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n51220), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_9 (.CI(n50415), .I0(GND_net), .I1(n12174), .CO(n50416));
    SB_LUT4 add_1100_8_lut (.I0(GND_net), .I1(GND_net), .I2(n12176), .I3(n50414), 
            .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5721), .I3(n50528), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n50880), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_24 (.CI(n51081), .I0(n2612), 
            .I1(VCC_net), .CO(n51082));
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n50292), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n50297), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_8 (.CI(n50297), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n50298));
    SB_CARRY add_1100_8 (.CI(n50414), .I0(GND_net), .I1(n12176), .CO(n50415));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n50528), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5721), .CO(n50529));
    SB_CARRY encoder0_position_30__I_0_add_2106_11 (.CI(n51220), .I0(n3125), 
            .I1(VCC_net), .CO(n51221));
    SB_CARRY encoder0_position_30__I_0_add_1503_4 (.CI(n50880), .I0(n2232), 
            .I1(GND_net), .CO(n50881));
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5707), .I1(current_limit[9]), 
            .I2(n19), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5710));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n50308), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n50879), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n50662));
    SB_LUT4 encoder0_position_30__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n51080), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_3 (.CI(n50879), .I0(n2233), 
            .I1(VCC_net), .CO(n50880));
    SB_CARRY add_151_19 (.CI(n50308), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n50309));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n50296), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_14_lut (.I0(n70042), .I1(n1422), 
            .I2(VCC_net), .I3(n50661), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5720), .I3(n50527), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_7_lut (.I0(GND_net), .I1(GND_net), .I2(n12178), .I3(n50413), 
            .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n50527), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5720), .CO(n50528));
    SB_CARRY encoder0_position_30__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n50879));
    SB_LUT4 encoder0_position_30__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n50660), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n51219), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52955_3_lut (.I0(n4_adj_5710), .I1(current_limit[5]), .I2(n11_adj_5705), 
            .I3(GND_net), .O(n68681));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52955_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1771_23 (.CI(n51080), .I0(n2613), 
            .I1(VCC_net), .CO(n51081));
    SB_CARRY encoder0_position_30__I_0_add_967_13 (.CI(n50660), .I0(n1423), 
            .I1(VCC_net), .CO(n50661));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5719), .I3(n50526), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_10 (.CI(n51219), .I0(n3126), 
            .I1(VCC_net), .CO(n51220));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n50526), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5719), .CO(n50527));
    SB_CARRY add_1100_7 (.CI(n50413), .I0(GND_net), .I1(n12178), .CO(n50414));
    SB_LUT4 encoder0_position_30__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n50659), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n51079), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n51218), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n50307), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1100_6_lut (.I0(GND_net), .I1(GND_net), .I2(n12180), .I3(n50412), 
            .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_9 (.CI(n51218), .I0(n3127), 
            .I1(VCC_net), .CO(n51219));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5717), .I3(n50525), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_22 (.CI(n51079), .I0(n2614), 
            .I1(VCC_net), .CO(n51080));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n50525), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5717), .CO(n50526));
    SB_LUT4 encoder0_position_30__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n51217), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_3 (.CI(n50292), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n50293));
    SB_LUT4 encoder0_position_30__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n51078), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_8 (.CI(n51217), .I0(n3128), 
            .I1(VCC_net), .CO(n51218));
    SB_CARRY encoder0_position_30__I_0_add_1771_21 (.CI(n51078), .I0(n2615), 
            .I1(VCC_net), .CO(n51079));
    SB_LUT4 i52956_3_lut (.I0(n68681), .I1(current_limit[6]), .I2(n13_adj_5703), 
            .I3(GND_net), .O(n68682));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n51077), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n51216), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_20 (.CI(n51077), .I0(n2616), 
            .I1(VCC_net), .CO(n51078));
    SB_LUT4 encoder0_position_30__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n51076), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_19 (.CI(n51076), .I0(n2617), 
            .I1(VCC_net), .CO(n51077));
    SB_CARRY encoder0_position_30__I_0_add_2106_7 (.CI(n51216), .I0(n3129), 
            .I1(GND_net), .CO(n51217));
    SB_LUT4 encoder0_position_30__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n51075), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n51215), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1945 (.I0(\data_in_frame[16] [3]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[3]), .O(n57219));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1945.LUT_INIT = 16'h3a0a;
    SB_CARRY add_151_7 (.CI(n50296), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n50297));
    SB_CARRY encoder0_position_30__I_0_add_967_12 (.CI(n50659), .I0(n1424), 
            .I1(VCC_net), .CO(n50660));
    SB_LUT4 encoder0_position_30__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n50658), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_6 (.CI(n50412), .I0(GND_net), .I1(n12180), .CO(n50413));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5716), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_18 (.CI(n51075), .I0(n2618), 
            .I1(VCC_net), .CO(n51076));
    SB_CARRY encoder0_position_30__I_0_add_967_11 (.CI(n50658), .I0(n1425), 
            .I1(VCC_net), .CO(n50659));
    SB_LUT4 add_1100_5_lut (.I0(GND_net), .I1(GND_net), .I2(n10), .I3(n50411), 
            .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5716), .CO(n50525));
    SB_CARRY encoder0_position_30__I_0_add_2106_6 (.CI(n51215), .I0(n3130), 
            .I1(GND_net), .CO(n51216));
    SB_LUT4 i12_4_lut_adj_1946 (.I0(\data_in_frame[16] [2]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[2]), .O(n57221));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1946.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n50657), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_10 (.CI(n50657), .I0(n1426), 
            .I1(VCC_net), .CO(n50658));
    SB_CARRY add_1100_5 (.CI(n50411), .I0(GND_net), .I1(n10), .CO(n50412));
    SB_LUT4 add_1100_4_lut (.I0(GND_net), .I1(GND_net), .I2(n12184), .I3(n50410), 
            .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n51074), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_4 (.CI(n50410), .I0(GND_net), .I1(n12184), .CO(n50411));
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n51214), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_17 (.CI(n51074), .I0(n2619), 
            .I1(VCC_net), .CO(n51075));
    SB_CARRY add_151_18 (.CI(n50307), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n50308));
    SB_LUT4 encoder0_position_30__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n50656), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_9 (.CI(n50656), .I0(n1427), 
            .I1(VCC_net), .CO(n50657));
    SB_LUT4 add_1100_3_lut (.I0(GND_net), .I1(GND_net), .I2(n12186), .I3(n50409), 
            .O(n4929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_3 (.CI(n50409), .I0(GND_net), .I1(n12186), .CO(n50410));
    SB_CARRY encoder0_position_30__I_0_add_2106_5 (.CI(n51214), .I0(n3131), 
            .I1(VCC_net), .CO(n51215));
    SB_LUT4 add_1100_2_lut (.I0(GND_net), .I1(GND_net), .I2(n5), .I3(VCC_net), 
            .O(n4930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1100_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n50655), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_8 (.CI(n50655), .I0(n1428), 
            .I1(VCC_net), .CO(n50656));
    SB_LUT4 encoder0_position_30__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n51213), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1100_2 (.CI(VCC_net), .I0(GND_net), .I1(n5), .CO(n50409));
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n50295), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n51073), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_16 (.CI(n51073), .I0(n2620), 
            .I1(VCC_net), .CO(n51074));
    SB_CARRY encoder0_position_30__I_0_add_2106_4 (.CI(n51213), .I0(n3132), 
            .I1(GND_net), .CO(n51214));
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n50306), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n51072), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n51212), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_3 (.CI(n51212), .I0(n3133), 
            .I1(VCC_net), .CO(n51213));
    SB_CARRY encoder0_position_30__I_0_add_1771_15 (.CI(n51072), .I0(n2621), 
            .I1(VCC_net), .CO(n51073));
    SB_LUT4 encoder0_position_30__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n50654), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n51071), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_14 (.CI(n51071), .I0(n2622), 
            .I1(VCC_net), .CO(n51072));
    SB_LUT4 encoder0_position_30__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n50292));
    SB_CARRY encoder0_position_30__I_0_add_967_7 (.CI(n50654), .I0(n1429), 
            .I1(GND_net), .CO(n50655));
    SB_LUT4 encoder0_position_30__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n51070), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n51212));
    SB_CARRY encoder0_position_30__I_0_add_1771_13 (.CI(n51070), .I0(n2623), 
            .I1(VCC_net), .CO(n51071));
    SB_LUT4 encoder0_position_30__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n51069), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_12 (.CI(n51069), .I0(n2624), 
            .I1(VCC_net), .CO(n51070));
    SB_CARRY add_151_17 (.CI(n50306), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n50307));
    SB_LUT4 encoder0_position_30__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n51068), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n50305), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n50653), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_6 (.CI(n50653), .I0(n1430), 
            .I1(GND_net), .CO(n50654));
    SB_LUT4 encoder0_position_30__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n50652), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_30_lut (.I0(n69620), .I1(n3006), 
            .I2(VCC_net), .I3(n51211), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n51210), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_5 (.CI(n50652), .I0(n1431), 
            .I1(VCC_net), .CO(n50653));
    SB_CARRY encoder0_position_30__I_0_add_1771_11 (.CI(n51068), .I0(n2625), 
            .I1(VCC_net), .CO(n51069));
    SB_LUT4 encoder0_position_30__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n51067), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n50651), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_6 (.CI(n50295), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n50296));
    SB_CARRY encoder0_position_30__I_0_add_2039_29 (.CI(n51210), .I0(n3007), 
            .I1(VCC_net), .CO(n51211));
    SB_CARRY add_151_16 (.CI(n50305), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n50306));
    SB_CARRY encoder0_position_30__I_0_add_1771_10 (.CI(n51067), .I0(n2626), 
            .I1(VCC_net), .CO(n51068));
    SB_CARRY encoder0_position_30__I_0_add_967_4 (.CI(n50651), .I0(n1432), 
            .I1(GND_net), .CO(n50652));
    SB_LUT4 encoder0_position_30__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n51209), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n51066), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1947 (.I0(\data_in_frame[16] [1]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[1]), .O(n57223));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1947.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n50650), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_9 (.CI(n51066), .I0(n2627), 
            .I1(VCC_net), .CO(n51067));
    SB_CARRY encoder0_position_30__I_0_add_967_3 (.CI(n50650), .I0(n1433), 
            .I1(VCC_net), .CO(n50651));
    SB_LUT4 encoder0_position_30__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n50650));
    SB_LUT4 encoder0_position_30__I_0_add_900_13_lut (.I0(n70007), .I1(n1323), 
            .I2(VCC_net), .I3(n50649), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n50648), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_12 (.CI(n50648), .I0(n1324), 
            .I1(VCC_net), .CO(n50649));
    SB_CARRY encoder0_position_30__I_0_add_2039_28 (.CI(n51209), .I0(n3008), 
            .I1(VCC_net), .CO(n51210));
    SB_LUT4 encoder0_position_30__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n28910));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n51065), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n51208), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_27 (.CI(n51208), .I0(n3009), 
            .I1(VCC_net), .CO(n51209));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n50304), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n51207), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_8 (.CI(n51065), .I0(n2628), 
            .I1(VCC_net), .CO(n51066));
    SB_LUT4 encoder0_position_30__I_0_add_1436_21_lut (.I0(n69845), .I1(n2115), 
            .I2(VCC_net), .I3(n50854), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n51064), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n50853), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_26 (.CI(n51207), .I0(n3010), 
            .I1(VCC_net), .CO(n51208));
    SB_LUT4 encoder0_position_30__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n51206), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_7 (.CI(n51064), .I0(n2629), 
            .I1(GND_net), .CO(n51065));
    SB_CARRY encoder0_position_30__I_0_add_2039_25 (.CI(n51206), .I0(n3011), 
            .I1(VCC_net), .CO(n51207));
    SB_CARRY encoder0_position_30__I_0_add_1436_20 (.CI(n50853), .I0(n2116), 
            .I1(VCC_net), .CO(n50854));
    SB_LUT4 encoder0_position_30__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n51063), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_6 (.CI(n51063), .I0(n2630), 
            .I1(GND_net), .CO(n51064));
    SB_LUT4 i53811_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n62046), 
            .O(n2346));
    defparam i53811_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_1949 (.I0(n8_adj_5790), .I1(n40525), .I2(GND_net), 
            .I3(GND_net), .O(n28310));
    defparam i1_2_lut_adj_1949.LUT_INIT = 16'hbbbb;
    SB_LUT4 i51407_4_lut (.I0(n17), .I1(n15_adj_5702), .I2(n13_adj_5703), 
            .I3(n67151), .O(n67133));
    defparam i51407_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53336_4_lut (.I0(n16), .I1(n6), .I2(n19), .I3(n67123), 
            .O(n69062));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53336_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51793_3_lut (.I0(n68682), .I1(current_limit[7]), .I2(n15_adj_5702), 
            .I3(GND_net), .O(n67519));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n51062), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_15 (.CI(n50304), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n50305));
    SB_CARRY encoder0_position_30__I_0_add_1771_5 (.CI(n51062), .I0(n2631), 
            .I1(VCC_net), .CO(n51063));
    SB_LUT4 encoder0_position_30__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n51061), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n50852), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_19 (.CI(n50852), .I0(n2117), 
            .I1(VCC_net), .CO(n50853));
    SB_LUT4 encoder0_position_30__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n50851), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_4 (.CI(n51061), .I0(n2632), 
            .I1(GND_net), .CO(n51062));
    SB_CARRY encoder0_position_30__I_0_add_1436_18 (.CI(n50851), .I0(n2118), 
            .I1(VCC_net), .CO(n50852));
    SB_LUT4 encoder0_position_30__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n50647), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n51205), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_24 (.CI(n51205), .I0(n3012), 
            .I1(VCC_net), .CO(n51206));
    SB_LUT4 encoder0_position_30__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n51060), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n51204), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_11 (.CI(n50647), .I0(n1325), 
            .I1(VCC_net), .CO(n50648));
    SB_LUT4 i53496_4_lut (.I0(n67519), .I1(n69062), .I2(n19), .I3(n67133), 
            .O(n69222));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53496_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53497_3_lut (.I0(n69222), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n69223));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53497_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_1771_3 (.CI(n51060), .I0(n2633), 
            .I1(VCC_net), .CO(n51061));
    SB_LUT4 encoder0_position_30__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n50850), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_17 (.CI(n50850), .I0(n2119), 
            .I1(VCC_net), .CO(n50851));
    SB_CARRY encoder0_position_30__I_0_add_2039_23 (.CI(n51204), .I0(n3013), 
            .I1(VCC_net), .CO(n51205));
    SB_CARRY encoder0_position_30__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n51060));
    SB_LUT4 encoder0_position_30__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n50849), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53426_3_lut (.I0(n69223), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n69152));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53426_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_14_i26_3_lut (.I0(n69152), .I1(current_limit[12]), 
            .I2(current[15]), .I3(GND_net), .O(n26_adj_5701));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_1436_16 (.CI(n50849), .I0(n2120), 
            .I1(VCC_net), .CO(n50850));
    SB_LUT4 encoder0_position_30__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n50848), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n50646), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n51203), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_10 (.CI(n50646), .I0(n1326), 
            .I1(VCC_net), .CO(n50647));
    SB_LUT4 encoder0_position_30__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n50645), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_22 (.CI(n51203), .I0(n3014), 
            .I1(VCC_net), .CO(n51204));
    SB_LUT4 encoder0_position_30__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1950 (.I0(n2427), .I1(n2425), .I2(n2426), .I3(n2424), 
            .O(n62514));
    defparam i1_4_lut_adj_1950.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1951 (.I0(\data_in_frame[16] [0]), .I1(n28310), 
            .I2(n28365), .I3(rx_data[0]), .O(n57225));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1951.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n57764));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n57765));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5715));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n57766));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n57767));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(duty[11]), .I1(n299), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5723));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(duty[10]), .I1(n300), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5788));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5718));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32_3_lut (.I0(n4), .I1(duty[2]), .I2(n308), .I3(GND_net), 
            .O(n26));   // verilog/TinyFPGA_B.v(96[21:25])
    defparam i32_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n57768));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n57769));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n51202), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_21 (.CI(n51202), .I0(n3015), 
            .I1(VCC_net), .CO(n51203));
    SB_LUT4 i23041_3_lut (.I0(n307), .I1(duty[3]), .I2(n26), .I3(GND_net), 
            .O(n8_adj_5700));   // verilog/TinyFPGA_B.v(96[21:25])
    defparam i23041_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n57770));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 i52965_3_lut (.I0(n8_adj_5700), .I1(n303), .I2(n15), .I3(GND_net), 
            .O(n68691));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n51201), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n57771));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_LUT4 i52966_3_lut (.I0(n68691), .I1(n302), .I2(n17_adj_5718), .I3(GND_net), 
            .O(n68692));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52966_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2039_20 (.CI(n51201), .I0(n3016), 
            .I1(VCC_net), .CO(n51202));
    SB_CARRY encoder0_position_30__I_0_add_1436_15 (.CI(n50848), .I0(n2121), 
            .I1(VCC_net), .CO(n50849));
    SB_LUT4 encoder0_position_30__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n50847), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n51200), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_14 (.CI(n50847), .I0(n2122), 
            .I1(VCC_net), .CO(n50848));
    SB_CARRY encoder0_position_30__I_0_add_2039_19 (.CI(n51200), .I0(n3017), 
            .I1(VCC_net), .CO(n51201));
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n57772));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n51199), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_18 (.CI(n51199), .I0(n3018), 
            .I1(VCC_net), .CO(n51200));
    SB_CARRY encoder0_position_30__I_0_add_900_9 (.CI(n50645), .I0(n1327), 
            .I1(VCC_net), .CO(n50646));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n57773));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n304), .I1(n300), .I2(n21_adj_5788), 
            .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n50644), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n51198), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n50846), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_13 (.CI(n50846), .I0(n2123), 
            .I1(VCC_net), .CO(n50847));
    SB_CARRY encoder0_position_30__I_0_add_900_8 (.CI(n50644), .I0(n1328), 
            .I1(VCC_net), .CO(n50645));
    SB_CARRY encoder0_position_30__I_0_add_2039_17 (.CI(n51198), .I0(n3019), 
            .I1(VCC_net), .CO(n51199));
    SB_LUT4 encoder0_position_30__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n51197), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n306), .I1(n305), .I2(n11), .I3(GND_net), 
            .O(n10_adj_5699));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i20_3_lut (.I0(n12), .I1(n299), .I2(n23_adj_5723), 
            .I3(GND_net), .O(n20_adj_5727));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n57774));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n57775));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 i51539_4_lut (.I0(n15), .I1(n13), .I2(n11), .I3(n9), .O(n67265));
    defparam i51539_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51474_4_lut (.I0(n21_adj_5788), .I1(n19_adj_5715), .I2(n17_adj_5718), 
            .I3(n67265), .O(n67200));
    defparam i51474_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52823_4_lut (.I0(n20_adj_5727), .I1(n10_adj_5699), .I2(n23_adj_5723), 
            .I3(n67196), .O(n68549));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52823_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51783_3_lut (.I0(n68692), .I1(n301), .I2(n19_adj_5715), .I3(GND_net), 
            .O(n67509));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53352_4_lut (.I0(n67509), .I1(n68549), .I2(n23_adj_5723), 
            .I3(n67200), .O(n69078));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53352_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47603_3_lut (.I0(duty[22]), .I1(duty[17]), .I2(n294), .I3(GND_net), 
            .O(n63312));
    defparam i47603_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i53353_3_lut (.I0(n69078), .I1(n298), .I2(duty[12]), .I3(GND_net), 
            .O(n69079));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53353_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47607_3_lut (.I0(duty[13]), .I1(duty[21]), .I2(n294), .I3(GND_net), 
            .O(n63316));
    defparam i47607_3_lut.LUT_INIT = 16'h7e7e;
    SB_CARRY encoder0_position_30__I_0_add_2039_16 (.CI(n51197), .I0(n3020), 
            .I1(VCC_net), .CO(n51198));
    SB_LUT4 i29098_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n43025));
    defparam i29098_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n57776));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n57777));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n57778));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n57779));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n28893));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n57899));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n50845), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_12 (.CI(n50845), .I0(n2124), 
            .I1(VCC_net), .CO(n50846));
    SB_LUT4 encoder0_position_30__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n51196), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47816_4_lut (.I0(duty[15]), .I1(n63312), .I2(duty[20]), .I3(n294), 
            .O(n63533));
    defparam i47816_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i47599_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n294), .I3(GND_net), 
            .O(n63308));
    defparam i47599_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n57898));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i10_4_lut (.I0(n294), .I1(n63533), .I2(n63316), .I3(n69079), 
            .O(n22_adj_5934));
    defparam i10_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n57897));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n57896));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i47814_4_lut (.I0(duty[19]), .I1(n63308), .I2(duty[16]), .I3(n294), 
            .O(n63531));
    defparam i47814_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i52230_3_lut (.I0(n15_adj_5760), .I1(n13_adj_5761), .I2(n11_adj_5762), 
            .I3(GND_net), .O(n67956));
    defparam i52230_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_30__I_0_add_2039_15 (.CI(n51196), .I0(n3021), 
            .I1(VCC_net), .CO(n51197));
    SB_LUT4 i52158_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n67956), .O(n67884));
    defparam i52158_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n57895));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51301_4_lut (.I0(n21_adj_5756), .I1(n19_adj_5757), .I2(n17_adj_5758), 
            .I3(n9_adj_5764), .O(n67027));
    defparam i51301_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_30__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n51195), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52250_4_lut (.I0(n9_adj_5764), .I1(n7_adj_5766), .I2(current[2]), 
            .I3(duty[2]), .O(n67976));
    defparam i52250_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n57894));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i52717_4_lut (.I0(n15_adj_5760), .I1(n13_adj_5761), .I2(n11_adj_5762), 
            .I3(n67976), .O(n68443));
    defparam i52717_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52697_4_lut (.I0(n21_adj_5756), .I1(n19_adj_5757), .I2(n17_adj_5758), 
            .I3(n68443), .O(n68423));
    defparam i52697_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 encoder0_position_30__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n50844), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_14 (.CI(n51195), .I0(n3022), 
            .I1(VCC_net), .CO(n51196));
    SB_CARRY encoder0_position_30__I_0_add_1436_11 (.CI(n50844), .I0(n2125), 
            .I1(VCC_net), .CO(n50845));
    SB_LUT4 encoder0_position_30__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n51194), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53262_4_lut (.I0(current[15]), .I1(n23_adj_5755), .I2(duty[12]), 
            .I3(n68423), .O(n68988));
    defparam i53262_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i52164_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n68988), .O(n67890));
    defparam i52164_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n57893));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n57892));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n57891));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5768));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i52947_3_lut (.I0(n4_adj_5768), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n68673));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52947_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52120_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5760), .O(n67846));
    defparam i52120_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i1_4_lut_adj_1978 (.I0(n62514), .I1(n2421), .I2(n2423), .I3(n2428), 
            .O(n62518));
    defparam i1_4_lut_adj_1978.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n57890));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n50643), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5754));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i51254_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n67884), .O(n66980));
    defparam i51254_4_lut.LUT_INIT = 16'h5adb;
    SB_CARRY encoder0_position_30__I_0_add_2039_13 (.CI(n51194), .I0(n3023), 
            .I1(VCC_net), .CO(n51195));
    SB_LUT4 encoder0_position_30__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n51193), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_12 (.CI(n51193), .I0(n3024), 
            .I1(VCC_net), .CO(n51194));
    SB_CARRY encoder0_position_30__I_0_add_900_7 (.CI(n50643), .I0(n1329), 
            .I1(GND_net), .CO(n50644));
    SB_LUT4 LessThan_11_i35_rep_84_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n70569));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_84_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n50843), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53338_3_lut (.I0(n30_adj_5754), .I1(n10_adj_5763), .I2(n67846), 
            .I3(GND_net), .O(n69064));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51799_4_lut (.I0(n68673), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n67525));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51799_4_lut.LUT_INIT = 16'h8f0e;
    SB_CARRY encoder0_position_30__I_0_add_1436_10 (.CI(n50843), .I0(n2126), 
            .I1(VCC_net), .CO(n50844));
    SB_LUT4 encoder0_position_30__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n50842), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n51192), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_9 (.CI(n50842), .I0(n2127), 
            .I1(VCC_net), .CO(n50843));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n57889));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2039_11 (.CI(n51192), .I0(n3025), 
            .I1(VCC_net), .CO(n51193));
    SB_LUT4 encoder0_position_30__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n50642), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n50841), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_6 (.CI(n50642), .I0(n1330), 
            .I1(GND_net), .CO(n50643));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n57888));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i52945_3_lut (.I0(n6_adj_5767), .I1(duty[10]), .I2(n21_adj_5756), 
            .I3(GND_net), .O(n68671));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52946_3_lut (.I0(n68671), .I1(duty[11]), .I2(n23_adj_5755), 
            .I3(GND_net), .O(n68672));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n51191), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52689_4_lut (.I0(current[15]), .I1(n23_adj_5755), .I2(duty[12]), 
            .I3(n67027), .O(n68415));
    defparam i52689_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5765), .I1(duty[9]), .I2(n19_adj_5757), 
            .I3(GND_net), .O(n16_adj_5759));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1436_8 (.CI(n50841), .I0(n2128), 
            .I1(VCC_net), .CO(n50842));
    SB_LUT4 encoder0_position_30__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n50840), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_10 (.CI(n51191), .I0(n3026), 
            .I1(VCC_net), .CO(n51192));
    SB_LUT4 i51801_3_lut (.I0(n68672), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n67527));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51801_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n50641), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n57887));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1436_7 (.CI(n50840), .I0(n2129), 
            .I1(GND_net), .CO(n50841));
    SB_CARRY encoder0_position_30__I_0_add_900_5 (.CI(n50641), .I0(n1331), 
            .I1(VCC_net), .CO(n50642));
    SB_LUT4 encoder0_position_30__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n51190), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n50839), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_6 (.CI(n50839), .I0(n2130), 
            .I1(GND_net), .CO(n50840));
    SB_LUT4 encoder0_position_30__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n50838), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_9 (.CI(n51190), .I0(n3027), 
            .I1(VCC_net), .CO(n51191));
    SB_LUT4 encoder0_position_30__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n51189), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_5 (.CI(n50838), .I0(n2131), 
            .I1(VCC_net), .CO(n50839));
    SB_CARRY encoder0_position_30__I_0_add_2039_8 (.CI(n51189), .I0(n3028), 
            .I1(VCC_net), .CO(n51190));
    SB_LUT4 encoder0_position_30__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n50640), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n50837), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_4 (.CI(n50640), .I0(n1332), 
            .I1(GND_net), .CO(n50641));
    SB_LUT4 encoder0_position_30__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n51188), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_7 (.CI(n51188), .I0(n3029), 
            .I1(GND_net), .CO(n51189));
    SB_CARRY encoder0_position_30__I_0_add_1436_4 (.CI(n50837), .I0(n2132), 
            .I1(GND_net), .CO(n50838));
    SB_LUT4 encoder0_position_30__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n51187), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_6 (.CI(n51187), .I0(n3030), 
            .I1(GND_net), .CO(n51188));
    SB_LUT4 encoder0_position_30__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n51186), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n50639), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_5 (.CI(n51186), .I0(n3031), 
            .I1(VCC_net), .CO(n51187));
    SB_LUT4 i53023_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n67890), .O(n68749));
    defparam i53023_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n57886));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_900_3 (.CI(n50639), .I0(n1333), 
            .I1(VCC_net), .CO(n50640));
    SB_LUT4 encoder0_position_30__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n50836), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_3 (.CI(n50836), .I0(n2133), 
            .I1(VCC_net), .CO(n50837));
    SB_LUT4 encoder0_position_30__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n50836));
    SB_LUT4 encoder0_position_30__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n51185), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n50639));
    SB_CARRY encoder0_position_30__I_0_add_2039_4 (.CI(n51185), .I0(n3032), 
            .I1(GND_net), .CO(n51186));
    SB_LUT4 encoder0_position_30__I_0_add_833_12_lut (.I0(n69991), .I1(n1224_adj_5836), 
            .I2(VCC_net), .I3(n50638), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n51184), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225_adj_5837), 
            .I2(VCC_net), .I3(n50637), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_3 (.CI(n51184), .I0(n3033), 
            .I1(VCC_net), .CO(n51185));
    SB_CARRY encoder0_position_30__I_0_add_833_11 (.CI(n50637), .I0(n1225_adj_5837), 
            .I1(VCC_net), .CO(n50638));
    SB_LUT4 encoder0_position_30__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226_adj_5838), 
            .I2(VCC_net), .I3(n50636), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n51184));
    SB_LUT4 encoder0_position_30__I_0_add_1972_29_lut (.I0(n69587), .I1(n2907), 
            .I2(VCC_net), .I3(n51183), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_833_10 (.CI(n50636), .I0(n1226_adj_5838), 
            .I1(VCC_net), .CO(n50637));
    SB_LUT4 encoder0_position_30__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n51182), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227_adj_5839), 
            .I2(VCC_net), .I3(n50635), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_28 (.CI(n51182), .I0(n2908), 
            .I1(VCC_net), .CO(n51183));
    SB_CARRY encoder0_position_30__I_0_add_833_9 (.CI(n50635), .I0(n1227_adj_5839), 
            .I1(VCC_net), .CO(n50636));
    SB_LUT4 encoder0_position_30__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n51181), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_27 (.CI(n51181), .I0(n2909), 
            .I1(VCC_net), .CO(n51182));
    SB_LUT4 encoder0_position_30__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n51180), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228_adj_5840), 
            .I2(VCC_net), .I3(n50634), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_26 (.CI(n51180), .I0(n2910), 
            .I1(VCC_net), .CO(n51181));
    SB_LUT4 encoder0_position_30__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n51179), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_8 (.CI(n50634), .I0(n1228_adj_5840), 
            .I1(VCC_net), .CO(n50635));
    SB_LUT4 encoder0_position_30__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229_adj_5841), 
            .I2(GND_net), .I3(n50633), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53498_4_lut (.I0(n67525), .I1(n69064), .I2(n70569), .I3(n66980), 
            .O(n69224));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53498_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n57885));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i52527_3_lut (.I0(n67527), .I1(n16_adj_5759), .I2(n68415), 
            .I3(GND_net), .O(n68253));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52527_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53552_4_lut (.I0(n68253), .I1(n69224), .I2(n70569), .I3(n68749), 
            .O(n69278));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53552_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53553_3_lut (.I0(n69278), .I1(duty[18]), .I2(current[15]), 
            .I3(GND_net), .O(n69279));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53553_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53134_4_lut (.I0(n69279), .I1(duty[20]), .I2(current[15]), 
            .I3(duty[19]), .O(n68860));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53134_4_lut.LUT_INIT = 16'h8f0e;
    SB_CARRY encoder0_position_30__I_0_add_1972_25 (.CI(n51179), .I0(n2911), 
            .I1(VCC_net), .CO(n51180));
    SB_CARRY encoder0_position_30__I_0_add_833_7 (.CI(n50633), .I0(n1229_adj_5841), 
            .I1(GND_net), .CO(n50634));
    SB_LUT4 encoder0_position_30__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230_adj_5842), 
            .I2(GND_net), .I3(n50632), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n51178), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1985 (.I0(n18_adj_5862), .I1(n68860), .I2(duty[21]), 
            .I3(current[15]), .O(n6_adj_5936));
    defparam i2_4_lut_adj_1985.LUT_INIT = 16'heafe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n57884));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_833_6 (.CI(n50632), .I0(n1230_adj_5842), 
            .I1(GND_net), .CO(n50633));
    SB_LUT4 encoder0_position_30__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231_adj_5843), 
            .I2(VCC_net), .I3(n50631), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_5 (.CI(n50631), .I0(n1231_adj_5843), 
            .I1(VCC_net), .CO(n50632));
    SB_LUT4 i7_4_lut_adj_1987 (.I0(duty[22]), .I1(duty[23]), .I2(n6_adj_5936), 
            .I3(current[15]), .O(n11573));
    defparam i7_4_lut_adj_1987.LUT_INIT = 16'h3332;
    SB_LUT4 encoder0_position_30__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232_adj_5844), 
            .I2(GND_net), .I3(n50630), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_24 (.CI(n51178), .I0(n2912), 
            .I1(VCC_net), .CO(n51179));
    SB_CARRY encoder0_position_30__I_0_add_833_4 (.CI(n50630), .I0(n1232_adj_5844), 
            .I1(GND_net), .CO(n50631));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n57883));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233_adj_5845), 
            .I2(VCC_net), .I3(n50629), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n51177), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n50303), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_3 (.CI(n50629), .I0(n1233_adj_5845), 
            .I1(VCC_net), .CO(n50630));
    SB_LUT4 encoder0_position_30__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n57882));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n57881));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n57880));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n57879));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n29037));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n57780));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n57781));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_23 (.CI(n51177), .I0(n2913), 
            .I1(VCC_net), .CO(n51178));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n57782));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n57783));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n57878));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n29035));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n29034));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n57877));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n29032));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n57876));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n29030));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n57875));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n57874));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n57873));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n57872));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n57871));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n57870));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2011 (.I0(n2429), .I1(n43025), .I2(n2430), .I3(n2431), 
            .O(n59736));
    defparam i1_4_lut_adj_2011.LUT_INIT = 16'ha080;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n57869));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n57868));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n57867));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n57866));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2016 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n57865));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2016.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n57864));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2018 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n57784));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2018.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2019 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n57785));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2019.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2020 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n57786));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2020.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2021 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n57787));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2021.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n57788));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2023 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n57789));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2023.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2024 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n57790));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2024.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2025 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n57791));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2025.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2026 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n57792));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2026.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2027 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n57793));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2027.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n57794));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2029 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n57795));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2029.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n57796));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2031 (.I0(n2417), .I1(n59736), .I2(n2420), .I3(n62518), 
            .O(n62524));
    defparam i1_4_lut_adj_2031.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n29017));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2033 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n29016));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2033.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2034 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n29015));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2034.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2035 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n57862));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2035.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n57797));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h2300;
    SB_LUT4 i6514_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6514_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2037 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n57733));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2037.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n57798));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h2300;
    SB_LUT4 i6512_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6512_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2039 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n57799));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2039.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2040 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n57800));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2040.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5941), 
            .I2(commutation_state_prev[0]), .I3(dti_N_404), .O(n27624));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2041 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n57801));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2041.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n57802));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5826));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n29013));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n29012));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_adj_2045 (.I0(commutation_state[0]), .I1(n4_adj_5941), 
            .I2(commutation_state_prev[0]), .I3(n42275), .O(n27779));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_2045.LUT_INIT = 16'hffde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n57861));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h2300;
    SB_LUT4 i16245_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30276));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15028_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5941), 
            .I2(commutation_state_prev[0]), .I3(n42275), .O(n29059));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i15028_2_lut_4_lut.LUT_INIT = 16'h00de;
    SB_LUT4 i16254_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30285));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16254_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16748_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n30779));   // verilog/coms.v(130[12] 305[6])
    defparam i16748_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16255_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30286));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16255_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16256_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30287));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16256_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16257_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30288));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16258_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30289));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16260_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30291));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16261_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30292));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2047 (.I0(n244), .I1(Ki[1]), .I2(GND_net), .I3(GND_net), 
            .O(n113));
    defparam i1_2_lut_adj_2047.LUT_INIT = 16'h8888;
    SB_LUT4 i16262_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30293));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1920_3_lut (.I0(n2821_adj_5856), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16263_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n30294));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2048 (.I0(n244), .I1(Ki[2]), .I2(GND_net), .I3(GND_net), 
            .O(n186));
    defparam i1_2_lut_adj_2048.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_2049 (.I0(n244), .I1(Ki[3]), .I2(GND_net), .I3(GND_net), 
            .O(n259));
    defparam i1_2_lut_adj_2049.LUT_INIT = 16'h8888;
    SB_LUT4 i15411_3_lut (.I0(\data_in_frame[0] [5]), .I1(rx_data[5]), .I2(n58008), 
            .I3(GND_net), .O(n29442));   // verilog/coms.v(130[12] 305[6])
    defparam i15411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_2050 (.I0(n25771), .I1(n58169), .I2(\data_in_frame[11] [2]), 
            .I3(n53323), .O(n58561));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_4_lut_adj_2050.LUT_INIT = 16'h6996;
    SB_LUT4 i16747_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n30778));   // verilog/coms.v(130[12] 305[6])
    defparam i16747_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_2051 (.I0(n25771), .I1(n58169), .I2(\data_in_frame[11] [2]), 
            .I3(n25961), .O(Kp_23__N_1301));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_4_lut_adj_2051.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_2052 (.I0(n244), .I1(Ki[4]), .I2(GND_net), .I3(GND_net), 
            .O(n332));
    defparam i1_2_lut_adj_2052.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_2053 (.I0(\data_in_frame[18] [0]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[0]), .O(n57183));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2053.LUT_INIT = 16'h3a0a;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5932));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 encoder0_position_30__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_2054 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42168), .O(n24_adj_5930));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_adj_2054.LUT_INIT = 16'hffbf;
    SB_LUT4 i15382_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n28358), .I3(GND_net), .O(n29413));   // verilog/coms.v(130[12] 305[6])
    defparam i15382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2055 (.I0(n244), .I1(Ki[5]), .I2(GND_net), .I3(GND_net), 
            .O(n405_adj_5857));
    defparam i1_2_lut_adj_2055.LUT_INIT = 16'h8888;
    SB_LUT4 i15379_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n28358), .I3(GND_net), .O(n29410));   // verilog/coms.v(130[12] 305[6])
    defparam i15379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15870_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n58897), 
            .I3(GND_net), .O(n29901));   // verilog/coms.v(130[12] 305[6])
    defparam i15870_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15867_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n58897), 
            .I3(GND_net), .O(n29898));   // verilog/coms.v(130[12] 305[6])
    defparam i15867_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2056 (.I0(n244), .I1(Ki[6]), .I2(GND_net), .I3(GND_net), 
            .O(n478_adj_5846));
    defparam i1_2_lut_adj_2056.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_2057 (.I0(n244), .I1(Ki[7]), .I2(GND_net), .I3(GND_net), 
            .O(n551));
    defparam i1_2_lut_adj_2057.LUT_INIT = 16'h8888;
    SB_LUT4 i15667_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n58009), 
            .I3(GND_net), .O(n29698));   // verilog/coms.v(130[12] 305[6])
    defparam i15667_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2058 (.I0(n244), .I1(Ki[8]), .I2(GND_net), .I3(GND_net), 
            .O(n624));
    defparam i1_2_lut_adj_2058.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_2059 (.I0(n2418), .I1(n2419), .I2(n2422), .I3(GND_net), 
            .O(n62620));
    defparam i1_3_lut_adj_2059.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27722), .O(n53943));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i16358_3_lut_4_lut (.I0(baudrate[9]), .I1(data_adj_6002[1]), 
            .I2(n48949), .I3(n114), .O(n30389));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16358_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i16357_3_lut_4_lut (.I0(baudrate[10]), .I1(data_adj_6002[2]), 
            .I2(n48949), .I3(n114), .O(n30388));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16357_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i16356_3_lut_4_lut (.I0(baudrate[11]), .I1(data_adj_6002[3]), 
            .I2(n48949), .I3(n114), .O(n30387));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16356_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i16355_3_lut_4_lut (.I0(baudrate[12]), .I1(data_adj_6002[4]), 
            .I2(n48949), .I3(n114), .O(n30386));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16355_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i16354_3_lut_4_lut (.I0(baudrate[13]), .I1(data_adj_6002[5]), 
            .I2(n48949), .I3(n114), .O(n30385));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16354_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(reset), .I1(n40525), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n7_adj_5831), .O(n28361));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(reset), .I1(n40525), .I2(n8_adj_5790), 
            .I3(GND_net), .O(n28365));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 mux_245_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_2060 (.I0(reset), .I1(n40525), .I2(n8_adj_5704), 
            .I3(GND_net), .O(n28363));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut_adj_2060.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_2061 (.I0(reset), .I1(n40525), .I2(n8_adj_5779), 
            .I3(GND_net), .O(n28355));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut_adj_2061.LUT_INIT = 16'h0404;
    SB_LUT4 i15373_3_lut (.I0(\data_in_frame[0] [4]), .I1(rx_data[4]), .I2(n58008), 
            .I3(GND_net), .O(n29404));   // verilog/coms.v(130[12] 305[6])
    defparam i15373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16324_3_lut (.I0(current[11]), .I1(data_adj_6010[11]), .I2(n27704), 
            .I3(GND_net), .O(n30355));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16325_3_lut (.I0(current[10]), .I1(data_adj_6010[10]), .I2(n27704), 
            .I3(GND_net), .O(n30356));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16326_3_lut (.I0(current[9]), .I1(data_adj_6010[9]), .I2(n27704), 
            .I3(GND_net), .O(n30357));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16327_3_lut (.I0(current[8]), .I1(data_adj_6010[8]), .I2(n27704), 
            .I3(GND_net), .O(n30358));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16328_3_lut (.I0(current[7]), .I1(data_adj_6010[7]), .I2(n27704), 
            .I3(GND_net), .O(n30359));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16329_3_lut (.I0(current[6]), .I1(data_adj_6010[6]), .I2(n27704), 
            .I3(GND_net), .O(n30360));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16330_3_lut (.I0(current[5]), .I1(data_adj_6010[5]), .I2(n27704), 
            .I3(GND_net), .O(n30361));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16331_3_lut (.I0(current[4]), .I1(data_adj_6010[4]), .I2(n27704), 
            .I3(GND_net), .O(n30362));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16332_3_lut (.I0(current[3]), .I1(data_adj_6010[3]), .I2(n27704), 
            .I3(GND_net), .O(n30363));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16333_3_lut (.I0(current[2]), .I1(data_adj_6010[2]), .I2(n27704), 
            .I3(GND_net), .O(n30364));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16334_3_lut (.I0(current[1]), .I1(data_adj_6010[1]), .I2(n27704), 
            .I3(GND_net), .O(n30365));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16336_3_lut (.I0(baudrate[31]), .I1(data_adj_6002[7]), .I2(n27922), 
            .I3(GND_net), .O(n30367));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16337_3_lut (.I0(baudrate[30]), .I1(data_adj_6002[6]), .I2(n27922), 
            .I3(GND_net), .O(n30368));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16338_3_lut (.I0(baudrate[29]), .I1(data_adj_6002[5]), .I2(n27922), 
            .I3(GND_net), .O(n30369));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16339_3_lut (.I0(baudrate[28]), .I1(data_adj_6002[4]), .I2(n27922), 
            .I3(GND_net), .O(n30370));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16340_3_lut (.I0(baudrate[27]), .I1(data_adj_6002[3]), .I2(n27922), 
            .I3(GND_net), .O(n30371));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16341_3_lut (.I0(baudrate[26]), .I1(data_adj_6002[2]), .I2(n27922), 
            .I3(GND_net), .O(n30372));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16342_3_lut (.I0(baudrate[25]), .I1(data_adj_6002[1]), .I2(n27922), 
            .I3(GND_net), .O(n30373));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6504_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6504_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i16343_3_lut (.I0(baudrate[24]), .I1(data_adj_6002[0]), .I2(n27922), 
            .I3(GND_net), .O(n30374));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6506_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6506_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i6508_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i6508_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i16359_3_lut (.I0(baudrate[8]), .I1(data_adj_6002[0]), .I2(n27924), 
            .I3(GND_net), .O(n30390));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6510_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i6510_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i23046_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), .I3(GND_net), 
            .O(n5));
    defparam i23046_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1587_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n12186));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_2062 (.I0(n62620), .I1(n2415), .I2(n62524), .I3(n2416), 
            .O(n62528));
    defparam i1_4_lut_adj_2062.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5767));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_1587_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n12184));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i23053_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), .I3(GND_net), 
            .O(n10));
    defparam i23053_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5763));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5765));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_4_lut (.I0(n260), .I1(n63531), .I2(duty[23]), .I3(n22_adj_5934), 
            .O(n11571));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h1505;
    SB_LUT4 encoder0_position_30__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5716));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51470_2_lut_4_lut (.I0(duty[10]), .I1(n300), .I2(duty[6]), 
            .I3(n304), .O(n67196));
    defparam i51470_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i15363_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n28358), .I3(GND_net), .O(n29394));   // verilog/coms.v(130[12] 305[6])
    defparam i15363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16537_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n30568));   // verilog/coms.v(130[12] 305[6])
    defparam i16537_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15360_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n28358), .I3(GND_net), .O(n29391));   // verilog/coms.v(130[12] 305[6])
    defparam i15360_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15864_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n58897), 
            .I3(GND_net), .O(n29895));   // verilog/coms.v(130[12] 305[6])
    defparam i15864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_2063 (.I0(\data_in_frame[18] [1]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[1]), .O(n57179));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2063.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15357_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n28358), .I3(GND_net), .O(n29388));   // verilog/coms.v(130[12] 305[6])
    defparam i15357_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5717));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1587_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n12180));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15354_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n28358), .I3(GND_net), .O(n29385));   // verilog/coms.v(130[12] 305[6])
    defparam i15354_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5719));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut_adj_2064 (.I0(\data_in_frame[18] [7]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[7]), .O(n57229));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2064.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2065 (.I0(\data_in_frame[18] [5]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[5]), .O(n57233));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2065.LUT_INIT = 16'h3a0a;
    SB_LUT4 mux_1587_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n12178));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i28235_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i28235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16394_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n20897), .I3(n4_adj_5937), .O(n30425));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i16394_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i15857_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n58897), 
            .I3(GND_net), .O(n29888));   // verilog/coms.v(130[12] 305[6])
    defparam i15857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5827));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut_adj_2066 (.I0(\data_in_frame[18] [4]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[4]), .O(n57235));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2066.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5720));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51045_3_lut (.I0(enable_slow_N_4214), .I1(n11_adj_5773), .I2(state_7__N_4111[0]), 
            .I3(GND_net), .O(n66471));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i51045_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i16_4_lut (.I0(state_adj_6035[0]), .I1(n66471), .I2(n6429), 
            .I3(n42234), .O(n8_adj_5938));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5721));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16398_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[0]), 
            .I2(n10_adj_5729), .I3(n25532), .O(n30429));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16398_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1587_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n12176));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1587_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n12174));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1587_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n12172));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12_4_lut_adj_2067 (.I0(\data_in_frame[18] [3]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[3]), .O(n57237));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2067.LUT_INIT = 16'h3a0a;
    SB_LUT4 i16405_3_lut (.I0(n58988), .I1(r_Bit_Index[0]), .I2(n27845), 
            .I3(GND_net), .O(n30436));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16405_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 mux_1587_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n12170));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i53981_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n62528), 
            .O(n2445));
    defparam i53981_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51397_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n67123));
    defparam i51397_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5707));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2068 (.I0(n2523), .I1(n2527), .I2(n2526), .I3(n2524), 
            .O(n62172));
    defparam i1_4_lut_adj_2068.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2069 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61718), .O(n61724));
    defparam i1_4_lut_adj_2069.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2070 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61724), .O(n61730));
    defparam i1_4_lut_adj_2070.LUT_INIT = 16'hfffe;
    SB_LUT4 i16409_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n61730), 
            .I3(n27), .O(n30440));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16409_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16410_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n58008), 
            .I3(GND_net), .O(n30441));   // verilog/coms.v(130[12] 305[6])
    defparam i16410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16414_4_lut (.I0(CS_MISO_c), .I1(data_adj_6010[0]), .I2(n11_adj_5791), 
            .I3(state_7__N_4320), .O(n30445));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16414_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1587_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n12168));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1587_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n12166));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_3_lut_adj_2071 (.I0(n62172), .I1(n2528), .I2(n2525), .I3(GND_net), 
            .O(n62174));
    defparam i1_3_lut_adj_2071.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_2072 (.I0(n8_adj_5807), .I1(n40525), .I2(GND_net), 
            .I3(GND_net), .O(n28304));
    defparam i1_2_lut_adj_2072.LUT_INIT = 16'hbbbb;
    SB_LUT4 i16421_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n22773), .I3(GND_net), .O(n30452));   // verilog/coms.v(130[12] 305[6])
    defparam i16421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1587_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n12164));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i51628_4_lut (.I0(data_ready), .I1(n6619), .I2(n24_adj_5930), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n66441));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i51628_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i51590_2_lut (.I0(n24_adj_5930), .I1(n6619), .I2(GND_net), 
            .I3(GND_net), .O(n66444));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i51590_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5722));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1587_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n12162));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i49_4_lut (.I0(n66444), .I1(n66441), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5932), .O(n56399));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i16156_4_lut_4_lut (.I0(n27799), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n30187));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16156_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5800));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1587_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n12160));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5801));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1587_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n12158));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1587_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n12156));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5802));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1587_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n12154));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_2_lut (.I0(n187), .I1(n135), .I2(GND_net), .I3(GND_net), 
            .O(n41));
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5828));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1587_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n12152));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i53611_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42168), .I3(GND_net), .O(n27735));
    defparam i53611_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 mux_1587_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n12150));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1587_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5811));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51682_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n66302));
    defparam i51682_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i28365_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42168), .I3(GND_net), .O(n42285));
    defparam i28365_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut (.I0(state[0]), .I1(bit_ctr[4]), .I2(n42981), 
            .I3(GND_net), .O(n4_adj_5926));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd5d5;
    SB_LUT4 i28355_2_lut (.I0(n22841), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n42275));
    defparam i28355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_2073 (.I0(hall2), .I1(commutation_state_7__N_27[2]), 
            .I2(GND_net), .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_adj_2073.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut_adj_2074 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_2074.LUT_INIT = 16'h1414;
    SB_LUT4 i16530_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n30561));   // verilog/coms.v(130[12] 305[6])
    defparam i16530_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54394_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5942));
    defparam i54394_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 i29168_4_lut (.I0(n950), .I1(n2531), .I2(n2532), .I3(n2533), 
            .O(n43095));
    defparam i29168_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1858_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42168), .O(n6619));   // verilog/TinyFPGA_B.v(362[5] 388[12])
    defparam i1858_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(reset), .I1(rx_data[2]), .I2(\data_in_frame[1] [2]), 
            .I3(n28338), .O(n57383));   // verilog/coms.v(94[13:20])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hf0e4;
    SB_LUT4 i14767_2_lut (.I0(n27648), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28804));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14767_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_2075 (.I0(n2519), .I1(n2520), .I2(n62174), .I3(n2521), 
            .O(n62180));
    defparam i1_4_lut_adj_2075.LUT_INIT = 16'hfffe;
    SB_LUT4 i53554_4_lut (.I0(commutation_state[1]), .I1(n22841), .I2(dti), 
            .I3(commutation_state[2]), .O(n27648));
    defparam i53554_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i1_4_lut_adj_2076 (.I0(n2529), .I1(n62180), .I2(n43095), .I3(n2530), 
            .O(n62182));
    defparam i1_4_lut_adj_2076.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2077 (.I0(n2516), .I1(n2515), .I2(n2518), .I3(n2522), 
            .O(n61008));
    defparam i1_4_lut_adj_2077.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2078 (.I0(n61008), .I1(n2514), .I2(n2517), .I3(n62182), 
            .O(n62188));
    defparam i1_4_lut_adj_2078.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_4306_i24_3_lut (.I0(encoder0_position[23]), .I1(n9_adj_5750), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n934));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231_adj_5843));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i842_3_lut (.I0(n1231_adj_5843), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2079 (.I0(\data_in_frame[8] [6]), .I1(n26306), 
            .I2(GND_net), .I3(GND_net), .O(n58169));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_2079.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54074_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n62188), 
            .O(n2544));
    defparam i54074_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_2080 (.I0(hall1), .I1(hall2), .I2(n20897), 
            .I3(GND_net), .O(n4_adj_5937));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_2080.LUT_INIT = 16'hf2f2;
    SB_LUT4 encoder0_position_30__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2081 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n57860));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2081.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2082 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n57859));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2082.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2083 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n57858));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2083.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2084 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n57857));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2084.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2085 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n57900));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2085.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2086 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n57856));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2086.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2087 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n57863));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2087.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2088 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n57855));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2088.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2089 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n57854));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2089.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2090 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n57853));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2090.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5829));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2091 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n57852));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2091.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36293_3_lut_4_lut (.I0(n37050), .I1(Ki[2]), .I2(n50204), 
            .I3(n20194), .O(n4_adj_5918));
    defparam i36293_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut (.I0(n37050), .I1(Ki[2]), .I2(n50204), .I3(n20194), 
            .O(n20185));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2092 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n57851));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2092.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2093 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n57850));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2093.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2094 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n28997));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2094.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2095 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n57849));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2095.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2096 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n57848));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2096.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2097 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n57847));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2097.LUT_INIT = 16'h2300;
    SB_LUT4 i29166_4_lut (.I0(n951), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n43093));
    defparam i29166_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i36117_3_lut_4_lut (.I0(n37154), .I1(Ki[3]), .I2(n4_adj_5915), 
            .I3(n20158), .O(n6_adj_5916));
    defparam i36117_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 encoder0_position_30__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_2098 (.I0(control_mode[1]), .I1(control_mode[0]), 
            .I2(n37407), .I3(GND_net), .O(n15_adj_5806));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_3_lut_adj_2098.LUT_INIT = 16'hfdfd;
    SB_LUT4 encoder0_position_30__I_0_i1773_3_lut (.I0(n2610), .I1(n2677), 
            .I2(n2643), .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2099 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n57846));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2099.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2100 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n57845));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2100.LUT_INIT = 16'h2300;
    SB_LUT4 i43128_3_lut (.I0(n3), .I1(n7445), .I2(n58792), .I3(GND_net), 
            .O(n58793));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43129_3_lut (.I0(encoder0_position[29]), .I1(n58793), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_2101 (.I0(n37154), .I1(Ki[3]), .I2(n4_adj_5915), 
            .I3(n20158), .O(n20112));
    defparam i1_3_lut_4_lut_adj_2101.LUT_INIT = 16'h8778;
    SB_LUT4 encoder0_position_30__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2102 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n57844));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2102.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225_adj_5837));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i836_3_lut (.I0(n1225_adj_5837), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2103 (.I0(n2619), .I1(n2627), .I2(n2625), .I3(n2623), 
            .O(n62554));
    defparam i1_4_lut_adj_2103.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2104 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n57843));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2104.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2105 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n57842));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2105.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2106 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n28988));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2106.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2107 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n57841));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2107.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2108 (.I0(n2629), .I1(n62554), .I2(n43093), .I3(n2630), 
            .O(n62556));
    defparam i1_4_lut_adj_2108.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_4_lut_adj_2109 (.I0(n37154), .I1(Ki[2]), .I2(n50001), 
            .I3(n20159), .O(n20113));
    defparam i1_3_lut_4_lut_adj_2109.LUT_INIT = 16'h8778;
    SB_LUT4 encoder0_position_30__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36109_3_lut_4_lut (.I0(n37154), .I1(Ki[2]), .I2(n50001), 
            .I3(n20159), .O(n4_adj_5915));
    defparam i36109_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2110 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n57840));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2110.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2111 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n57839));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2111.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2112 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n57838));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2112.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2113 (.I0(n2615), .I1(n2616), .I2(n2617), .I3(n62556), 
            .O(n62562));
    defparam i1_4_lut_adj_2113.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1840_3_lut (.I0(n2709), .I1(n2776), 
            .I2(n2742), .I3(GND_net), .O(n2808));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i18_3_lut (.I0(encoder0_position[17]), .I1(n15_adj_5743), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2114 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n57837));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2114.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2115 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n57836));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2115.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2116 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n57835));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2116.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43136_3_lut (.I0(n7_adj_5752), .I1(n7449), .I2(n58792), .I3(GND_net), 
            .O(n58801));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2117 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n57834));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2117.LUT_INIT = 16'h2300;
    SB_LUT4 i43137_3_lut (.I0(encoder0_position[25]), .I1(n58801), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2118 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n57833));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2118.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2119 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n57832));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2119.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2120 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n57831));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2120.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_2121 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n57927));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_2121.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_2122 (.I0(n2624), .I1(n2621), .I2(GND_net), .I3(GND_net), 
            .O(n62540));
    defparam i1_2_lut_adj_2122.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_2123 (.I0(n2626), .I1(n2622), .I2(n2628), .I3(GND_net), 
            .O(n62542));
    defparam i1_3_lut_adj_2123.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2124 (.I0(n2612), .I1(n2613), .I2(n2614), .I3(n62562), 
            .O(n62568));
    defparam i1_4_lut_adj_2124.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229_adj_5841));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2125 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n57830));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2125.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2126 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n57829));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2126.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i840_3_lut (.I0(n1229_adj_5841), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_4_lut_adj_2127 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n42168), .O(n56483));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_4_lut_4_lut_adj_2127.LUT_INIT = 16'hb1f1;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2128 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n57828));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2128.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2129 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61798), .O(n61804));
    defparam i1_4_lut_adj_2129.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2130 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61804), .O(n61810));
    defparam i1_4_lut_adj_2130.LUT_INIT = 16'hfffe;
    SB_LUT4 i15526_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n61810), 
            .I3(n27), .O(n29557));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15526_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2131 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61782), .O(n61788));
    defparam i1_4_lut_adj_2131.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2132 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61788), .O(n61794));
    defparam i1_4_lut_adj_2132.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2133 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n57827));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2133.LUT_INIT = 16'h2300;
    SB_LUT4 i15527_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n61794), 
            .I3(n27), .O(n29558));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15527_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2134 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n57826));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2134.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2135 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n57825));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2135.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2136 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n57824));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2136.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2137 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n57823));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2137.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2138 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61766), .O(n61772));
    defparam i1_4_lut_adj_2138.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2139 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61772), .O(n61778));
    defparam i1_4_lut_adj_2139.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2140 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n57822));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2140.LUT_INIT = 16'h2300;
    SB_LUT4 i15528_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n61778), 
            .I3(n27), .O(n29559));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15528_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2141 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61814), .O(n61820));
    defparam i1_4_lut_adj_2141.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2142 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61820), .O(n61826));
    defparam i1_4_lut_adj_2142.LUT_INIT = 16'hfffe;
    SB_LUT4 i15559_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n61826), 
            .I3(n27), .O(n29590));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15559_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2143 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n57821));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2143.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2144 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n57820));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2144.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2145 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61734), .O(n61740));
    defparam i1_4_lut_adj_2145.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2146 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61740), .O(n61746));
    defparam i1_4_lut_adj_2146.LUT_INIT = 16'hfffe;
    SB_LUT4 i15560_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n61746), 
            .I3(n27), .O(n29591));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15560_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2147 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61750), .O(n61756));
    defparam i1_4_lut_adj_2147.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2148 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61756), .O(n61762));
    defparam i1_4_lut_adj_2148.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15564_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n61762), 
            .I3(n27), .O(n29595));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15564_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2149 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n57819));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2149.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2150 (.I0(o_Rx_DV_N_3488[12]), .I1(n4939), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n61702), .O(n61708));
    defparam i1_4_lut_adj_2150.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2151 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5728), 
            .I3(n61708), .O(n61714));
    defparam i1_4_lut_adj_2151.LUT_INIT = 16'hfffe;
    SB_LUT4 i15565_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n61714), 
            .I3(n27), .O(n29596));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15565_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2152 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n57818));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2152.LUT_INIT = 16'h2300;
    SB_LUT4 i15584_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n22760), .I3(GND_net), .O(n29615));   // verilog/coms.v(130[12] 305[6])
    defparam i15584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23050_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n22773), .I3(GND_net), .O(n29617));
    defparam i23050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2153 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n57817));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2153.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2154 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n57734));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2154.LUT_INIT = 16'h2300;
    SB_LUT4 i15676_3_lut_4_lut (.I0(n1742), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3837), .O(n29707));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15676_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i43134_3_lut (.I0(n6_adj_5753), .I1(n7448), .I2(n58792), .I3(GND_net), 
            .O(n58799));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43135_3_lut (.I0(encoder0_position[26]), .I1(n58799), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228_adj_5840));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2155 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n57816));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2155.LUT_INIT = 16'h2300;
    SB_LUT4 i15671_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29702));   // verilog/coms.v(130[12] 305[6])
    defparam i15671_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i839_3_lut (.I0(n1228_adj_5840), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2156 (.I0(n2618), .I1(n62542), .I2(n2620), .I3(n62540), 
            .O(n62548));
    defparam i1_4_lut_adj_2156.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2157 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n28960));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2157.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1174_3_lut (.I0(n1723), .I1(n1790_adj_5848), 
            .I2(n1752), .I3(GND_net), .O(n1822_adj_5852));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5830));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1241_3_lut (.I0(n1822_adj_5852), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2158 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n57815));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2158.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5833));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_4_lut_adj_2159 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2821), .O(n25_adj_5928));   // verilog/TinyFPGA_B.v(377[7:11])
    defparam i1_4_lut_4_lut_adj_2159.LUT_INIT = 16'h5450;
    SB_LUT4 mux_4306_i26_3_lut (.I0(encoder0_position[25]), .I1(n7_adj_5752), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2160 (.I0(n4_adj_5776), .I1(n5_adj_5775), .I2(n731), 
            .I3(n6_adj_5753), .O(n5_adj_5929));
    defparam i1_4_lut_adj_2160.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_2161 (.I0(n3), .I1(n2_adj_5778), .I2(n5_adj_5929), 
            .I3(GND_net), .O(n58792));
    defparam i1_3_lut_adj_2161.LUT_INIT = 16'h8080;
    SB_LUT4 i43132_3_lut (.I0(n5_adj_5775), .I1(n7447), .I2(n58792), .I3(GND_net), 
            .O(n58797));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43133_3_lut (.I0(encoder0_position[27]), .I1(n58797), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i43133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47939_3_lut (.I0(n4910), .I1(duty[20]), .I2(n11573), .I3(GND_net), 
            .O(n63665));
    defparam i47939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47941_3_lut (.I0(n63665), .I1(n63663), .I2(n11571), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i47941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227_adj_5839));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i838_3_lut (.I0(n1227_adj_5839), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2162 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n57814));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2162.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2163 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n57813));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2163.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i25_3_lut (.I0(encoder0_position[24]), .I1(n8_adj_5751), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15594_3_lut (.I0(current[0]), .I1(data_adj_6010[0]), .I2(n27704), 
            .I3(GND_net), .O(n29625));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47936_3_lut (.I0(n4909), .I1(duty[21]), .I2(n11573), .I3(GND_net), 
            .O(n63662));
    defparam i47936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230_adj_5842));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i841_3_lut (.I0(n1230_adj_5842), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47938_3_lut (.I0(n63662), .I1(n63663), .I2(n11571), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i47938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1176_3_lut (.I0(n1725), .I1(n1792_adj_5849), 
            .I2(n1752), .I3(GND_net), .O(n1824_adj_5853));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47937_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n11573), 
            .I3(GND_net), .O(n63663));
    defparam i47937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47933_3_lut (.I0(n4908), .I1(duty[22]), .I2(n11573), .I3(GND_net), 
            .O(n63659));
    defparam i47933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47935_3_lut (.I0(n63659), .I1(n63663), .I2(n11571), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i47935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1243_3_lut (.I0(n1824_adj_5853), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7219_3_lut (.I0(n4907), .I1(current[15]), .I2(n11571), .I3(GND_net), 
            .O(n20935));
    defparam i7219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7220_3_lut (.I0(n20935), .I1(duty[23]), .I2(n11573), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i7220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2164 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n57812));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2164.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_4306_i10_3_lut (.I0(encoder0_position[9]), .I1(n23_adj_5735), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i9_3_lut (.I0(encoder0_position[8]), .I1(n24_adj_5734), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i8_3_lut (.I0(encoder0_position[7]), .I1(n25_adj_5733), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5914));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i23_3_lut (.I0(encoder0_position[22]), .I1(n10_adj_5748), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n935));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i709_3_lut (.I0(n935), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5913));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2165 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n57811));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2165.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232_adj_5844));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i843_3_lut (.I0(n1232_adj_5844), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1178_3_lut (.I0(n1727), .I1(n1794_adj_5850), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(0)  quad_counter1 (.a_prev(a_prev_adj_5782), .b_prev(b_prev_adj_5783), 
            .a_new({a_new_adj_5988[1], Open_0}), .b_new({b_new_adj_5989[1], 
            Open_1}), .position_31__N_3837(position_31__N_3837_adj_5785), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1779(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .n1786(n1786), .GND_net(GND_net), .n1788(n1788), .n1790(n1790), 
            .n1792(n1792), .n1794(n1794), .n1796(n1796), .\encoder1_position[25] (encoder1_position[25]), 
            .\encoder1_position[24] (encoder1_position[24]), .\encoder1_position[23] (encoder1_position[23]), 
            .\encoder1_position[22] (encoder1_position[22]), .\encoder1_position[21] (encoder1_position[21]), 
            .\encoder1_position[20] (encoder1_position[20]), .\encoder1_position[19] (encoder1_position[19]), 
            .\encoder1_position[18] (encoder1_position[18]), .\encoder1_position[17] (encoder1_position[17]), 
            .\encoder1_position[16] (encoder1_position[16]), .\encoder1_position[15] (encoder1_position[15]), 
            .\encoder1_position[14] (encoder1_position[14]), .\encoder1_position[13] (encoder1_position[13]), 
            .\encoder1_position[12] (encoder1_position[12]), .\encoder1_position[11] (encoder1_position[11]), 
            .\encoder1_position[10] (encoder1_position[10]), .\encoder1_position[9] (encoder1_position[9]), 
            .\encoder1_position[8] (encoder1_position[8]), .\encoder1_position[7] (encoder1_position[7]), 
            .\encoder1_position[6] (encoder1_position[6]), .\encoder1_position[5] (encoder1_position[5]), 
            .\encoder1_position[4] (encoder1_position[4]), .n29664(n29664), 
            .n1784(n1784), .\encoder1_position[3] (encoder1_position[3]), 
            .n29656(n29656), .\encoder1_position[2] (encoder1_position[2]), 
            .n1822(n1822), .n1824(n1824), .VCC_net(VCC_net), .n29397(n29397), 
            .debounce_cnt_N_3834(debounce_cnt_N_3834_adj_5784)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 encoder0_position_30__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i22_3_lut (.I0(encoder0_position[21]), .I1(n11_adj_5747), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n936));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233_adj_5845));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i844_3_lut (.I0(n1233_adj_5845), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5912));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28234_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i28234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28360_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i28360_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2166 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n57810));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2166.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5803));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2167 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n57809));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2167.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(\data_out_frame[9] [0]), .O(n10_adj_5726));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2168 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n57808));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2168.LUT_INIT = 16'h2300;
    SB_LUT4 i15599_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n22773), .I3(GND_net), .O(n29630));   // verilog/coms.v(130[12] 305[6])
    defparam i15599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2169 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n57807));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2169.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2170 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n57806));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2170.LUT_INIT = 16'h2300;
    SB_LUT4 mux_4306_i19_3_lut (.I0(encoder0_position[18]), .I1(n14_adj_5744), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5804));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5805));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2171 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n57805));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2171.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i16_3_lut (.I0(encoder0_position[15]), .I1(n17_adj_5741), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.clk16MHz(clk16MHz), .enable_slow_N_4214(enable_slow_N_4214), 
           .GND_net(GND_net), .\state[0] (state_adj_6035[0]), .\state_7__N_3919[0] (state_7__N_3919[0]), 
           .data_ready(data_ready), .ID({ID}), .baudrate({baudrate}), 
           .n30390(n30390), .n30389(n30389), .n30388(n30388), .n30387(n30387), 
           .n30386(n30386), .n30385(n30385), .n30374(n30374), .n30373(n30373), 
           .n30372(n30372), .n30371(n30371), .n30370(n30370), .n30369(n30369), 
           .n30368(n30368), .n30367(n30367), .n114(n114), .data({data_adj_6002}), 
           .n27922(n27922), .n48949(n48949), .n27924(n27924), .\state_7__N_4111[0] (state_7__N_4111[0]), 
           .scl_enable(scl_enable), .VCC_net(VCC_net), .sda_enable(sda_enable), 
           .sda_out(sda_out), .n29653(n29653), .n29652(n29652), .n29646(n29646), 
           .n29645(n29645), .n29640(n29640), .n29639(n29639), .n29637(n29637), 
           .n6429(n6429), .n30429(n30429), .n8(n8_adj_5938), .n11(n11_adj_5773), 
           .scl(scl), .n42234(n42234), .\state_7__N_4127[3] (state_7__N_4127[3]), 
           .n10(n10_adj_5729), .n4(n4_adj_5771), .n4_adj_26(n4_adj_5772), 
           .n25532(n25532), .n25568(n25568), .n42355(n42355)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(391[10] 403[6])
    SB_LUT4 i3_4_lut_adj_2172 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n61190));
    defparam i3_4_lut_adj_2172.LUT_INIT = 16'h0004;
    SB_LUT4 encoder0_position_30__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15606_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[1]), 
            .I2(n10_adj_5729), .I3(n25568), .O(n29637));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15606_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15608_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[2]), 
            .I2(n4_adj_5771), .I3(n25532), .O(n29639));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15608_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2173 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n57804));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2173.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15609_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[3]), 
            .I2(n4_adj_5771), .I3(n25568), .O(n29640));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i13_3_lut (.I0(encoder0_position[12]), .I1(n20_adj_5738), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54043_4_lut (.I0(n2610), .I1(n62548), .I2(n62568), .I3(n2611), 
            .O(n2643));
    defparam i54043_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i20_3_lut (.I0(encoder0_position[19]), .I1(n13_adj_5745), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n938));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15633_3_lut_4_lut (.I0(n1784), .I1(b_prev_adj_5783), .I2(a_new_adj_5988[1]), 
            .I3(position_31__N_3837_adj_5785), .O(n29664));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15633_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i15613_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n31_adj_5935), .I3(GND_net), .O(n29644));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15613_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15614_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[4]), 
            .I2(n4_adj_5772), .I3(n25532), .O(n29645));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15614_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15615_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[5]), 
            .I2(n4_adj_5772), .I3(n25568), .O(n29646));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15615_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5810), .I3(n15_adj_5806), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i7_3_lut (.I0(encoder0_position[6]), .I1(n26_adj_5732), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i6_3_lut (.I0(encoder0_position[5]), .I1(n27_adj_5731), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2174 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n57803));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2174.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i5_3_lut (.I0(encoder0_position[4]), .I1(n28), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_4306_i12_3_lut (.I0(encoder0_position[11]), .I1(n21_adj_5737), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15619_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n22760), .I3(GND_net), .O(n29650));   // verilog/coms.v(130[12] 305[6])
    defparam i15619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5911));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i17_3_lut (.I0(encoder0_position[16]), .I1(n16_adj_5742), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15620_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n22760), .I3(GND_net), .O(n29651));   // verilog/coms.v(130[12] 305[6])
    defparam i15620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2175 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n57735));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2175.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2176 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n57736));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2176.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15621_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[6]), 
            .I2(n42355), .I3(n25532), .O(n29652));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15621_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53741_1_lut (.I0(n43071), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69467));
    defparam i53741_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2177 (.I0(n3217), .I1(n29_adj_5924), .I2(n3284), 
            .I3(n3237), .O(n62218));
    defparam i1_4_lut_adj_2177.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2178 (.I0(n3216), .I1(n62218), .I2(n3283), .I3(n3237), 
            .O(n62220));
    defparam i1_4_lut_adj_2178.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2179 (.I0(n3213), .I1(n62220), .I2(n3280), .I3(n3237), 
            .O(n62222));
    defparam i1_4_lut_adj_2179.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2180 (.I0(n3212), .I1(n62222), .I2(n3279), .I3(n3237), 
            .O(n62224));
    defparam i1_4_lut_adj_2180.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2190_3_lut (.I0(n3219), .I1(n3286), 
            .I2(n3237), .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2181 (.I0(n15_adj_5920), .I1(n19_adj_5922), .I2(n13_adj_5919), 
            .I3(n33), .O(n62380));
    defparam i1_4_lut_adj_2181.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2182 (.I0(n3215), .I1(n62380), .I2(n3282), .I3(n3237), 
            .O(n62382));
    defparam i1_4_lut_adj_2182.LUT_INIT = 16'heefc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2183 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n57737));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2183.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2184 (.I0(n3211), .I1(n62382), .I2(n3278), .I3(n3237), 
            .O(n62384));
    defparam i1_4_lut_adj_2184.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2185 (.I0(n3209), .I1(n62384), .I2(n3276), .I3(n3237), 
            .O(n62386));
    defparam i1_4_lut_adj_2185.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2186 (.I0(n3223), .I1(n31_adj_5925), .I2(n3290), 
            .I3(n3237), .O(n62330));
    defparam i1_4_lut_adj_2186.LUT_INIT = 16'heefc;
    SB_LUT4 i16_4_lut_adj_2187 (.I0(n3231), .I1(n66396), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5869));
    defparam i16_4_lut_adj_2187.LUT_INIT = 16'hac0c;
    coms neopxl_color_23__I_0 (.n29606(n29606), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .clk16MHz(clk16MHz), .n29891(n29891), .VCC_net(VCC_net), .\data_in_frame[7] ({Open_2, 
         Open_3, \data_in_frame[7] [5:0]}), .GND_net(GND_net), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .n29888(n29888), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n2874(n2874), .\data_out_frame[8] ({\data_out_frame[8] }), .n57860(n57860), 
         .n57859(n57859), .n29885(n29885), .\data_in_frame[8] ({Open_4, 
         Open_5, Open_6, \data_in_frame[8] [4], Open_7, \data_in_frame[8] [2], 
         Open_8, Open_9}), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .n58651(n58651), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .n58570(n58570), .n25705(n25705), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), .pwm_setpoint({pwm_setpoint}), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .current_limit({Open_10, Open_11, Open_12, Open_13, Open_14, 
         current_limit[10], Open_15, Open_16, Open_17, current_limit[6], 
         Open_18, Open_19, Open_20, Open_21, Open_22, Open_23}), 
         .n22773(n22773), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .n58099(n58099), .\data_out_frame[4] ({\data_out_frame[4] }), .n25676(n25676), 
         .n29881(n29881), .n29878(n29878), .n29875(n29875), .n29872(n29872), 
         .n29869(n29869), .n29866(n29866), .n29863(n29863), .n29860(n29860), 
         .n29857(n29857), .\data_in_frame[5] ({\data_in_frame[5] }), .n29854(n29854), 
         .n29851(n29851), .n29848(n29848), .n29621(n29621), .n29844(n29844), 
         .\data_in_frame[0] ({Open_24, Open_25, Open_26, Open_27, \data_in_frame[0] [3:1], 
         Open_28}), .n29841(n29841), .n29838(n29838), .n26306(n26306), 
         .n29818(n29818), .n25666(n25666), .n34(n34), .\data_in_frame[0][5] (\data_in_frame[0] [5]), 
         .n26111(n26111), .n2076(n2076), .encoder1_position_scaled({encoder1_position_scaled}), 
         .displacement({displacement}), .n15(n15_adj_5810), .n15_adj_7(n15_adj_5806), 
         .\data_in_frame[3] ({Open_29, Open_30, Open_31, Open_32, \data_in_frame[3] [3], 
         Open_33, \data_in_frame[3] [1], Open_34}), .\data_in_frame[2][1] (\data_in_frame[2] [1]), 
         .\data_in_frame[0][0] (\data_in_frame[0] [0]), .\data_in_frame[2][5] (\data_in_frame[2] [5]), 
         .\data_in_frame[3][0] (\data_in_frame[3] [0]), .n58498(n58498), 
         .\data_in_frame[1] ({Open_35, Open_36, \data_in_frame[1] [5], 
         Open_37, Open_38, Open_39, Open_40, Open_41}), .\data_in_frame[3][7] (\data_in_frame[3] [7]), 
         .n29641(n29641), .neopxl_color({neopxl_color}), .n29657(n29657), 
         .n58075(n58075), .encoder0_position_scaled({encoder0_position_scaled}), 
         .\data_in_frame[1][6] (\data_in_frame[1] [6]), .n29813(n29813), 
         .n57858(n57858), .\data_in_frame[1][7] (\data_in_frame[1] [7]), 
         .\data_in_frame[8][3] (\data_in_frame[8] [3]), .n57857(n57857), 
         .reset(reset), .setpoint({setpoint}), .\data_in_frame[1][2] (\data_in_frame[1] [2]), 
         .deadband({deadband}), .\data_in_frame[2][0] (\data_in_frame[2] [0]), 
         .\data_in_frame[3][5] (\data_in_frame[3] [5]), .n29698(n29698), 
         .\data_in_frame[2][3] (\data_in_frame[2] [3]), .n57900(n57900), 
         .control_mode({control_mode[7:5], Open_42, Open_43, Open_44, 
         Open_45, Open_46}), .n57856(n57856), .\data_in_frame[8][6] (\data_in_frame[8] [6]), 
         .\control_mode[1] (control_mode[1]), .\data_in_frame[20][4] (\data_in_frame[20] [4]), 
         .\control_mode[0] (control_mode[0]), .\data_in_frame[21][2] (\data_in_frame[21] [2]), 
         .\data_in_frame[21][3] (\data_in_frame[21] [3]), .\data_in_frame[18] ({Open_47, 
         Open_48, \data_in_frame[18] [5], Open_49, Open_50, Open_51, 
         Open_52, Open_53}), .n57863(n57863), .n57855(n57855), .n57854(n57854), 
         .n57853(n57853), .n57852(n57852), .n57851(n57851), .n57850(n57850), 
         .n28997(n28997), .n57849(n57849), .n57848(n57848), .n57847(n57847), 
         .n57846(n57846), .n57845(n57845), .n57844(n57844), .n57843(n57843), 
         .n57842(n57842), .\data_in_frame[22][5] (\data_in_frame[22] [5]), 
         .\data_in_frame[20][3] (\data_in_frame[20] [3]), .\data_in_frame[22][4] (\data_in_frame[22] [4]), 
         .\data_in_frame[20][0] (\data_in_frame[20] [0]), .\data_in_frame[21][1] (\data_in_frame[21] [1]), 
         .\data_in_frame[21][5] (\data_in_frame[21] [5]), .\data_in_frame[19] ({\data_in_frame[19] [7:6], 
         Open_54, Open_55, \data_in_frame[19] [3:0]}), .\data_in_frame[22][1] (\data_in_frame[22] [1]), 
         .n28988(n28988), .n57841(n57841), .n57840(n57840), .n57839(n57839), 
         .n57838(n57838), .n57837(n57837), .n57836(n57836), .n57835(n57835), 
         .\data_in_frame[22][7] (\data_in_frame[22] [7]), .n57834(n57834), 
         .n57833(n57833), .n57832(n57832), .n57831(n57831), .n57830(n57830), 
         .n57829(n57829), .n57828(n57828), .\data_in_frame[17] ({\data_in_frame[17] [7], 
         Open_56, Open_57, Open_58, Open_59, Open_60, Open_61, \data_in_frame[17] [0]}), 
         .\data_in_frame[22][2] (\data_in_frame[22] [2]), .n57827(n57827), 
         .\data_in_frame[20][1] (\data_in_frame[20] [1]), .\data_in_frame[22][3] (\data_in_frame[22] [3]), 
         .n57826(n57826), .n57825(n57825), .n57824(n57824), .n57823(n57823), 
         .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .n4942(n4942), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
         .n29(n29), .n23(n23_adj_5728), .n27(n27), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
         .n57822(n57822), .n57821(n57821), .n57820(n57820), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .n37407(n37407), .n57819(n57819), .n57818(n57818), .n57817(n57817), 
         .n57734(n57734), .n57816(n57816), .n28960(n28960), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .\data_out_frame[3][1] (\data_out_frame[3] [1]), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .n57815(n57815), .n29703(n29703), .n57814(n57814), .IntegralLimit({IntegralLimit}), 
         .n57813(n57813), .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), .ID({ID}), 
         .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), 
         .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), 
         .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), 
         .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .n29709(n29709), .\Kp[15] (Kp[15]), 
         .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), 
         .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .n8(n8_adj_5790), 
         .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), 
         .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
         .n29729(n29729), .n29728(n29728), .n29727(n29727), .n29726(n29726), 
         .n29725(n29725), .n29724(n29724), .n29723(n29723), .n29722(n29722), 
         .n29721(n29721), .n29720(n29720), .n150(n150), .n36515(n36515), 
         .n29719(n29719), .n29718(n29718), .n29717(n29717), .n29716(n29716), 
         .n29715(n29715), .n29714(n29714), .n58897(n58897), .n29713(n29713), 
         .n29712(n29712), .n29708(n29708), .n29702(n29702), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n29701(n29701), 
         .n29697(n29697), .\current_limit[2] (current_limit[2]), .\data_out_frame[3][6] (\data_out_frame[3] [6]), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .PWMLimit({PWMLimit}), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .n57812(n57812), 
         .n57811(n57811), .n57810(n57810), .n57809(n57809), .rx_data({rx_data}), 
         .n58929(n58929), .n57808(n57808), .n57807(n57807), .n57806(n57806), 
         .n57805(n57805), .n29677(n29677), .\current_limit[12] (current_limit[12]), 
         .n57804(n57804), .n57803(n57803), .n29676(n29676), .\current_limit[11] (current_limit[11]), 
         .n29674(n29674), .\current_limit[9] (current_limit[9]), .n29673(n29673), 
         .\current_limit[8] (current_limit[8]), .n29671(n29671), .\current_limit[7] (current_limit[7]), 
         .n57735(n57735), .n57736(n57736), .n57737(n57737), .n57738(n57738), 
         .n29669(n29669), .\current_limit[5] (current_limit[5]), .n57739(n57739), 
         .n29666(n29666), .\current_limit[3] (current_limit[3]), .n57740(n57740), 
         .\data_out_frame[1][7] (\data_out_frame[1] [7]), .n28940(n28940), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .n29655(n29655), 
         .n29654(n29654), .n57741(n57741), .n57742(n57742), .n57743(n57743), 
         .n29651(n29651), .n29650(n29650), .n57744(n57744), .n57745(n57745), 
         .n29630(n29630), .n7(n7_adj_5939), .n57746(n57746), .n57747(n57747), 
         .n30552(n30552), .n28932(n28932), .n57748(n57748), .n8_adj_8(n8_adj_5704), 
         .n29617(n29617), .\current_limit[0] (current_limit[0]), .n29615(n29615), 
         .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n57749(n57749), .n57750(n57750), 
         .n57751(n57751), .n57752(n57752), .n57753(n57753), .n57754(n57754), 
         .n30561(n30561), .n28924(n28924), .n57755(n57755), .n57756(n57756), 
         .n57757(n57757), .n57758(n57758), .n57759(n57759), .n57760(n57760), 
         .n30568(n30568), .n28917(n28917), .n41(n41_adj_5917), .n57761(n57761), 
         .n57762(n57762), .n57763(n57763), .n25(n25_adj_5724), .n28911(n28911), 
         .n28910(n28910), .n57764(n57764), .n57765(n57765), .n57766(n57766), 
         .n57767(n57767), .n57768(n57768), .n57769(n57769), .n57770(n57770), 
         .n57771(n57771), .n57772(n57772), .n57773(n57773), .n57774(n57774), 
         .n57775(n57775), .n57776(n57776), .n57777(n57777), .n57778(n57778), 
         .n57779(n57779), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n28893(n28893), .rx_data_ready(rx_data_ready), .n57899(n57899), 
         .\data_out_frame[0][3] (\data_out_frame[0] [3]), .n57898(n57898), 
         .n58008(n58008), .n30452(n30452), .\current_limit[4] (current_limit[4]), 
         .n30441(n30441), .n57237(n57237), .\data_in_frame[18][3] (\data_in_frame[18] [3]), 
         .n57235(n57235), .\data_in_frame[18][4] (\data_in_frame[18] [4]), 
         .n57233(n57233), .n8_adj_9(n8_adj_5779), .n58010(n58010), .n57229(n57229), 
         .\data_in_frame[18][7] (\data_in_frame[18] [7]), .n29385(n29385), 
         .n29388(n29388), .n57179(n57179), .\data_in_frame[18][1] (\data_in_frame[18] [1]), 
         .n29895(n29895), .n29391(n29391), .n29394(n29394), .n29404(n29404), 
         .\data_in_frame[0][4] (\data_in_frame[0] [4]), .n29898(n29898), 
         .n29901(n29901), .n29410(n29410), .n29413(n29413), .n57183(n57183), 
         .\data_in_frame[18][0] (\data_in_frame[18] [0]), .n29442(n29442), 
         .n57383(n57383), .\data_in_frame[9][7] (\data_in_frame[9] [7]), 
         .\data_in_frame[11][2] (\data_in_frame[11] [2]), .\data_in_frame[12] ({Open_62, 
         Open_63, Open_64, Open_65, Open_66, Open_67, Open_68, \data_in_frame[12] [0]}), 
         .\data_out_frame[1][5] (\data_out_frame[1] [5]), .n58011(n58011), 
         .n57225(n57225), .\data_in_frame[16] ({\data_in_frame[16] }), .n57223(n57223), 
         .n57221(n57221), .n57219(n57219), .n57215(n57215), .n57211(n57211), 
         .n57207(n57207), .n57203(n57203), .n30149(n30149), .n58009(n58009), 
         .n57199(n57199), .\data_in_frame[17][3] (\data_in_frame[17] [3]), 
         .n57195(n57195), .\data_in_frame[17][4] (\data_in_frame[17] [4]), 
         .n57191(n57191), .\data_in_frame[17][5] (\data_in_frame[17] [5]), 
         .n30169(n30169), .\data_in_frame[17][6] (\data_in_frame[17] [6]), 
         .n57187(n57187), .n57117(n57117), .\data_in_frame[21][0] (\data_in_frame[21] [0]), 
         .n57169(n57169), .n57167(n57167), .n57163(n57163), .n57159(n57159), 
         .\data_in_frame[21][4] (\data_in_frame[21] [4]), .n57155(n57155), 
         .\data_in_frame[21][7] (\data_in_frame[21] [7]), .n29502(n29502), 
         .n29505(n29505), .n29508(n29508), .n29511(n29511), .n29514(n29514), 
         .n29520(n29520), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n57897(n57897), .n29538(n29538), .n29541(n29541), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n57896(n57896), .n29560(n29560), .n57895(n57895), .n29566(n29566), 
         .\data_out_frame[1][3] (\data_out_frame[1] [3]), .n57894(n57894), 
         .n57893(n57893), .n29575(n29575), .n29578(n29578), .n29581(n29581), 
         .\data_in_frame[3][2] (\data_in_frame[3] [2]), .n29584(n29584), 
         .n57892(n57892), .n57891(n57891), .n29592(n29592), .n57890(n57890), 
         .n57889(n57889), .n57888(n57888), .n57887(n57887), .n57886(n57886), 
         .n57885(n57885), .n57884(n57884), .n29600(n29600), .n29423(n29423), 
         .n40525(n40525), .n28352(n28352), .n57883(n57883), .n57882(n57882), 
         .n57881(n57881), .n57880(n57880), .n57879(n57879), .LED_c(LED_c), 
         .n29603(n29603), .n30680(n30680), .n29037(n29037), .n57780(n57780), 
         .n57781(n57781), .n57782(n57782), .n28355(n28355), .n57783(n57783), 
         .n57878(n57878), .n30686(n30686), .n29035(n29035), .n30687(n30687), 
         .n29034(n29034), .n57877(n57877), .n30689(n30689), .n29032(n29032), 
         .n57876(n57876), .n30691(n30691), .n29030(n29030), .n57875(n57875), 
         .n57874(n57874), .n57873(n57873), .n57872(n57872), .n57871(n57871), 
         .n57870(n57870), .n57869(n57869), .n57868(n57868), .n57867(n57867), 
         .n57866(n57866), .n57865(n57865), .n57864(n57864), .n29403(n29403), 
         .n57784(n57784), .n29401(n29401), .\current_limit[1] (current_limit[1]), 
         .n57785(n57785), .n57786(n57786), .n57787(n57787), .n57788(n57788), 
         .n57789(n57789), .n57790(n57790), .n57791(n57791), .n57792(n57792), 
         .n57793(n57793), .n57794(n57794), .n57795(n57795), .n57796(n57796), 
         .n30717(n30717), .n29017(n29017), .n30718(n30718), .n29016(n29016), 
         .n30719(n30719), .n29015(n29015), .n57862(n57862), .n57797(n57797), 
         .n57733(n57733), .n57798(n57798), .n57799(n57799), .n57800(n57800), 
         .n57801(n57801), .n57802(n57802), .DE_c(DE_c), .n26(n26_adj_5701), 
         .n18(n18_adj_5862), .n28363(n28363), .n30778(n30778), .n29013(n29013), 
         .n30779(n30779), .n29012(n29012), .n57861(n57861), .\current[15] (current[15]), 
         .n260(n260), .n58520(n58520), .n28358(n28358), .n28338(n28338), 
         .n15_adj_10(n15_adj_5808), .n25961(n25961), .Kp_23__N_1301(Kp_23__N_1301), 
         .n58561(n58561), .n8_adj_11(n8_adj_5807), .n58766(n58766), .n17(n17_adj_5868), 
         .n18_adj_12(n18_adj_5854), .\motor_state_23__N_91[1] (motor_state_23__N_91[1]), 
         .\motor_state[1] (motor_state[1]), .\motor_state_23__N_91[2] (motor_state_23__N_91[2]), 
         .\motor_state[2] (motor_state[2]), .\motor_state_23__N_91[3] (motor_state_23__N_91[3]), 
         .\motor_state[3] (motor_state[3]), .\motor_state_23__N_91[4] (motor_state_23__N_91[4]), 
         .\motor_state[4] (motor_state[4]), .\motor_state_23__N_91[5] (motor_state_23__N_91[5]), 
         .\motor_state[5] (motor_state[5]), .\motor_state_23__N_91[6] (motor_state_23__N_91[6]), 
         .\motor_state[6] (motor_state[6]), .\motor_state_23__N_91[7] (motor_state_23__N_91[7]), 
         .\motor_state[7] (motor_state[7]), .n28361(n28361), .n10(n10_adj_5940), 
         .\motor_state_23__N_91[9] (motor_state_23__N_91[9]), .\motor_state[9] (motor_state[9]), 
         .\motor_state_23__N_91[10] (motor_state_23__N_91[10]), .\motor_state[10] (motor_state[10]), 
         .\motor_state_23__N_91[11] (motor_state_23__N_91[11]), .\motor_state[11] (motor_state[11]), 
         .\motor_state_23__N_91[12] (motor_state_23__N_91[12]), .\motor_state[12] (motor_state[12]), 
         .\motor_state_23__N_91[13] (motor_state_23__N_91[13]), .\motor_state[13] (motor_state[13]), 
         .\motor_state_23__N_91[14] (motor_state_23__N_91[14]), .\motor_state[14] (motor_state[14]), 
         .n7_adj_13(n7_adj_5831), .\motor_state_23__N_91[21] (motor_state_23__N_91[21]), 
         .\motor_state[21] (motor_state[21]), .n28304(n28304), .\motor_state_23__N_91[17] (motor_state_23__N_91[17]), 
         .\motor_state[17] (motor_state[17]), .n53323(n53323), .\motor_state_23__N_91[19] (motor_state_23__N_91[19]), 
         .\motor_state[19] (motor_state[19]), .\motor_state_23__N_91[20] (motor_state_23__N_91[20]), 
         .\motor_state[20] (motor_state[20]), .n25771(n25771), .\current[7] (current[7]), 
         .\motor_state_23__N_91[22] (motor_state_23__N_91[22]), .\motor_state[22] (motor_state[22]), 
         .\motor_state_23__N_91[23] (motor_state_23__N_91[23]), .\motor_state[23] (motor_state[23]), 
         .n7_adj_14(n7_adj_5858), .\motor_state_23__N_91[15] (motor_state_23__N_91[15]), 
         .\motor_state[15] (motor_state[15]), .\motor_state_23__N_91[18] (motor_state_23__N_91[18]), 
         .\motor_state[18] (motor_state[18]), .n58169(n58169), .n58405(n58405), 
         .n58556(n58556), .\current[6] (current[6]), .\current[5] (current[5]), 
         .\current[4] (current[4]), .\current[3] (current[3]), .\current[2] (current[2]), 
         .\current[1] (current[1]), .\current[0] (current[0]), .\current[11] (current[11]), 
         .\current[10] (current[10]), .\current[9] (current[9]), .\current[8] (current[8]), 
         .n22760(n22760), .n52894(n52894), .n14(n14_adj_5835), .n58366(n58366), 
         .n66452(n66452), .n58711(n58711), .n25819(n25819), .n26235(n26235), 
         .n26405(n26405), .n70252(n70252), .n58046(n58046), .n63899(n63899), 
         .n63900(n63900), .n60683(n60683), .n69300(n69300), .n60931(n60931), 
         .n63903(n63903), .n63902(n63902), .tx_o(tx_o), .r_Clock_Count({r_Clock_Count_adj_6024}), 
         .tx_enable(tx_enable), .baudrate({baudrate}), .n27845(n27845), 
         .n58988(n58988), .\r_SM_Main[2] (r_SM_Main[2]), .r_Rx_Data(r_Rx_Data), 
         .RX_N_2(RX_N_2), .r_Clock_Count_adj_23({r_Clock_Count}), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), 
         .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), 
         .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), 
         .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .n61478(n61478), .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), 
         .\r_SM_Main[1] (r_SM_Main[1]), .n4939(n4939), .n25566(n25566), 
         .n29596(n29596), .n29595(n29595), .n29591(n29591), .n29590(n29590), 
         .n29559(n29559), .n29558(n29558), .n29557(n29557), .\r_Bit_Index[0] (r_Bit_Index[0]), 
         .n61043(n61043), .n30440(n30440), .n53943(n53943), .n30436(n30436), 
         .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), .n61750(n61750), .n61702(n61702), 
         .n61734(n61734), .n61814(n61814), .n61782(n61782), .n61766(n61766), 
         .n61798(n61798), .n61718(n61718), .n57927(n57927), .n27722(n27722)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i51158_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n66388));
    defparam i51158_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_4_lut_adj_2188 (.I0(n3222), .I1(n17_adj_5921), .I2(n3289), 
            .I3(n3237), .O(n62332));
    defparam i1_4_lut_adj_2188.LUT_INIT = 16'heefc;
    SB_LUT4 i11_2_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26235));   // verilog/coms.v(100[12:26])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_2189 (.I0(n3225), .I1(n23_adj_5923), .I2(n3292), 
            .I3(n3237), .O(n62334));
    defparam i1_4_lut_adj_2189.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2190 (.I0(n66388), .I1(n5_adj_5869), .I2(n66389), 
            .I3(n3237), .O(n54403));
    defparam i1_4_lut_adj_2190.LUT_INIT = 16'h88c0;
    SB_LUT4 i1_4_lut_adj_2191 (.I0(n3218), .I1(n62330), .I2(n3285), .I3(n3237), 
            .O(n62338));
    defparam i1_4_lut_adj_2191.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2192 (.I0(n62338), .I1(n54403), .I2(n62334), 
            .I3(n62332), .O(n62342));
    defparam i1_4_lut_adj_2192.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2193 (.I0(n3214), .I1(n62342), .I2(n3281), .I3(n3237), 
            .O(n62344));
    defparam i1_4_lut_adj_2193.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2194 (.I0(n3207), .I1(n62344), .I2(n3274), .I3(n3237), 
            .O(n62346));
    defparam i1_4_lut_adj_2194.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2195 (.I0(n3210), .I1(n62224), .I2(n3277), .I3(n3237), 
            .O(n62226));
    defparam i1_4_lut_adj_2195.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_2196 (.I0(n62386), .I1(n3208), .I2(n3275), .I3(n3237), 
            .O(n61041));
    defparam i1_4_lut_adj_2196.LUT_INIT = 16'heefa;
    SB_LUT4 i1_4_lut_adj_2197 (.I0(n62346), .I1(n3206), .I2(n3273), .I3(n3237), 
            .O(n61029));
    defparam i1_4_lut_adj_2197.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_30__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2198 (.I0(n61), .I1(n61029), .I2(n61041), .I3(n62226), 
            .O(n62232));
    defparam i1_4_lut_adj_2198.LUT_INIT = 16'hfffe;
    SB_LUT4 i53744_4_lut (.I0(n62232), .I1(n3204), .I2(n3271), .I3(n3237), 
            .O(n43071));
    defparam i53744_4_lut.LUT_INIT = 16'h1105;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2199 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n57738));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2199.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2200 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n57739));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2200.LUT_INIT = 16'h2300;
    TLI4970 tli (.GND_net(GND_net), .n29837(n29837), .\data[15] (data_adj_6010[15]), 
            .n29836(n29836), .\data[12] (data_adj_6010[12]), .n29835(n29835), 
            .\data[11] (data_adj_6010[11]), .n29834(n29834), .\data[10] (data_adj_6010[10]), 
            .n29833(n29833), .\data[9] (data_adj_6010[9]), .n29832(n29832), 
            .\data[8] (data_adj_6010[8]), .n29831(n29831), .\data[7] (data_adj_6010[7]), 
            .n29830(n29830), .\data[6] (data_adj_6010[6]), .n29829(n29829), 
            .\data[5] (data_adj_6010[5]), .n29828(n29828), .\data[4] (data_adj_6010[4]), 
            .n29827(n29827), .\data[3] (data_adj_6010[3]), .n29826(n29826), 
            .\data[2] (data_adj_6010[2]), .n29825(n29825), .\data[1] (data_adj_6010[1]), 
            .clk16MHz(clk16MHz), .VCC_net(VCC_net), .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), 
            .n29625(n29625), .\current[0] (current[0]), .n30445(n30445), 
            .\data[0] (data_adj_6010[0]), .n30365(n30365), .\current[1] (current[1]), 
            .n30364(n30364), .\current[2] (current[2]), .n30363(n30363), 
            .\current[3] (current[3]), .n30362(n30362), .\current[4] (current[4]), 
            .n30361(n30361), .\current[5] (current[5]), .n30360(n30360), 
            .\current[6] (current[6]), .n30359(n30359), .\current[7] (current[7]), 
            .n30358(n30358), .\current[8] (current[8]), .n30357(n30357), 
            .\current[9] (current[9]), .n30356(n30356), .\current[10] (current[10]), 
            .n30355(n30355), .\current[11] (current[11]), .n6(n6_adj_5809), 
            .n6_adj_4(n6_adj_5777), .n5(n5_adj_5812), .n5_adj_5(n5_adj_5789), 
            .n6_adj_6(n6_adj_5774), .state_7__N_4320(state_7__N_4320), .n42331(n42331), 
            .n27704(n27704), .\current[15] (current[15]), .n25555(n25555), 
            .n25573(n25573), .n25579(n25579), .n25563(n25563), .n25544(n25544), 
            .n11(n11_adj_5791)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(405[11] 411[4])
    SB_LUT4 i15622_4_lut (.I0(state_7__N_4127[3]), .I1(data_adj_6002[7]), 
            .I2(n42355), .I3(n25568), .O(n29653));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15622_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15623_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n22760), .I3(GND_net), .O(n29654));   // verilog/coms.v(130[12] 305[6])
    defparam i15623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15624_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n22760), .I3(GND_net), .O(n29655));   // verilog/coms.v(130[12] 305[6])
    defparam i15624_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(0)_U0  quad_counter0 (.\a_new[1] (a_new[1]), .\b_new[1] (b_new[1]), 
            .debounce_cnt_N_3834(debounce_cnt_N_3834), .a_prev(a_prev), 
            .b_prev(b_prev), .position_31__N_3837(position_31__N_3837), 
            .GND_net(GND_net), .ENCODER0_B_N_keep(ENCODER0_B_N), .n1779(clk16MHz), 
            .ENCODER0_A_N_keep(ENCODER0_A_N), .n29707(n29707), .n1742(n1742), 
            .n29706(n29706), .n29672(n29672), .n1744(n1744), .\encoder0_position[30] (encoder0_position[30]), 
            .\encoder0_position[29] (encoder0_position[29]), .\encoder0_position[28] (encoder0_position[28]), 
            .\encoder0_position[27] (encoder0_position[27]), .\encoder0_position[26] (encoder0_position[26]), 
            .\encoder0_position[25] (encoder0_position[25]), .\encoder0_position[24] (encoder0_position[24]), 
            .\encoder0_position[23] (encoder0_position[23]), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(305[27] 311[6])
    SB_LUT4 i15625_3_lut (.I0(a_prev_adj_5782), .I1(a_new_adj_5988[1]), 
            .I2(debounce_cnt_N_3834_adj_5784), .I3(GND_net), .O(n29656));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4306_i1_3_lut (.I0(encoder0_position[0]), .I1(n32), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_4306_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53735_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69461));
    defparam i53735_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_2201 (.I0(n3220), .I1(n3218), .I2(n3225), .I3(GND_net), 
            .O(n62660));
    defparam i1_3_lut_adj_2201.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2202 (.I0(n3215), .I1(n3217), .I2(n3224), .I3(n3228), 
            .O(n62752));
    defparam i1_4_lut_adj_2202.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2203 (.I0(n3226), .I1(n3223), .I2(n3222), .I3(n3227), 
            .O(n62676));
    defparam i1_4_lut_adj_2203.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2204 (.I0(n3209), .I1(n3213), .I2(n62676), .I3(GND_net), 
            .O(n62680));
    defparam i1_3_lut_adj_2204.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2205 (.I0(n3210), .I1(n3211), .I2(n3214), .I3(n62752), 
            .O(n62758));
    defparam i1_4_lut_adj_2205.LUT_INIT = 16'hfffe;
    SB_LUT4 i29124_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n43051));
    defparam i29124_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2206 (.I0(n62660), .I1(n3216), .I2(n3221), .I3(n3219), 
            .O(n62664));
    defparam i1_4_lut_adj_2206.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2207 (.I0(n3229), .I1(n43051), .I2(n3230), .I3(n3231), 
            .O(n59785));
    defparam i1_4_lut_adj_2207.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut_adj_2208 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[16] [0]), .I3(\data_out_frame[18] [2]), 
            .O(n60683));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_2208.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2209 (.I0(n3207), .I1(n62758), .I2(n62680), .I3(n3208), 
            .O(n62684));
    defparam i1_4_lut_adj_2209.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2210 (.I0(n3205), .I1(n3212), .I2(n59785), .I3(n62664), 
            .O(n62670));
    defparam i1_4_lut_adj_2210.LUT_INIT = 16'hfffe;
    SB_LUT4 i53740_4_lut (.I0(n3206), .I1(n62670), .I2(n62684), .I3(n3204), 
            .O(n3237));
    defparam i53740_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5910));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_2211 (.I0(\data_out_frame[18] [1]), .I1(n26111), 
            .I2(n58651), .I3(n2076), .O(n20_adj_5864));
    defparam i8_4_lut_adj_2211.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_2212 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[19] [4]), 
            .I2(n58570), .I3(n52894), .O(n19_adj_5865));
    defparam i7_4_lut_adj_2212.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n60931), .I1(n25819), .I2(n26405), .I3(n69300), 
            .O(n21_adj_5863));
    defparam i9_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i11_3_lut (.I0(n21_adj_5863), .I1(n19_adj_5865), .I2(n20_adj_5864), 
            .I3(GND_net), .O(n58366));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2213 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n57740));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2213.LUT_INIT = 16'h2300;
    pwm PWM (.GND_net(GND_net), .n2874(n2874), .pwm_out(pwm_out), .clk32MHz(clk32MHz), 
        .reset(reset), .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2214 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n28940));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2214.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2215 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n57741));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2215.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5909));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16688_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n30719));   // verilog/coms.v(130[12] 305[6])
    defparam i16688_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16687_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n30718));   // verilog/coms.v(130[12] 305[6])
    defparam i16687_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16686_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n30717));   // verilog/coms.v(130[12] 305[6])
    defparam i16686_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16660_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n30691));   // verilog/coms.v(130[12] 305[6])
    defparam i16660_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    motorControl control (.GND_net(GND_net), .n182(n182), .IntegralLimit({IntegralLimit}), 
            .n156(n156), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), 
            .\Ki[7] (Ki[7]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .\Ki[8] (Ki[8]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Ki[9] (Ki[9]), 
            .\Ki[1] (Ki[1]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .n150(n150), .\Ki[0] (Ki[0]), 
            .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .n6(n6_adj_5916), .n37154(n37154), 
            .n20194(n20194), .\Kp[13] (Kp[13]), .n20185(n20185), .n214(n214), 
            .\Ki[6] (Ki[6]), .\Kp[14] (Kp[14]), .clk16MHz(clk16MHz), .duty({duty}), 
            .reset(reset), .n37050(n37050), .n4(n4_adj_5918), .\Kp[11] (Kp[11]), 
            .\Kp[12] (Kp[12]), .PWMLimit({PWMLimit}), .n406(n406), .setpoint({setpoint}), 
            .n15(n15_adj_5808), .n405(n405), .\Kp[15] (Kp[15]), .n478(n478), 
            .n135(n135), .n500(n500), .\Ki[10] (Ki[10]), .VCC_net(VCC_net), 
            .n187(n187), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .n41(n41_adj_5867), 
            .deadband({deadband}), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .n219(n219), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .n20112(n20112), .n20113(n20113), .n7(n7_adj_5858), .n56(n56), 
            .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .\motor_state[13] (motor_state[13]), .\motor_state[12] (motor_state[12]), 
            .\motor_state[11] (motor_state[11]), .\motor_state[10] (motor_state[10]), 
            .\motor_state[9] (motor_state[9]), .n10(n10_adj_5940), .\motor_state[7] (motor_state[7]), 
            .\motor_state[6] (motor_state[6]), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .\motor_state[1] (motor_state[1]), 
            .n18(n18_adj_5854), .\duty_23__N_3602[7] (duty_23__N_3602[7]), 
            .\duty_23__N_3602[4] (duty_23__N_3602[4]), .n624(n624), .n551(n551), 
            .n478_adj_1(n478_adj_5846), .n405_adj_2(n405_adj_5857), .n332(n332), 
            .n259(n259), .n186(n186), .n113(n113), .n244(n244), .n36515(n36515), 
            .n41_adj_3(n41), .\data_in_frame[9][7] (\data_in_frame[9] [7]), 
            .\data_in_frame[6][3] (\data_in_frame[6] [3]), .\data_in_frame[8][4] (\data_in_frame[8] [4]), 
            .\data_in_frame[8][2] (\data_in_frame[8] [2]), .n58520(n58520), 
            .\data_in_frame[4][2] (\data_in_frame[4] [2]), .\data_in_frame[8][6] (\data_in_frame[8] [6]), 
            .\data_in_frame[1][6] (\data_in_frame[1] [6]), .\data_in_frame[12][0] (\data_in_frame[12] [0]), 
            .n58075(n58075), .n58405(n58405), .n58556(n58556), .\data_in_frame[3][7] (\data_in_frame[3] [7]), 
            .\data_in_frame[4][1] (\data_in_frame[4] [1]), .\data_in_frame[8][3] (\data_in_frame[8] [3]), 
            .n58766(n58766), .n50204(n50204), .n50001(n50001), .n62(n62_adj_5866), 
            .n20158(n20158), .n20159(n20159), .n42880(n42880)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 303[4])
    SB_LUT4 i16658_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n30689));   // verilog/coms.v(130[12] 305[6])
    defparam i16658_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16656_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n30687));   // verilog/coms.v(130[12] 305[6])
    defparam i16656_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16655_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n30686));   // verilog/coms.v(130[12] 305[6])
    defparam i16655_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, VCC_net, timer, 
            GND_net, \neo_pixel_transmitter.t0 , n29644, n27799, \bit_ctr[4] , 
            n30294, n30293, n30292, n30291, n30289, n30288, n30287, 
            n30286, n30285, n30276, n30187, \bit_ctr[1] , n56711, 
            state, neopxl_color, \bit_ctr[0] , NEOPXL_c, n110, LED_c, 
            n42981, n52805, n66110, \color_bit_N_502[1] , n31) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    input VCC_net;
    output [10:0]timer;
    input GND_net;
    output [10:0]\neo_pixel_transmitter.t0 ;
    input n29644;
    output n27799;
    output \bit_ctr[4] ;
    input n30294;
    input n30293;
    input n30292;
    input n30291;
    input n30289;
    input n30288;
    input n30287;
    input n30286;
    input n30285;
    input n30276;
    input n30187;
    output \bit_ctr[1] ;
    input n56711;
    output [1:0]state;
    input [23:0]neopxl_color;
    output \bit_ctr[0] ;
    output NEOPXL_c;
    output n110;
    input LED_c;
    output n42981;
    output n52805;
    output n66110;
    output \color_bit_N_502[1] ;
    output n31;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n57942, \neo_pixel_transmitter.done , 
        start_N_507, n7, start;
    wire [10:0]n13;
    
    wire n50330;
    wire [10:0]n49;
    
    wire n51547, n51548, n51546, n51545, n51544, n50331;
    wire [31:0]n137;
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    
    wire n29094;
    wire [10:0]one_wire_N_479;
    
    wire n50339, n50338, n103, n52285, n4, n57_adj_5690, n117, 
        n47, n66450, n40200, n63857, n63858, n1, n27789, n28808;
    wire [1:0]state_1__N_440;
    
    wire n27803, n29098, n63894, n63893, \neo_pixel_transmitter.done_N_524 , 
        n68502, n61219, n50337, n50336, n50335, n50334, n50333, 
        n50332, n4_adj_5693, n70183, n51553, n51552, n51551, n51550, 
        n51549, n70189, n70489, n57_adj_5694;
    wire [5:0]color_bit_N_502;
    
    wire n66108, n6893, n8_adj_5695, n59002, n4_adj_5696, n31_c, 
        n94, n66448, n10_adj_5697, n69306, n58905, n37, n58885, 
        n68501, n52829, n42983, n63816, n63815, n70276, n63817, 
        n63840, n70192, n70492, n63839, n70186, n63841, n60564, 
        n60563, n70273, n16, n63537, n61178;
    
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n57942), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 116[6])
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n50330));
    SB_LUT4 timer_1939_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n51547), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_6 (.CI(n51547), .I0(GND_net), .I1(timer[4]), 
            .CO(n51548));
    SB_LUT4 timer_1939_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n51546), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_5 (.CI(n51546), .I0(GND_net), .I1(timer[3]), 
            .CO(n51547));
    SB_LUT4 timer_1939_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n51545), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_4 (.CI(n51545), .I0(GND_net), .I1(timer[2]), 
            .CO(n51546));
    SB_LUT4 timer_1939_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n51544), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_3 (.CI(n50330), .I0(timer[1]), .I1(n13[1]), 
            .CO(n50331));
    SB_CARRY timer_1939_add_4_3 (.CI(n51544), .I0(GND_net), .I1(timer[1]), 
            .CO(n51545));
    SB_LUT4 timer_1939_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n51544));
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29644));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF timer_1939__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr[2]), .C(clk16MHz), .E(n27799), .D(n137[2]), 
            .R(n29094));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr[3]), .C(clk16MHz), .E(n27799), .D(n137[3]), 
            .R(n29094));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i4 (.Q(\bit_ctr[4] ), .C(clk16MHz), .E(n27799), 
            .D(n137[4]), .R(n29094));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF timer_1939__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1939__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n30294));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n30293));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n30292));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n30291));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n30289));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n30288));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n30287));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n30286));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n30285));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n30276));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF bit_ctr_i1 (.Q(\bit_ctr[1] ), .C(clk16MHz), .D(n30187));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n56711));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n50339), .O(one_wire_N_479[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n13[9]), 
            .I3(n50338), .O(one_wire_N_479[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i43195_4_lut (.I0(n103), .I1(n52285), .I2(n4), .I3(state[0]), 
            .O(n57_adj_5690));   // verilog/neopixel.v(16[11:16])
    defparam i43195_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_2_lut (.I0(n117), .I1(one_wire_N_479[10]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/neopixel.v(6[16:24])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut (.I0(n66450), .I1(n40200), .I2(state[1]), .I3(state[0]), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i53615_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 115[11])
    defparam i53615_2_lut.LUT_INIT = 16'hdddd;
    SB_CARRY sub_67_add_2_11 (.CI(n50338), .I0(timer[9]), .I1(n13[9]), 
            .CO(n50339));
    SB_LUT4 i48131_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n63857));
    defparam i48131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48132_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n63858));
    defparam i48132_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_i0 (.Q(\bit_ctr[0] ), .C(clk16MHz), .E(n27789), 
            .D(n1), .R(n28808));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n27803), .D(state_1__N_440[0]), 
            .S(n29098));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i48168_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n63894));
    defparam i48168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48167_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n63893));
    defparam i48167_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n68502), .D(\neo_pixel_transmitter.done_N_524 ), 
            .R(n61219));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n50337), .O(one_wire_N_479[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n50337), .I0(timer[8]), .I1(n13[8]), 
            .CO(n50338));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n50336), .O(one_wire_N_479[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n50336), .I0(timer[7]), .I1(n13[7]), 
            .CO(n50337));
    SB_LUT4 sub_67_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n13[6]), 
            .I3(n50335), .O(one_wire_N_479[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_8 (.CI(n50335), .I0(timer[6]), .I1(n13[6]), 
            .CO(n50336));
    SB_LUT4 sub_67_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n13[5]), 
            .I3(n50334), .O(one_wire_N_479[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_7 (.CI(n50334), .I0(timer[5]), .I1(n13[5]), 
            .CO(n50335));
    SB_LUT4 sub_67_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n13[4]), 
            .I3(n50333), .O(one_wire_N_479[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_6 (.CI(n50333), .I0(timer[4]), .I1(n13[4]), 
            .CO(n50334));
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n50332), .O(one_wire_N_479[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_5 (.CI(n50332), .I0(timer[3]), .I1(n13[3]), 
            .CO(n50333));
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n50331), .O(one_wire_N_479[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_4 (.CI(n50331), .I0(timer[2]), .I1(n13[2]), 
            .CO(n50332));
    SB_LUT4 sub_67_add_2_3_lut (.I0(one_wire_N_479[2]), .I1(timer[1]), .I2(n13[1]), 
            .I3(n50330), .O(n4_adj_5693)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 bit_ctr_0__bdd_4_lut_54452_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(\bit_ctr[1] ), .O(n70183));
    defparam bit_ctr_0__bdd_4_lut_54452_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 timer_1939_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n51553), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1939_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n51552), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_11 (.CI(n51552), .I0(GND_net), .I1(timer[9]), 
            .CO(n51553));
    SB_LUT4 timer_1939_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n51551), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_10 (.CI(n51551), .I0(GND_net), .I1(timer[8]), 
            .CO(n51552));
    SB_LUT4 timer_1939_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n51550), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_9 (.CI(n51550), .I0(GND_net), .I1(timer[7]), 
            .CO(n51551));
    SB_LUT4 timer_1939_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n51549), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_8 (.CI(n51549), .I0(GND_net), .I1(timer[6]), 
            .CO(n51550));
    SB_LUT4 timer_1939_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n51548), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1939_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1939_add_4_7 (.CI(n51548), .I0(GND_net), .I1(timer[5]), 
            .CO(n51549));
    SB_LUT4 bit_ctr_0__bdd_4_lut_54697_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(\bit_ctr[1] ), .O(n70189));
    defparam bit_ctr_0__bdd_4_lut_54697_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n47), .I3(\neo_pixel_transmitter.done_N_524 ), 
            .O(n61219));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_4_lut_4_lut (.I0(n110), .I1(state[1]), .I2(n40200), .I3(state[0]), 
            .O(n27803));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'heee2;
    SB_LUT4 i1_2_lut_3_lut (.I0(n110), .I1(state[1]), .I2(n27789), .I3(GND_net), 
            .O(n27799));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(\bit_ctr[1] ), .O(n70489));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n57_adj_5694), .I2(LED_c), 
            .I3(state[1]), .O(n27789));   // verilog/neopixel.v(35[4] 115[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_LUT4 i14777_2_lut_4_lut (.I0(state[0]), .I1(n57_adj_5694), .I2(LED_c), 
            .I3(state[1]), .O(n28808));   // verilog/neopixel.v(35[4] 115[11])
    defparam i14777_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 sub_67_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29055_2_lut_3_lut_4_lut (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), 
            .I2(bit_ctr[3]), .I3(bit_ctr[2]), .O(n42981));
    defparam i29055_2_lut_3_lut_4_lut.LUT_INIT = 16'hf0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), 
            .I2(bit_ctr[3]), .I3(bit_ctr[2]), .O(n52805));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0f1e;
    SB_LUT4 i1_2_lut_3_lut_adj_1775 (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), 
            .I2(bit_ctr[2]), .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1775.LUT_INIT = 16'h1e1e;
    SB_LUT4 i50382_2_lut_3_lut (.I0(\bit_ctr[4] ), .I1(n42981), .I2(n52805), 
            .I3(GND_net), .O(n66108));   // verilog/neopixel.v(21[26:38])
    defparam i50382_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i2107_3_lut_4_lut (.I0(bit_ctr[2]), .I1(n6893), .I2(bit_ctr[3]), 
            .I3(\bit_ctr[4] ), .O(n137[4]));   // verilog/neopixel.v(68[23:32])
    defparam i2107_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i2093_2_lut_3_lut (.I0(bit_ctr[2]), .I1(\bit_ctr[1] ), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n137[2]));   // verilog/neopixel.v(68[23:32])
    defparam i2093_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_3_lut_4_lut (.I0(color_bit_N_502[2]), .I1(\bit_ctr[4] ), 
            .I2(n42981), .I3(\bit_ctr[0] ), .O(n8_adj_5695));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hffeb;
    SB_LUT4 i44_3_lut_4_lut (.I0(one_wire_N_479[3]), .I1(n4_adj_5693), .I2(one_wire_N_479[2]), 
            .I3(\neo_pixel_transmitter.done ), .O(n59002));
    defparam i44_3_lut_4_lut.LUT_INIT = 16'hfa88;
    SB_LUT4 i1_2_lut_3_lut_adj_1776 (.I0(n103), .I1(start), .I2(state[1]), 
            .I3(GND_net), .O(n4_adj_5696));
    defparam i1_2_lut_3_lut_adj_1776.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_3_lut (.I0(n103), .I1(one_wire_N_479[2]), .I2(one_wire_N_479[3]), 
            .I3(GND_net), .O(n31_c));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1777 (.I0(one_wire_N_479[3]), .I1(n4_adj_5693), 
            .I2(n103), .I3(GND_net), .O(n94));
    defparam i1_2_lut_3_lut_adj_1777.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2100_2_lut_3_lut_4_lut (.I0(bit_ctr[2]), .I1(\bit_ctr[1] ), 
            .I2(\bit_ctr[0] ), .I3(bit_ctr[3]), .O(n137[3]));   // verilog/neopixel.v(68[23:32])
    defparam i2100_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i50901_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n117), 
            .I3(one_wire_N_479[10]), .O(n66448));   // verilog/neopixel.v(34[12] 116[6])
    defparam i50901_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_adj_1778 (.I0(one_wire_N_479[9]), .I1(one_wire_N_479[8]), 
            .I2(GND_net), .I3(GND_net), .O(n117));
    defparam i1_2_lut_adj_1778.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_479[3]), .I1(n4_adj_5693), .I2(GND_net), 
            .I3(GND_net), .O(n52285));   // verilog/neopixel.v(101[14:24])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1779 (.I0(one_wire_N_479[2]), .I1(one_wire_N_479[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1779.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_479[5]), .I1(one_wire_N_479[4]), .I2(n117), 
            .I3(one_wire_N_479[7]), .O(n10_adj_5697));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(one_wire_N_479[6]), .I1(n10_adj_5697), .I2(one_wire_N_479[10]), 
            .I3(GND_net), .O(n103));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i53580_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n69306));
    defparam i53580_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i43232_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n58905));
    defparam i43232_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut (.I0(n94), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n37));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i54366_4_lut (.I0(n37), .I1(n58905), .I2(n31_c), .I3(n69306), 
            .O(n57942));
    defparam i54366_4_lut.LUT_INIT = 16'hdddc;
    SB_LUT4 i26251_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(16[11:16])
    defparam i26251_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 sub_67_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1780 (.I0(\neo_pixel_transmitter.done ), .I1(n117), 
            .I2(one_wire_N_479[10]), .I3(GND_net), .O(n40200));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_3_lut_adj_1780.LUT_INIT = 16'h4040;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45_4_lut (.I0(n31_c), .I1(n47), .I2(state[1]), .I3(start), 
            .O(n58885));
    defparam i45_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52775_4_lut (.I0(n58885), .I1(n94), .I2(\neo_pixel_transmitter.done ), 
            .I3(n58905), .O(n68501));
    defparam i52775_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i52776_4_lut (.I0(n68501), .I1(n59002), .I2(state[0]), .I3(n4_adj_5696), 
            .O(n68502));
    defparam i52776_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 i2_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_524 ));
    defparam i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50384_2_lut_3_lut (.I0(\bit_ctr[4] ), .I1(n42981), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n66110));
    defparam i50384_2_lut_3_lut.LUT_INIT = 16'h0606;
    SB_LUT4 i1_2_lut_adj_1781 (.I0(\bit_ctr[4] ), .I1(n42981), .I2(GND_net), 
            .I3(GND_net), .O(n52829));
    defparam i1_2_lut_adj_1781.LUT_INIT = 16'h6666;
    SB_LUT4 i29057_2_lut (.I0(\bit_ctr[4] ), .I1(n42981), .I2(GND_net), 
            .I3(GND_net), .O(n42983));
    defparam i29057_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1782 (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_502[1] ));
    defparam i1_2_lut_adj_1782.LUT_INIT = 16'h6666;
    SB_LUT4 i1082_4_lut (.I0(\color_bit_N_502[1] ), .I1(n42983), .I2(n8_adj_5695), 
            .I3(n52805), .O(n57_adj_5694));   // verilog/neopixel.v(21[26:38])
    defparam i1082_4_lut.LUT_INIT = 16'h3233;
    SB_LUT4 i2088_2_lut (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n6893));   // verilog/neopixel.v(68[23:32])
    defparam i2088_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15063_2_lut (.I0(n27799), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29094));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15063_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14_4_lut (.I0(n66448), .I1(n57_adj_5690), .I2(\neo_pixel_transmitter.done ), 
            .I3(n58905), .O(n29098));   // verilog/neopixel.v(34[12] 116[6])
    defparam i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i48090_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n63816));
    defparam i48090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48089_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n63815));
    defparam i48089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48091_4_lut (.I0(n63816), .I1(n70276), .I2(n52829), .I3(n52805), 
            .O(n63817));
    defparam i48091_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48114_4_lut (.I0(n63817), .I1(n63815), .I2(n52829), .I3(\color_bit_N_502[1] ), 
            .O(n63840));
    defparam i48114_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i48113_3_lut (.I0(n70192), .I1(n70492), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n63839));
    defparam i48113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48115_3_lut (.I0(n63840), .I1(n70186), .I2(n66110), .I3(GND_net), 
            .O(n63841));
    defparam i48115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28250_4_lut (.I0(n63841), .I1(n57_adj_5694), .I2(n63839), 
            .I3(n66108), .O(state_1__N_440[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i28250_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut (.I0(start), .I1(n31_c), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n60564));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_3_lut_adj_1783 (.I0(n94), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(GND_net), .O(n60563));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_3_lut_adj_1783.LUT_INIT = 16'hf7f7;
    SB_LUT4 state_1__I_0_102_Mux_0_i1_4_lut (.I0(n60563), .I1(n60564), .I2(state[0]), 
            .I3(\bit_ctr[0] ), .O(n1));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_102_Mux_0_i1_4_lut.LUT_INIT = 16'hca35;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(\color_bit_N_502[1] ), .I1(n63893), 
            .I2(n63894), .I3(color_bit_N_502[2]), .O(n70273));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70273_bdd_4_lut (.I0(n70273), .I1(n63858), .I2(n63857), .I3(color_bit_N_502[2]), 
            .O(n70276));
    defparam n70273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n70489_bdd_4_lut (.I0(n70489), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(\color_bit_N_502[1] ), .O(n70492));
    defparam n70489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1784 (.I0(\neo_pixel_transmitter.done ), .I1(n57_adj_5690), 
            .I2(start), .I3(GND_net), .O(n110));   // verilog/neopixel.v(16[11:16])
    defparam i1_2_lut_3_lut_adj_1784.LUT_INIT = 16'h0808;
    SB_LUT4 i51587_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n57_adj_5690), 
            .I2(start), .I3(GND_net), .O(n66450));   // verilog/neopixel.v(16[11:16])
    defparam i51587_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i6_4_lut (.I0(n69306), .I1(one_wire_N_479[6]), .I2(one_wire_N_479[10]), 
            .I3(one_wire_N_479[4]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i47820_4_lut (.I0(one_wire_N_479[3]), .I1(one_wire_N_479[5]), 
            .I2(one_wire_N_479[9]), .I3(one_wire_N_479[7]), .O(n63537));
    defparam i47820_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n63537), .I1(one_wire_N_479[2]), .I2(n16), .I3(one_wire_N_479[8]), 
            .O(n61178));
    defparam i9_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(start), .I2(n61178), .I3(n37), 
            .O(n31));
    defparam i1_4_lut.LUT_INIT = 16'hbbba;
    SB_LUT4 n70189_bdd_4_lut (.I0(n70189), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(\color_bit_N_502[1] ), .O(n70192));
    defparam n70189_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n70183_bdd_4_lut (.I0(n70183), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(\color_bit_N_502[1] ), .O(n70186));
    defparam n70183_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (a_prev, b_prev, a_new, b_new, position_31__N_3837, 
            ENCODER1_B_N_keep, n1779, ENCODER1_A_N_keep, n1786, GND_net, 
            n1788, n1790, n1792, n1794, n1796, \encoder1_position[25] , 
            \encoder1_position[24] , \encoder1_position[23] , \encoder1_position[22] , 
            \encoder1_position[21] , \encoder1_position[20] , \encoder1_position[19] , 
            \encoder1_position[18] , \encoder1_position[17] , \encoder1_position[16] , 
            \encoder1_position[15] , \encoder1_position[14] , \encoder1_position[13] , 
            \encoder1_position[12] , \encoder1_position[11] , \encoder1_position[10] , 
            \encoder1_position[9] , \encoder1_position[8] , \encoder1_position[7] , 
            \encoder1_position[6] , \encoder1_position[5] , \encoder1_position[4] , 
            n29664, n1784, \encoder1_position[3] , n29656, \encoder1_position[2] , 
            n1822, n1824, VCC_net, n29397, debounce_cnt_N_3834) /* synthesis lattice_noprune=1 */ ;
    output a_prev;
    output b_prev;
    output [1:0]a_new;
    output [1:0]b_new;
    output position_31__N_3837;
    input ENCODER1_B_N_keep;
    input n1779;
    input ENCODER1_A_N_keep;
    output n1786;
    input GND_net;
    output n1788;
    output n1790;
    output n1792;
    output n1794;
    output n1796;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    input n29664;
    output n1784;
    output \encoder1_position[3] ;
    input n29656;
    output \encoder1_position[2] ;
    output n1822;
    output n1824;
    input VCC_net;
    input n29397;
    output debounce_cnt_N_3834;
    
    wire [1:0]b_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3841, n51676, n51675, n51674, n51673, n51672, 
        n51671, n51670, n51669, n51668, n51667, n51666, n51665, 
        n51664, n51663, n51662, n51661, n51660, n51659, n51658, 
        n51657, n51656, n51655, n51654, n51653, n51652, n51651, 
        n51650, n51649, n51648, n51647, n51646;
    
    SB_LUT4 position_31__I_938_4_lut (.I0(a_prev), .I1(b_prev), .I2(a_new[1]), 
            .I3(b_new[1]), .O(position_31__N_3837));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_938_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF b_new_i0 (.Q(b_new_c[0]), .C(n1779), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1779), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1945_add_4_33_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1786), .I3(n51676), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1945_add_4_32_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1788), .I3(n51675), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_32 (.CI(n51675), .I0(direction_N_3841), 
            .I1(n1788), .CO(n51676));
    SB_LUT4 position_1945_add_4_31_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1790), .I3(n51674), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_31 (.CI(n51674), .I0(direction_N_3841), 
            .I1(n1790), .CO(n51675));
    SB_LUT4 position_1945_add_4_30_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1792), .I3(n51673), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_30 (.CI(n51673), .I0(direction_N_3841), 
            .I1(n1792), .CO(n51674));
    SB_LUT4 position_1945_add_4_29_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1794), .I3(n51672), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_29 (.CI(n51672), .I0(direction_N_3841), 
            .I1(n1794), .CO(n51673));
    SB_LUT4 position_1945_add_4_28_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1796), .I3(n51671), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_28 (.CI(n51671), .I0(direction_N_3841), 
            .I1(n1796), .CO(n51672));
    SB_LUT4 position_1945_add_4_27_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[25] ), .I3(n51670), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_27 (.CI(n51670), .I0(direction_N_3841), 
            .I1(\encoder1_position[25] ), .CO(n51671));
    SB_LUT4 position_1945_add_4_26_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[24] ), .I3(n51669), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_26 (.CI(n51669), .I0(direction_N_3841), 
            .I1(\encoder1_position[24] ), .CO(n51670));
    SB_LUT4 position_1945_add_4_25_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[23] ), .I3(n51668), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_25 (.CI(n51668), .I0(direction_N_3841), 
            .I1(\encoder1_position[23] ), .CO(n51669));
    SB_LUT4 position_1945_add_4_24_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[22] ), .I3(n51667), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_24 (.CI(n51667), .I0(direction_N_3841), 
            .I1(\encoder1_position[22] ), .CO(n51668));
    SB_LUT4 position_1945_add_4_23_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[21] ), .I3(n51666), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_23 (.CI(n51666), .I0(direction_N_3841), 
            .I1(\encoder1_position[21] ), .CO(n51667));
    SB_LUT4 position_1945_add_4_22_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[20] ), .I3(n51665), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_22 (.CI(n51665), .I0(direction_N_3841), 
            .I1(\encoder1_position[20] ), .CO(n51666));
    SB_LUT4 position_1945_add_4_21_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[19] ), .I3(n51664), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_21 (.CI(n51664), .I0(direction_N_3841), 
            .I1(\encoder1_position[19] ), .CO(n51665));
    SB_LUT4 position_1945_add_4_20_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[18] ), .I3(n51663), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_20 (.CI(n51663), .I0(direction_N_3841), 
            .I1(\encoder1_position[18] ), .CO(n51664));
    SB_LUT4 position_1945_add_4_19_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[17] ), .I3(n51662), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_19 (.CI(n51662), .I0(direction_N_3841), 
            .I1(\encoder1_position[17] ), .CO(n51663));
    SB_LUT4 position_1945_add_4_18_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[16] ), .I3(n51661), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_18 (.CI(n51661), .I0(direction_N_3841), 
            .I1(\encoder1_position[16] ), .CO(n51662));
    SB_LUT4 position_1945_add_4_17_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[15] ), .I3(n51660), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_17 (.CI(n51660), .I0(direction_N_3841), 
            .I1(\encoder1_position[15] ), .CO(n51661));
    SB_LUT4 position_1945_add_4_16_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[14] ), .I3(n51659), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_16 (.CI(n51659), .I0(direction_N_3841), 
            .I1(\encoder1_position[14] ), .CO(n51660));
    SB_LUT4 position_1945_add_4_15_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[13] ), .I3(n51658), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_15 (.CI(n51658), .I0(direction_N_3841), 
            .I1(\encoder1_position[13] ), .CO(n51659));
    SB_LUT4 position_1945_add_4_14_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[12] ), .I3(n51657), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_14 (.CI(n51657), .I0(direction_N_3841), 
            .I1(\encoder1_position[12] ), .CO(n51658));
    SB_LUT4 position_1945_add_4_13_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[11] ), .I3(n51656), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_13 (.CI(n51656), .I0(direction_N_3841), 
            .I1(\encoder1_position[11] ), .CO(n51657));
    SB_LUT4 position_1945_add_4_12_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[10] ), .I3(n51655), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_12 (.CI(n51655), .I0(direction_N_3841), 
            .I1(\encoder1_position[10] ), .CO(n51656));
    SB_LUT4 position_1945_add_4_11_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[9] ), .I3(n51654), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_11 (.CI(n51654), .I0(direction_N_3841), 
            .I1(\encoder1_position[9] ), .CO(n51655));
    SB_LUT4 position_1945_add_4_10_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[8] ), .I3(n51653), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_10 (.CI(n51653), .I0(direction_N_3841), 
            .I1(\encoder1_position[8] ), .CO(n51654));
    SB_LUT4 position_1945_add_4_9_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[7] ), .I3(n51652), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_9 (.CI(n51652), .I0(direction_N_3841), 
            .I1(\encoder1_position[7] ), .CO(n51653));
    SB_LUT4 position_1945_add_4_8_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[6] ), .I3(n51651), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_8 (.CI(n51651), .I0(direction_N_3841), 
            .I1(\encoder1_position[6] ), .CO(n51652));
    SB_LUT4 position_1945_add_4_7_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[5] ), .I3(n51650), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_7 (.CI(n51650), .I0(direction_N_3841), 
            .I1(\encoder1_position[5] ), .CO(n51651));
    SB_LUT4 position_1945_add_4_6_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[4] ), .I3(n51649), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF direction_42 (.Q(n1784), .C(n1779), .D(n29664));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_1945_add_4_6 (.CI(n51649), .I0(direction_N_3841), 
            .I1(\encoder1_position[4] ), .CO(n51650));
    SB_LUT4 position_1945_add_4_5_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[3] ), .I3(n51648), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n29656));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_1945_add_4_5 (.CI(n51648), .I0(direction_N_3841), 
            .I1(\encoder1_position[3] ), .CO(n51649));
    SB_LUT4 position_1945_add_4_4_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder1_position[2] ), .I3(n51647), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_4 (.CI(n51647), .I0(direction_N_3841), 
            .I1(\encoder1_position[2] ), .CO(n51648));
    SB_LUT4 position_1945_add_4_3_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1822), .I3(n51646), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_3 (.CI(n51646), .I0(direction_N_3841), 
            .I1(n1822), .CO(n51647));
    SB_LUT4 position_1945_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1824), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1945_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1945_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n1824), 
            .CO(n51646));
    SB_DFFE position_1945__i0 (.Q(n1824), .C(n1779), .E(position_31__N_3837), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i31 (.Q(n1786), .C(n1779), .E(position_31__N_3837), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i30 (.Q(n1788), .C(n1779), .E(position_31__N_3837), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i29 (.Q(n1790), .C(n1779), .E(position_31__N_3837), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i28 (.Q(n1792), .C(n1779), .E(position_31__N_3837), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i27 (.Q(n1794), .C(n1779), .E(position_31__N_3837), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i26 (.Q(n1796), .C(n1779), .E(position_31__N_3837), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i25 (.Q(\encoder1_position[25] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i24 (.Q(\encoder1_position[24] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i23 (.Q(\encoder1_position[23] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i22 (.Q(\encoder1_position[22] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i21 (.Q(\encoder1_position[21] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i20 (.Q(\encoder1_position[20] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i19 (.Q(\encoder1_position[19] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i18 (.Q(\encoder1_position[18] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i17 (.Q(\encoder1_position[17] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i16 (.Q(\encoder1_position[16] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i15 (.Q(\encoder1_position[15] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i14 (.Q(\encoder1_position[14] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i13 (.Q(\encoder1_position[13] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i12 (.Q(\encoder1_position[12] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i11 (.Q(\encoder1_position[11] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i10 (.Q(\encoder1_position[10] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i9 (.Q(\encoder1_position[9] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i8 (.Q(\encoder1_position[8] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i7 (.Q(\encoder1_position[7] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i6 (.Q(\encoder1_position[6] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i5 (.Q(\encoder1_position[5] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i4 (.Q(\encoder1_position[4] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i3 (.Q(\encoder1_position[3] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i2 (.Q(\encoder1_position[2] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1945__i1 (.Q(n1822), .C(n1779), .E(position_31__N_3837), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1779), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1779), .D(b_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29397));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3841));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 debounce_cnt_I_937_4_lut (.I0(a_new_c[0]), .I1(b_new_c[0]), 
            .I2(a_new[1]), .I3(b_new[1]), .O(debounce_cnt_N_3834));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (clk16MHz, enable_slow_N_4214, GND_net, \state[0] , \state_7__N_3919[0] , 
            data_ready, ID, baudrate, n30390, n30389, n30388, n30387, 
            n30386, n30385, n30374, n30373, n30372, n30371, n30370, 
            n30369, n30368, n30367, n114, data, n27922, n48949, 
            n27924, \state_7__N_4111[0] , scl_enable, VCC_net, sda_enable, 
            sda_out, n29653, n29652, n29646, n29645, n29640, n29639, 
            n29637, n6429, n30429, n8, n11, scl, n42234, \state_7__N_4127[3] , 
            n10, n4, n4_adj_26, n25532, n25568, n42355) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output enable_slow_N_4214;
    input GND_net;
    output \state[0] ;
    input \state_7__N_3919[0] ;
    output data_ready;
    output [7:0]ID;
    output [31:0]baudrate;
    input n30390;
    input n30389;
    input n30388;
    input n30387;
    input n30386;
    input n30385;
    input n30374;
    input n30373;
    input n30372;
    input n30371;
    input n30370;
    input n30369;
    input n30368;
    input n30367;
    output n114;
    output [7:0]data;
    output n27922;
    output n48949;
    output n27924;
    output \state_7__N_4111[0] ;
    output scl_enable;
    input VCC_net;
    output sda_enable;
    output sda_out;
    input n29653;
    input n29652;
    input n29646;
    input n29645;
    input n29640;
    input n29639;
    input n29637;
    output n6429;
    input n30429;
    input n8;
    output n11;
    output scl;
    output n42234;
    input \state_7__N_4127[3] ;
    output n10;
    output n4;
    output n4_adj_26;
    output n25532;
    output n25568;
    output n42355;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n29824;
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    
    wire ready_prev;
    wire [0:0]n5723;
    
    wire enable;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n15, n48918, n25437;
    wire [15:0]n5115;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n28, n26, n27, n25, n52335;
    wire [7:0]state_adj_5689;   // verilog/i2c_controller.v(33[12:17])
    
    wire n63535, n66497, n58919, n17, n60624;
    wire [7:0]state_7__N_3886;
    wire [15:0]delay_counter_15__N_3957;
    
    wire n50575, n50574, n50573, n50572, n50571, n6689, n50570, 
        n6688, n50569, n6687, n50568, n6686, n50567, n6685, n50566, 
        n50565, n6683, n50564, n50563, n50562, n50561, n57143, 
        rw, n29624, n29620, n6758;
    wire [1:0]n6492;
    
    wire n60131;
    wire [2:0]n1;
    
    wire n27768, n29082, n52908, n57053, n30405, n30404, n30403, 
        n30402, n30401, n30400, n30399, n30398, n30397, n30396, 
        n30395, n30394, n30393, n30392, n30391, n30384, n30383, 
        n30382, n30381, n30380, n30379, n30378, n30377, n30376, 
        n30375, n37701, n42246, n58903, n47, n42846, n27693, n48930, 
        n29, n52059, n95, n111, n4_c, n4_adj_5683, n28406, n66458, 
        n10_c, n11_c, n10_adj_5684;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n57539;
    
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n29824));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4214));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5723[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n15));   // verilog/eeprom.v(30[11:23])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i18_2_lut (.I0(state[2]), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n48918));
    defparam i18_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i53626_2_lut (.I0(n25437), .I1(enable_slow_N_4214), .I2(GND_net), 
            .I3(GND_net), .O(n5115[13]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i53626_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[5]), .I1(delay_counter[12]), .I2(delay_counter[6]), 
            .I3(delay_counter[10]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[8]), .I1(delay_counter[11]), .I2(delay_counter[9]), 
            .I3(delay_counter[7]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[0]), .I2(delay_counter[13]), 
            .I3(delay_counter[2]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n25437));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(state[0]), .I1(enable_slow_N_4214), .I2(n25437), 
            .I3(GND_net), .O(n52335));
    defparam i2_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i47818_3_lut (.I0(\state[0] ), .I1(n25437), .I2(state_adj_5689[3]), 
            .I3(GND_net), .O(n63535));
    defparam i47818_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n66497), .I1(n58919), .I2(state[0]), .I3(n63535), 
            .O(n17));
    defparam i24_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i2_4_lut (.I0(n17), .I1(state[2]), .I2(\state_7__N_3919[0] ), 
            .I3(state[1]), .O(n60624));
    defparam i2_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i35054_4_lut (.I0(state[1]), .I1(n15), .I2(state[2]), .I3(state[0]), 
            .O(state_7__N_3886[1]));   // verilog/eeprom.v(27[11:16])
    defparam i35054_4_lut.LUT_INIT = 16'ha5ba;
    SB_LUT4 add_1106_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5115[13]), 
            .I3(n50575), .O(delay_counter_15__N_3957[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1106_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5115[13]), 
            .I3(n50574), .O(delay_counter_15__N_3957[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_16 (.CI(n50574), .I0(delay_counter[14]), .I1(n5115[13]), 
            .CO(n50575));
    SB_LUT4 add_1106_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5115[13]), 
            .I3(n50573), .O(delay_counter_15__N_3957[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_15 (.CI(n50573), .I0(delay_counter[13]), .I1(n5115[13]), 
            .CO(n50574));
    SB_LUT4 add_1106_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5115[13]), 
            .I3(n50572), .O(delay_counter_15__N_3957[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_14 (.CI(n50572), .I0(delay_counter[12]), .I1(n5115[13]), 
            .CO(n50573));
    SB_LUT4 add_1106_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5115[13]), 
            .I3(n50571), .O(delay_counter_15__N_3957[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_13 (.CI(n50571), .I0(delay_counter[11]), .I1(n5115[13]), 
            .CO(n50572));
    SB_LUT4 add_1106_12_lut (.I0(n48918), .I1(delay_counter[10]), .I2(n5115[13]), 
            .I3(n50570), .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1106_12 (.CI(n50570), .I0(delay_counter[10]), .I1(n5115[13]), 
            .CO(n50571));
    SB_LUT4 add_1106_11_lut (.I0(n48918), .I1(delay_counter[9]), .I2(n5115[13]), 
            .I3(n50569), .O(n6688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1106_11 (.CI(n50569), .I0(delay_counter[9]), .I1(n5115[13]), 
            .CO(n50570));
    SB_LUT4 add_1106_10_lut (.I0(n48918), .I1(delay_counter[8]), .I2(n5115[13]), 
            .I3(n50568), .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1106_10 (.CI(n50568), .I0(delay_counter[8]), .I1(n5115[13]), 
            .CO(n50569));
    SB_LUT4 add_1106_9_lut (.I0(n48918), .I1(delay_counter[7]), .I2(n5115[13]), 
            .I3(n50567), .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1106_9 (.CI(n50567), .I0(delay_counter[7]), .I1(n5115[13]), 
            .CO(n50568));
    SB_LUT4 add_1106_8_lut (.I0(n48918), .I1(delay_counter[6]), .I2(n5115[13]), 
            .I3(n50566), .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1106_8 (.CI(n50566), .I0(delay_counter[6]), .I1(n5115[13]), 
            .CO(n50567));
    SB_LUT4 add_1106_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5115[13]), 
            .I3(n50565), .O(delay_counter_15__N_3957[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_7 (.CI(n50565), .I0(delay_counter[5]), .I1(n5115[13]), 
            .CO(n50566));
    SB_LUT4 add_1106_6_lut (.I0(n48918), .I1(delay_counter[4]), .I2(n5115[13]), 
            .I3(n50564), .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1106_6 (.CI(n50564), .I0(delay_counter[4]), .I1(n5115[13]), 
            .CO(n50565));
    SB_LUT4 add_1106_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5115[13]), 
            .I3(n50563), .O(delay_counter_15__N_3957[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_5 (.CI(n50563), .I0(delay_counter[3]), .I1(n5115[13]), 
            .CO(n50564));
    SB_LUT4 add_1106_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5115[13]), 
            .I3(n50562), .O(delay_counter_15__N_3957[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_4 (.CI(n50562), .I0(delay_counter[2]), .I1(n5115[13]), 
            .CO(n50563));
    SB_LUT4 add_1106_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5115[13]), 
            .I3(n50561), .O(delay_counter_15__N_3957[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_3 (.CI(n50561), .I0(delay_counter[1]), .I1(n5115[13]), 
            .CO(n50562));
    SB_LUT4 add_1106_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5115[13]), 
            .I3(GND_net), .O(delay_counter_15__N_3957[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1106_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5115[13]), 
            .CO(n50561));
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n57143));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n29624));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29620));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state_adj_5689[3]), .I1(state_adj_5689[2]), 
            .I2(\state[0] ), .I3(GND_net), .O(n6758));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i53655_3_lut_4_lut (.I0(state_adj_5689[3]), .I1(state_adj_5689[2]), 
            .I2(\state[0] ), .I3(state_adj_5689[1]), .O(enable_slow_N_4214));
    defparam i53655_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_4_lut (.I0(state_adj_5689[3]), .I1(state_adj_5689[2]), 
            .I2(n6492[1]), .I3(state_adj_5689[1]), .O(n60131));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_DFFESR byte_counter_1946__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27768), .D(n1[1]), .R(n29082));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1946__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27768), .D(n1[2]), .R(n29082));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1946__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27768), .D(n52908), .R(n29082));   // verilog/eeprom.v(68[25:39])
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n57053));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30405));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30404));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30403));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30402));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30401));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30400));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30399));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30398));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30397));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30396));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30395));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30394));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30393));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30392));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30391));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30390));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30389));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30388));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30387));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n30386));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n30385));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n30384));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n30383));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30382));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30381));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30380));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30379));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30378));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30377));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30376));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30375));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30374));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30373));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30372));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30371));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30370));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30369));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30368));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30367));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n37701));   // verilog/eeprom.v(27[11:16])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28326_2_lut (.I0(enable_slow_N_4214), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n42246));
    defparam i28326_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n60624), .D(state_7__N_3886[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i2_3_lut_4_lut_adj_1760 (.I0(\state[0] ), .I1(state_adj_5689[3]), 
            .I2(n58903), .I3(n25437), .O(n47));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1761 (.I0(\state[0] ), .I1(state_adj_5689[3]), 
            .I2(state_adj_5689[2]), .I3(state_adj_5689[1]), .O(n42846));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_1761.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27693), 
            .D(delay_counter_15__N_3957[1]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27693), 
            .D(delay_counter_15__N_3957[2]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27693), 
            .D(delay_counter_15__N_3957[3]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27693), 
            .D(n6683), .S(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27693), 
            .D(delay_counter_15__N_3957[5]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27693), 
            .D(n6685), .S(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27693), 
            .D(n6686), .S(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27693), 
            .D(n6687), .S(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27693), 
            .D(n6688), .S(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27693), .D(n6689), .S(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27693), .D(delay_counter_15__N_3957[11]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27693), .D(delay_counter_15__N_3957[12]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27693), .D(delay_counter_15__N_3957[13]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27693), .D(delay_counter_15__N_3957[14]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27693), .D(delay_counter_15__N_3957[15]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27693), 
            .D(delay_counter_15__N_3957[0]), .R(n48930));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i16368_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[7]), .I3(ID[7]), 
            .O(n30399));
    defparam i16368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16369_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[6]), .I3(ID[6]), 
            .O(n30400));
    defparam i16369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16370_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[5]), .I3(ID[5]), 
            .O(n30401));
    defparam i16370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16371_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[4]), .I3(ID[4]), 
            .O(n30402));
    defparam i16371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16372_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[3]), .I3(ID[3]), 
            .O(n30403));
    defparam i16372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16373_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[2]), .I3(ID[2]), 
            .O(n30404));
    defparam i16373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16374_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[1]), .I3(ID[1]), 
            .O(n30405));
    defparam i16374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15589_3_lut_4_lut (.I0(n29), .I1(n114), .I2(data[0]), .I3(ID[0]), 
            .O(n29620));
    defparam i15589_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1762 (.I0(byte_counter[1]), .I1(n52059), 
            .I2(n114), .I3(byte_counter[2]), .O(n27922));
    defparam i2_3_lut_4_lut_adj_1762.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_adj_1763 (.I0(byte_counter[1]), .I1(n52059), 
            .I2(byte_counter[2]), .I3(GND_net), .O(n29));
    defparam i1_2_lut_3_lut_adj_1763.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(n37701), .I3(data_ready), 
            .O(n29624));   // verilog/eeprom.v(27[11:16])
    defparam i12_4_lut_4_lut.LUT_INIT = 16'hfa08;
    SB_LUT4 i1_4_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(\state_7__N_3919[0] ), 
            .I3(state[1]), .O(n27768));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h4410;
    SB_LUT4 i2_3_lut_4_lut_adj_1764 (.I0(state[2]), .I1(state[0]), .I2(\state_7__N_3919[0] ), 
            .I3(state[1]), .O(n29082));
    defparam i2_3_lut_4_lut_adj_1764.LUT_INIT = 16'h0010;
    SB_LUT4 i36260_3_lut_4_lut (.I0(n42246), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n1[2]));   // verilog/eeprom.v(68[25:39])
    defparam i36260_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i1_2_lut_3_lut_adj_1765 (.I0(enable_slow_N_4214), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n52908));
    defparam i1_2_lut_3_lut_adj_1765.LUT_INIT = 16'hd2d2;
    SB_LUT4 i43246_2_lut_3_lut (.I0(enable_slow_N_4214), .I1(ready_prev), 
            .I2(state[1]), .I3(GND_net), .O(n58919));
    defparam i43246_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1766 (.I0(n48949), .I1(state[2]), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n27924));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut_adj_1766.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_1767 (.I0(n48949), .I1(state[2]), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n95));   // verilog/eeprom.v(30[11:23])
    defparam i1_2_lut_3_lut_adj_1767.LUT_INIT = 16'hfdfd;
    SB_LUT4 i35049_4_lut_4_lut (.I0(data[7]), .I1(n48949), .I2(n114), 
            .I3(baudrate[15]), .O(n30383));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i35049_4_lut_4_lut.LUT_INIT = 16'hfb08;
    SB_LUT4 i36253_2_lut_3_lut_4_lut (.I0(enable_slow_N_4214), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n1[1]));   // verilog/eeprom.v(68[25:39])
    defparam i36253_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i35039_4_lut (.I0(data[6]), .I1(n95), .I2(baudrate[14]), .I3(n27924), 
            .O(n30384));   // verilog/TinyFPGA_B.v(253[15:23])
    defparam i35039_4_lut.LUT_INIT = 16'heae0;
    SB_LUT4 i2_3_lut_adj_1768 (.I0(byte_counter[2]), .I1(n52059), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n48949));
    defparam i2_3_lut_adj_1768.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_adj_1769 (.I0(state[2]), .I1(byte_counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n111));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_adj_1769.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(n15), .O(n27693));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h1416;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(n15), .O(n48930));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h1012;
    SB_LUT4 i1_2_lut_adj_1770 (.I0(\state_7__N_3919[0] ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_1770.LUT_INIT = 16'heeee;
    SB_LUT4 i53561_3_lut (.I0(n47), .I1(n42246), .I2(state[0]), .I3(GND_net), 
            .O(n4_adj_5683));
    defparam i53561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1771 (.I0(state[1]), .I1(state[2]), .I2(n4_adj_5683), 
            .I3(n4_c), .O(n28406));
    defparam i2_4_lut_adj_1771.LUT_INIT = 16'hecfd;
    SB_LUT4 i51141_3_lut (.I0(n28406), .I1(state[2]), .I2(\state_7__N_3919[0] ), 
            .I3(GND_net), .O(n66458));   // verilog/eeprom.v(27[11:16])
    defparam i51141_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i28_4_lut (.I0(n66458), .I1(n47), .I2(state[1]), .I3(n28406), 
            .O(n10_c));   // verilog/eeprom.v(27[11:16])
    defparam i28_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i27_4_lut (.I0(n10_c), .I1(n58919), .I2(state[0]), .I3(state[2]), 
            .O(n57053));   // verilog/eeprom.v(27[11:16])
    defparam i27_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(state_adj_5689[3]), 
            .I1(state_adj_5689[2]), .I2(\state[0] ), .I3(state_adj_5689[1]), 
            .O(n11_c));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(n42246), .O(n29824));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'ha8e8;
    SB_LUT4 i50827_2_lut_3_lut (.I0(state_adj_5689[2]), .I1(state_adj_5689[1]), 
            .I2(state[1]), .I3(GND_net), .O(n66497));
    defparam i50827_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 mux_1433_Mux_0_i3_3_lut_4_lut (.I0(state[0]), .I1(enable_slow_N_4214), 
            .I2(n25437), .I3(state[1]), .O(n5723[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1433_Mux_0_i3_3_lut_4_lut.LUT_INIT = 16'h04aa;
    SB_LUT4 i16367_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[0]), .I3(baudrate[0]), 
            .O(n30398));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16367_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16360_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[7]), .I3(baudrate[7]), 
            .O(n30391));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16360_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16361_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[6]), .I3(baudrate[6]), 
            .O(n30392));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16361_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16362_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[5]), .I3(baudrate[5]), 
            .O(n30393));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16362_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16363_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[4]), .I3(baudrate[4]), 
            .O(n30394));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16363_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16364_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[3]), .I3(baudrate[3]), 
            .O(n30395));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16364_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16365_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[2]), .I3(baudrate[2]), 
            .O(n30396));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16365_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16366_3_lut_4_lut (.I0(n29), .I1(n111), .I2(data[1]), .I3(baudrate[1]), 
            .O(n30397));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16366_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16351_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[0]), 
            .I3(baudrate[16]), .O(n30382));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16344_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[7]), 
            .I3(baudrate[23]), .O(n30375));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16344_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16345_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[6]), 
            .I3(baudrate[22]), .O(n30376));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16346_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[5]), 
            .I3(baudrate[21]), .O(n30377));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16347_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[4]), 
            .I3(baudrate[20]), .O(n30378));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16348_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[3]), 
            .I3(baudrate[19]), .O(n30379));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16349_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[2]), 
            .I3(baudrate[18]), .O(n30380));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16350_3_lut_4_lut (.I0(n48949), .I1(n111), .I2(data[1]), 
            .I3(baudrate[17]), .O(n30381));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut (.I0(ready_prev), .I1(n42846), .I2(state[0]), .I3(state[1]), 
            .O(n52059));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_adj_1772 (.I0(state[2]), .I1(byte_counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n114));
    defparam i1_2_lut_adj_1772.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(rw), .I2(n52335), .I3(state[2]), 
            .O(n10_adj_5684));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut.LUT_INIT = 16'h888a;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n10_adj_5684), .I1(rw), .I2(state[0]), 
            .I3(state[2]), .O(n57143));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'heeae;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n42846), .I1(saved_addr[0]), .I2(rw), 
            .I3(\state_7__N_4111[0] ), .O(n57539));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hd8cc;
    i2c_controller i2c (.clk16MHz(clk16MHz), .scl_enable(scl_enable), .\state_7__N_4111[0] (\state_7__N_4111[0] ), 
            .\state[2] (state_adj_5689[2]), .\state[1] (state_adj_5689[1]), 
            .n58903(n58903), .GND_net(GND_net), .VCC_net(VCC_net), .sda_enable(sda_enable), 
            .sda_out(sda_out), .n29653(n29653), .data({data}), .n29652(n29652), 
            .n29646(n29646), .n29645(n29645), .n29640(n29640), .n29639(n29639), 
            .n29637(n29637), .n57539(n57539), .\saved_addr[0] (saved_addr[0]), 
            .n6429(n6429), .\state[3] (state_adj_5689[3]), .n30429(n30429), 
            .n8(n8), .\state[0] (\state[0] ), .n60131(n60131), .enable_slow_N_4214(enable_slow_N_4214), 
            .n11(n11), .enable(enable), .scl(scl), .n42234(n42234), 
            .\state_7__N_4127[3] (\state_7__N_4127[3] ), .n11_adj_24(n11_c), 
            .n10(n10), .n6758(n6758), .sda_out_N_4209(n6492[1]), .n4(n4), 
            .n4_adj_25(n4_adj_26), .n25532(n25532), .n25568(n25568), .n42355(n42355)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (clk16MHz, scl_enable, \state_7__N_4111[0] , \state[2] , 
            \state[1] , n58903, GND_net, VCC_net, sda_enable, sda_out, 
            n29653, data, n29652, n29646, n29645, n29640, n29639, 
            n29637, n57539, \saved_addr[0] , n6429, \state[3] , n30429, 
            n8, \state[0] , n60131, enable_slow_N_4214, n11, enable, 
            scl, n42234, \state_7__N_4127[3] , n11_adj_24, n10, n6758, 
            sda_out_N_4209, n4, n4_adj_25, n25532, n25568, n42355) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output scl_enable;
    output \state_7__N_4111[0] ;
    output \state[2] ;
    output \state[1] ;
    output n58903;
    input GND_net;
    input VCC_net;
    output sda_enable;
    output sda_out;
    input n29653;
    output [7:0]data;
    input n29652;
    input n29646;
    input n29645;
    input n29640;
    input n29639;
    input n29637;
    input n57539;
    output \saved_addr[0] ;
    output n6429;
    output \state[3] ;
    input n30429;
    input n8;
    output \state[0] ;
    input n60131;
    input enable_slow_N_4214;
    output n11;
    input enable;
    output scl;
    output n42234;
    input \state_7__N_4127[3] ;
    input n11_adj_24;
    output n10;
    input n6758;
    output sda_out_N_4209;
    output n4;
    output n4_adj_25;
    output n25532;
    output n25568;
    output n42355;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire i2c_clk_N_4200, scl_enable_N_4201, enable_slow_N_4213, n27752;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n29060;
    wire [7:0]n119;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n50582, n50581, sda_out_adj_5670, n50580, n50579, n50578, 
        n50577, n50576;
    wire [5:0]n29;
    
    wire n27831, n28823, n5, n42759, n42506, n42757, n61159, n59916, 
        n11_c, n60981, n27751, n57265, n27749, n51709, n51708, 
        n51707, n51706, n51705, n11_adj_5671, n42842, n4_c, n9, 
        n15, n11_adj_5673, n6422, n9_adj_5675, n12, n4_adj_5677, 
        n66498, n28, n69308, n58895;
    
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4200));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4201));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4111[0] ), .C(clk16MHz), .E(n27752), 
            .D(enable_slow_N_4213));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i43230_2_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n58903));
    defparam i43230_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n29060));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29060), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4200));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n50582), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n50581), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2428_2_lut (.I0(sda_out_adj_5670), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2428_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_39_add_2_8 (.CI(n50581), .I0(counter[6]), .I1(VCC_net), 
            .CO(n50582));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n50580), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n50580), .I0(counter[5]), .I1(VCC_net), 
            .CO(n50581));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n50579), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n50579), .I0(counter[4]), .I1(VCC_net), 
            .CO(n50580));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n50578), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n50578), .I0(counter[3]), .I1(VCC_net), 
            .CO(n50579));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n50577), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n50577), .I0(counter[2]), .I1(VCC_net), 
            .CO(n50578));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n50576), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n50576), .I0(counter[1]), .I1(VCC_net), 
            .CO(n50577));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n50576));
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29653));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29652));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29646));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29645));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29640));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29639));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29637));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n57539));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1955_1956__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29060));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1955_1956__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29060));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1955_1956__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29060));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1955_1956__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29060));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1955_1956__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29060));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27831), .D(n119[1]), 
            .S(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27831), .D(n119[2]), 
            .S(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27831), .D(n119[3]), 
            .R(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27831), .D(n119[4]), 
            .R(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27831), .D(n119[5]), 
            .R(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27831), .D(n119[6]), 
            .R(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27831), .D(n119[7]), 
            .R(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6429), .D(n5), 
            .S(n42759));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6429), .D(n42506), 
            .S(n42757));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6429), .D(n61159), 
            .S(n59916));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1955_1956__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29060));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30429));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i54174_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6429), 
            .I3(\state[1] ), .O(n59916));   // verilog/i2c_controller.v(130[5:15])
    defparam i54174_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 equal_1520_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_c));   // verilog/i2c_controller.v(130[5:15])
    defparam equal_1520_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hdfff;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27751), 
            .D(n60981), .S(n57265));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_5670), .C(i2c_clk), .E(n27749), 
            .D(n60131), .S(n57265));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27831), .D(n119[0]), 
            .S(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_1955_1956_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n51709), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1955_1956_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1955_1956_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n51708), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1955_1956_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1955_1956_add_4_6 (.CI(n51708), .I0(GND_net), .I1(counter2[4]), 
            .CO(n51709));
    SB_LUT4 counter2_1955_1956_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n51707), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1955_1956_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1955_1956_add_4_5 (.CI(n51707), .I0(GND_net), .I1(counter2[3]), 
            .CO(n51708));
    SB_LUT4 counter2_1955_1956_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n51706), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1955_1956_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1955_1956_add_4_4 (.CI(n51706), .I0(GND_net), .I1(counter2[2]), 
            .CO(n51707));
    SB_LUT4 counter2_1955_1956_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n51705), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1955_1956_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1955_1956_add_4_3 (.CI(n51705), .I0(GND_net), .I1(counter2[1]), 
            .CO(n51706));
    SB_LUT4 counter2_1955_1956_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1955_1956_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1955_1956_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n51705));
    SB_LUT4 i53658_2_lut (.I0(enable_slow_N_4214), .I1(\state_7__N_4111[0] ), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(44[32:47])
    defparam i53658_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_5671));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i28920_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(GND_net), .O(n42842));
    defparam i28920_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9), .O(n61159));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf0f4;
    SB_LUT4 i2_3_lut_4_lut_adj_1752 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n60981));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_1752.LUT_INIT = 16'h1110;
    SB_LUT4 i14792_2_lut_4_lut (.I0(n27831), .I1(\state[3] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n28823));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14792_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(enable_slow_N_4214), .I2(\state_7__N_4111[0] ), 
            .I3(GND_net), .O(n27752));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i28347_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i28347_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28314_3_lut_4_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n42234));   // verilog/i2c_controller.v(130[5:15])
    defparam i28314_3_lut_4_lut_4_lut.LUT_INIT = 16'hfcfd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n15));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5673));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut (.I0(\state_7__N_4127[3] ), .I1(n11_adj_5671), .I2(n11_c), 
            .I3(enable), .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'h2a2f;
    SB_LUT4 i54182_3_lut (.I0(n6429), .I1(n15), .I2(n11), .I3(GND_net), 
            .O(n42757));
    defparam i54182_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i54150_2_lut (.I0(\state_7__N_4127[3] ), .I1(n11_adj_5671), 
            .I2(GND_net), .I3(GND_net), .O(n42506));
    defparam i54150_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i54183_4_lut (.I0(n6429), .I1(\state[0] ), .I2(n11_adj_24), 
            .I3(n58903), .O(n42759));
    defparam i54183_4_lut.LUT_INIT = 16'h0a8a;
    SB_LUT4 i53606_4_lut (.I0(\state[3] ), .I1(n6422), .I2(n42842), .I3(n42234), 
            .O(n6429));
    defparam i53606_4_lut.LUT_INIT = 16'h5f13;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n11_adj_5673), .I1(n11_adj_5671), .I2(\saved_addr[0] ), 
            .I3(\state_7__N_4127[3] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'h5575;
    SB_LUT4 equal_273_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5675));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_273_i9_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6422));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1754 (.I0(\state[3] ), .I1(n6422), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5677));
    defparam i1_2_lut_adj_1754.LUT_INIT = 16'hbbbb;
    SB_LUT4 i50828_4_lut (.I0(n58903), .I1(n4_adj_5677), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n66498));
    defparam i50828_4_lut.LUT_INIT = 16'hfcdd;
    SB_LUT4 i14_4_lut (.I0(n66498), .I1(n9_adj_5675), .I2(n6758), .I3(\state_7__N_4127[3] ), 
            .O(n27831));
    defparam i14_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'h5110;
    SB_LUT4 i53582_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n69308));
    defparam i53582_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n11_c), .I1(n69308), .I2(n28), .I3(n58895), 
            .O(n27749));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1732_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(sda_out_N_4209));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1732_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i29039_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n58895));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i29039_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[0] ), .I1(n58903), .I2(\state[3] ), .I3(n11_c), 
            .O(n57265));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n11_c), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n58895), .O(n27751));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'h0a22;
    SB_LUT4 i43331_3_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[1] ), 
            .I3(\state[3] ), .O(scl_enable_N_4201));
    defparam i43331_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_352_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_352_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_350_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_25));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_350_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1758 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n25532));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_1758.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1759 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n25568));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_1759.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28433_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n42355));
    defparam i28433_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n29606, \data_in_frame[4] , clk16MHz, n29891, VCC_net, 
            \data_in_frame[7] , GND_net, \data_out_frame[20] , \data_out_frame[22] , 
            n29888, \data_in_frame[6] , \data_out_frame[21] , n2874, 
            \data_out_frame[8] , n57860, n57859, n29885, \data_in_frame[8] , 
            \data_out_frame[24] , \data_out_frame[25] , \data_out_frame[19] , 
            \data_out_frame[15] , \data_out_frame[17] , \data_out_frame[18] , 
            n58651, \data_out_frame[13] , \data_out_frame[23] , n58570, 
            n25705, \FRAME_MATCHER.state[3] , \data_out_frame[12] , \data_out_frame[16] , 
            \FRAME_MATCHER.i_31__N_2509 , pwm_setpoint, \data_out_frame[10] , 
            \data_out_frame[5] , current_limit, n22773, \data_out_frame[14] , 
            \data_out_frame[11] , \data_out_frame[7] , \data_out_frame[9] , 
            \data_out_frame[6] , n58099, \data_out_frame[4] , n25676, 
            n29881, n29878, n29875, n29872, n29869, n29866, n29863, 
            n29860, n29857, \data_in_frame[5] , n29854, n29851, n29848, 
            n29621, n29844, \data_in_frame[0] , n29841, n29838, n26306, 
            n29818, n25666, n34, \data_in_frame[0][5] , n26111, n2076, 
            encoder1_position_scaled, displacement, n15, n15_adj_7, 
            \data_in_frame[3] , \data_in_frame[2][1] , \data_in_frame[0][0] , 
            \data_in_frame[2][5] , \data_in_frame[3][0] , n58498, \data_in_frame[1] , 
            \data_in_frame[3][7] , n29641, neopxl_color, n29657, n58075, 
            encoder0_position_scaled, \data_in_frame[1][6] , n29813, n57858, 
            \data_in_frame[1][7] , \data_in_frame[8][3] , n57857, reset, 
            setpoint, \data_in_frame[1][2] , deadband, \data_in_frame[2][0] , 
            \data_in_frame[3][5] , n29698, \data_in_frame[2][3] , n57900, 
            control_mode, n57856, \data_in_frame[8][6] , \control_mode[1] , 
            \data_in_frame[20][4] , \control_mode[0] , \data_in_frame[21][2] , 
            \data_in_frame[21][3] , \data_in_frame[18] , n57863, n57855, 
            n57854, n57853, n57852, n57851, n57850, n28997, n57849, 
            n57848, n57847, n57846, n57845, n57844, n57843, n57842, 
            \data_in_frame[22][5] , \data_in_frame[20][3] , \data_in_frame[22][4] , 
            \data_in_frame[20][0] , \data_in_frame[21][1] , \data_in_frame[21][5] , 
            \data_in_frame[19] , \data_in_frame[22][1] , n28988, n57841, 
            n57840, n57839, n57838, n57837, n57836, n57835, \data_in_frame[22][7] , 
            n57834, n57833, n57832, n57831, n57830, n57829, n57828, 
            \data_in_frame[17] , \data_in_frame[22][2] , n57827, \data_in_frame[20][1] , 
            \data_in_frame[22][3] , n57826, n57825, n57824, n57823, 
            \o_Rx_DV_N_3488[12] , n4942, \o_Rx_DV_N_3488[24] , n29, 
            n23, n27, \r_SM_Main_2__N_3536[1] , n57822, n57821, n57820, 
            \byte_transmit_counter[2] , n37407, n57819, n57818, n57817, 
            n57734, n57816, n28960, \data_out_frame[1][1] , \data_out_frame[3][1] , 
            \byte_transmit_counter[0] , n57815, n29703, n57814, IntegralLimit, 
            n57813, \FRAME_MATCHER.i[0] , ID, \Kp[1] , \Kp[2] , \Kp[3] , 
            \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , n29709, 
            \Kp[15] , \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , 
            \Ki[6] , \Ki[7] , n8, \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , 
            \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , n29729, n29728, 
            n29727, n29726, n29725, n29724, n29723, n29722, n29721, 
            n29720, n150, n36515, n29719, n29718, n29717, n29716, 
            n29715, n29714, n58897, n29713, n29712, n29708, n29702, 
            \FRAME_MATCHER.rx_data_ready_prev , \data_out_frame[3][7] , 
            n29701, n29697, \current_limit[2] , \data_out_frame[3][6] , 
            \data_out_frame[3][4] , PWMLimit, \data_out_frame[3][3] , 
            n57812, n57811, n57810, n57809, rx_data, n58929, n57808, 
            n57807, n57806, n57805, n29677, \current_limit[12] , n57804, 
            n57803, n29676, \current_limit[11] , n29674, \current_limit[9] , 
            n29673, \current_limit[8] , n29671, \current_limit[7] , 
            n57735, n57736, n57737, n57738, n29669, \current_limit[5] , 
            n57739, n29666, \current_limit[3] , n57740, \data_out_frame[1][7] , 
            n28940, \data_out_frame[1][6] , n29655, n29654, n57741, 
            n57742, n57743, n29651, n29650, n57744, n57745, n29630, 
            n7, n57746, n57747, n30552, n28932, n57748, n8_adj_8, 
            n29617, \current_limit[0] , n29615, \Ki[0] , \Kp[0] , 
            n57749, n57750, n57751, n57752, n57753, n57754, n30561, 
            n28924, n57755, n57756, n57757, n57758, n57759, n57760, 
            n30568, n28917, n41, n57761, n57762, n57763, n25, 
            n28911, n28910, n57764, n57765, n57766, n57767, n57768, 
            n57769, n57770, n57771, n57772, n57773, n57774, n57775, 
            n57776, n57777, n57778, n57779, \data_out_frame[0][2] , 
            n28893, rx_data_ready, n57899, \data_out_frame[0][3] , n57898, 
            n58008, n30452, \current_limit[4] , n30441, n57237, \data_in_frame[18][3] , 
            n57235, \data_in_frame[18][4] , n57233, n8_adj_9, n58010, 
            n57229, \data_in_frame[18][7] , n29385, n29388, n57179, 
            \data_in_frame[18][1] , n29895, n29391, n29394, n29404, 
            \data_in_frame[0][4] , n29898, n29901, n29410, n29413, 
            n57183, \data_in_frame[18][0] , n29442, n57383, \data_in_frame[9][7] , 
            \data_in_frame[11][2] , \data_in_frame[12] , \data_out_frame[1][5] , 
            n58011, n57225, \data_in_frame[16] , n57223, n57221, n57219, 
            n57215, n57211, n57207, n57203, n30149, n58009, n57199, 
            \data_in_frame[17][3] , n57195, \data_in_frame[17][4] , n57191, 
            \data_in_frame[17][5] , n30169, \data_in_frame[17][6] , n57187, 
            n57117, \data_in_frame[21][0] , n57169, n57167, n57163, 
            n57159, \data_in_frame[21][4] , n57155, \data_in_frame[21][7] , 
            n29502, n29505, n29508, n29511, n29514, n29520, \data_out_frame[0][4] , 
            n57897, n29538, n29541, \data_out_frame[1][0] , n57896, 
            n29560, n57895, n29566, \data_out_frame[1][3] , n57894, 
            n57893, n29575, n29578, n29581, \data_in_frame[3][2] , 
            n29584, n57892, n57891, n29592, n57890, n57889, n57888, 
            n57887, n57886, n57885, n57884, n29600, n29423, n40525, 
            n28352, n57883, n57882, n57881, n57880, n57879, LED_c, 
            n29603, n30680, n29037, n57780, n57781, n57782, n28355, 
            n57783, n57878, n30686, n29035, n30687, n29034, n57877, 
            n30689, n29032, n57876, n30691, n29030, n57875, n57874, 
            n57873, n57872, n57871, n57870, n57869, n57868, n57867, 
            n57866, n57865, n57864, n29403, n57784, n29401, \current_limit[1] , 
            n57785, n57786, n57787, n57788, n57789, n57790, n57791, 
            n57792, n57793, n57794, n57795, n57796, n30717, n29017, 
            n30718, n29016, n30719, n29015, n57862, n57797, n57733, 
            n57798, n57799, n57800, n57801, n57802, DE_c, n26, 
            n18, n28363, n30778, n29013, n30779, n29012, n57861, 
            \current[15] , n260, n58520, n28358, n28338, n15_adj_10, 
            n25961, Kp_23__N_1301, n58561, n8_adj_11, n58766, n17, 
            n18_adj_12, \motor_state_23__N_91[1] , \motor_state[1] , \motor_state_23__N_91[2] , 
            \motor_state[2] , \motor_state_23__N_91[3] , \motor_state[3] , 
            \motor_state_23__N_91[4] , \motor_state[4] , \motor_state_23__N_91[5] , 
            \motor_state[5] , \motor_state_23__N_91[6] , \motor_state[6] , 
            \motor_state_23__N_91[7] , \motor_state[7] , n28361, n10, 
            \motor_state_23__N_91[9] , \motor_state[9] , \motor_state_23__N_91[10] , 
            \motor_state[10] , \motor_state_23__N_91[11] , \motor_state[11] , 
            \motor_state_23__N_91[12] , \motor_state[12] , \motor_state_23__N_91[13] , 
            \motor_state[13] , \motor_state_23__N_91[14] , \motor_state[14] , 
            n7_adj_13, \motor_state_23__N_91[21] , \motor_state[21] , 
            n28304, \motor_state_23__N_91[17] , \motor_state[17] , n53323, 
            \motor_state_23__N_91[19] , \motor_state[19] , \motor_state_23__N_91[20] , 
            \motor_state[20] , n25771, \current[7] , \motor_state_23__N_91[22] , 
            \motor_state[22] , \motor_state_23__N_91[23] , \motor_state[23] , 
            n7_adj_14, \motor_state_23__N_91[15] , \motor_state[15] , 
            \motor_state_23__N_91[18] , \motor_state[18] , n58169, n58405, 
            n58556, \current[6] , \current[5] , \current[4] , \current[3] , 
            \current[2] , \current[1] , \current[0] , \current[11] , 
            \current[10] , \current[9] , \current[8] , n22760, n52894, 
            n14, n58366, n66452, n58711, n25819, n26235, n26405, 
            n70252, n58046, n63899, n63900, n60683, n69300, n60931, 
            n63903, n63902, tx_o, r_Clock_Count, tx_enable, baudrate, 
            n27845, n58988, \r_SM_Main[2] , r_Rx_Data, RX_N_2, r_Clock_Count_adj_23, 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[8] , \o_Rx_DV_N_3488[7] , n61478, \r_SM_Main_2__N_3446[1] , 
            \r_SM_Main[1] , n4939, n25566, n29596, n29595, n29591, 
            n29590, n29559, n29558, n29557, \r_Bit_Index[0] , n61043, 
            n30440, n53943, n30436, \o_Rx_DV_N_3488[0] , n61750, n61702, 
            n61734, n61814, n61782, n61766, n61798, n61718, n57927, 
            n27722) /* synthesis syn_module_defined=1 */ ;
    input n29606;
    output [7:0]\data_in_frame[4] ;
    input clk16MHz;
    input n29891;
    input VCC_net;
    output [7:0]\data_in_frame[7] ;
    input GND_net;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[22] ;
    input n29888;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_out_frame[21] ;
    input n2874;
    output [7:0]\data_out_frame[8] ;
    input n57860;
    input n57859;
    input n29885;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output n58651;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[23] ;
    output n58570;
    input n25705;
    output \FRAME_MATCHER.state[3] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[16] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]pwm_setpoint;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[5] ;
    output [15:0]current_limit;
    output n22773;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[6] ;
    output n58099;
    output [7:0]\data_out_frame[4] ;
    output n25676;
    input n29881;
    input n29878;
    input n29875;
    input n29872;
    input n29869;
    input n29866;
    input n29863;
    input n29860;
    input n29857;
    output [7:0]\data_in_frame[5] ;
    input n29854;
    input n29851;
    input n29848;
    input n29621;
    input n29844;
    output [7:0]\data_in_frame[0] ;
    input n29841;
    input n29838;
    output n26306;
    input n29818;
    output n25666;
    input n34;
    output \data_in_frame[0][5] ;
    output n26111;
    output n2076;
    input [23:0]encoder1_position_scaled;
    input [23:0]displacement;
    output n15;
    input n15_adj_7;
    output [7:0]\data_in_frame[3] ;
    output \data_in_frame[2][1] ;
    output \data_in_frame[0][0] ;
    output \data_in_frame[2][5] ;
    output \data_in_frame[3][0] ;
    input n58498;
    output [7:0]\data_in_frame[1] ;
    output \data_in_frame[3][7] ;
    input n29641;
    output [23:0]neopxl_color;
    input n29657;
    output n58075;
    input [23:0]encoder0_position_scaled;
    output \data_in_frame[1][6] ;
    input n29813;
    input n57858;
    output \data_in_frame[1][7] ;
    output \data_in_frame[8][3] ;
    input n57857;
    input reset;
    output [23:0]setpoint;
    output \data_in_frame[1][2] ;
    output [23:0]deadband;
    output \data_in_frame[2][0] ;
    output \data_in_frame[3][5] ;
    input n29698;
    output \data_in_frame[2][3] ;
    input n57900;
    output [7:0]control_mode;
    input n57856;
    output \data_in_frame[8][6] ;
    output \control_mode[1] ;
    output \data_in_frame[20][4] ;
    output \control_mode[0] ;
    output \data_in_frame[21][2] ;
    output \data_in_frame[21][3] ;
    output [7:0]\data_in_frame[18] ;
    input n57863;
    input n57855;
    input n57854;
    input n57853;
    input n57852;
    input n57851;
    input n57850;
    input n28997;
    input n57849;
    input n57848;
    input n57847;
    input n57846;
    input n57845;
    input n57844;
    input n57843;
    input n57842;
    output \data_in_frame[22][5] ;
    output \data_in_frame[20][3] ;
    output \data_in_frame[22][4] ;
    output \data_in_frame[20][0] ;
    output \data_in_frame[21][1] ;
    output \data_in_frame[21][5] ;
    output [7:0]\data_in_frame[19] ;
    output \data_in_frame[22][1] ;
    input n28988;
    input n57841;
    input n57840;
    input n57839;
    input n57838;
    input n57837;
    input n57836;
    input n57835;
    output \data_in_frame[22][7] ;
    input n57834;
    input n57833;
    input n57832;
    input n57831;
    input n57830;
    input n57829;
    input n57828;
    output [7:0]\data_in_frame[17] ;
    output \data_in_frame[22][2] ;
    input n57827;
    output \data_in_frame[20][1] ;
    output \data_in_frame[22][3] ;
    input n57826;
    input n57825;
    input n57824;
    input n57823;
    output \o_Rx_DV_N_3488[12] ;
    input n4942;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    output n27;
    input \r_SM_Main_2__N_3536[1] ;
    input n57822;
    input n57821;
    input n57820;
    output \byte_transmit_counter[2] ;
    output n37407;
    input n57819;
    input n57818;
    input n57817;
    input n57734;
    input n57816;
    input n28960;
    output \data_out_frame[1][1] ;
    output \data_out_frame[3][1] ;
    output \byte_transmit_counter[0] ;
    input n57815;
    input n29703;
    input n57814;
    output [23:0]IntegralLimit;
    input n57813;
    output \FRAME_MATCHER.i[0] ;
    input [7:0]ID;
    output \Kp[1] ;
    output \Kp[2] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output \Kp[5] ;
    output \Kp[6] ;
    output \Kp[7] ;
    output \Kp[8] ;
    output \Kp[9] ;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    output \Kp[13] ;
    output \Kp[14] ;
    input n29709;
    output \Kp[15] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output n8;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    output \Ki[14] ;
    output \Ki[15] ;
    input n29729;
    input n29728;
    input n29727;
    input n29726;
    input n29725;
    input n29724;
    input n29723;
    input n29722;
    input n29721;
    input n29720;
    input n150;
    output n36515;
    input n29719;
    input n29718;
    input n29717;
    input n29716;
    input n29715;
    input n29714;
    output n58897;
    input n29713;
    input n29712;
    input n29708;
    input n29702;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output \data_out_frame[3][7] ;
    input n29701;
    input n29697;
    output \current_limit[2] ;
    output \data_out_frame[3][6] ;
    output \data_out_frame[3][4] ;
    output [23:0]PWMLimit;
    output \data_out_frame[3][3] ;
    input n57812;
    input n57811;
    input n57810;
    input n57809;
    output [7:0]rx_data;
    output n58929;
    input n57808;
    input n57807;
    input n57806;
    input n57805;
    input n29677;
    output \current_limit[12] ;
    input n57804;
    input n57803;
    input n29676;
    output \current_limit[11] ;
    input n29674;
    output \current_limit[9] ;
    input n29673;
    output \current_limit[8] ;
    input n29671;
    output \current_limit[7] ;
    input n57735;
    input n57736;
    input n57737;
    input n57738;
    input n29669;
    output \current_limit[5] ;
    input n57739;
    input n29666;
    output \current_limit[3] ;
    input n57740;
    output \data_out_frame[1][7] ;
    input n28940;
    output \data_out_frame[1][6] ;
    input n29655;
    input n29654;
    input n57741;
    input n57742;
    input n57743;
    input n29651;
    input n29650;
    input n57744;
    input n57745;
    input n29630;
    output n7;
    input n57746;
    input n57747;
    input n30552;
    input n28932;
    input n57748;
    output n8_adj_8;
    input n29617;
    output \current_limit[0] ;
    input n29615;
    output \Ki[0] ;
    output \Kp[0] ;
    input n57749;
    input n57750;
    input n57751;
    input n57752;
    input n57753;
    input n57754;
    input n30561;
    input n28924;
    input n57755;
    input n57756;
    input n57757;
    input n57758;
    input n57759;
    input n57760;
    input n30568;
    input n28917;
    input n41;
    input n57761;
    input n57762;
    input n57763;
    input n25;
    input n28911;
    input n28910;
    input n57764;
    input n57765;
    input n57766;
    input n57767;
    input n57768;
    input n57769;
    input n57770;
    input n57771;
    input n57772;
    input n57773;
    input n57774;
    input n57775;
    input n57776;
    input n57777;
    input n57778;
    input n57779;
    output \data_out_frame[0][2] ;
    input n28893;
    output rx_data_ready;
    input n57899;
    output \data_out_frame[0][3] ;
    input n57898;
    output n58008;
    input n30452;
    output \current_limit[4] ;
    input n30441;
    input n57237;
    output \data_in_frame[18][3] ;
    input n57235;
    output \data_in_frame[18][4] ;
    input n57233;
    output n8_adj_9;
    output n58010;
    input n57229;
    output \data_in_frame[18][7] ;
    input n29385;
    input n29388;
    input n57179;
    output \data_in_frame[18][1] ;
    input n29895;
    input n29391;
    input n29394;
    input n29404;
    output \data_in_frame[0][4] ;
    input n29898;
    input n29901;
    input n29410;
    input n29413;
    input n57183;
    output \data_in_frame[18][0] ;
    input n29442;
    input n57383;
    output \data_in_frame[9][7] ;
    output \data_in_frame[11][2] ;
    output [7:0]\data_in_frame[12] ;
    output \data_out_frame[1][5] ;
    output n58011;
    input n57225;
    output [7:0]\data_in_frame[16] ;
    input n57223;
    input n57221;
    input n57219;
    input n57215;
    input n57211;
    input n57207;
    input n57203;
    input n30149;
    output n58009;
    input n57199;
    output \data_in_frame[17][3] ;
    input n57195;
    output \data_in_frame[17][4] ;
    input n57191;
    output \data_in_frame[17][5] ;
    input n30169;
    output \data_in_frame[17][6] ;
    input n57187;
    input n57117;
    output \data_in_frame[21][0] ;
    input n57169;
    input n57167;
    input n57163;
    input n57159;
    output \data_in_frame[21][4] ;
    input n57155;
    output \data_in_frame[21][7] ;
    input n29502;
    input n29505;
    input n29508;
    input n29511;
    input n29514;
    input n29520;
    output \data_out_frame[0][4] ;
    input n57897;
    input n29538;
    input n29541;
    output \data_out_frame[1][0] ;
    input n57896;
    input n29560;
    input n57895;
    input n29566;
    output \data_out_frame[1][3] ;
    input n57894;
    input n57893;
    input n29575;
    input n29578;
    input n29581;
    output \data_in_frame[3][2] ;
    input n29584;
    input n57892;
    input n57891;
    input n29592;
    input n57890;
    input n57889;
    input n57888;
    input n57887;
    input n57886;
    input n57885;
    input n57884;
    input n29600;
    input n29423;
    output n40525;
    output n28352;
    input n57883;
    input n57882;
    input n57881;
    input n57880;
    input n57879;
    output LED_c;
    input n29603;
    input n30680;
    input n29037;
    input n57780;
    input n57781;
    input n57782;
    input n28355;
    input n57783;
    input n57878;
    input n30686;
    input n29035;
    input n30687;
    input n29034;
    input n57877;
    input n30689;
    input n29032;
    input n57876;
    input n30691;
    input n29030;
    input n57875;
    input n57874;
    input n57873;
    input n57872;
    input n57871;
    input n57870;
    input n57869;
    input n57868;
    input n57867;
    input n57866;
    input n57865;
    input n57864;
    input n29403;
    input n57784;
    input n29401;
    output \current_limit[1] ;
    input n57785;
    input n57786;
    input n57787;
    input n57788;
    input n57789;
    input n57790;
    input n57791;
    input n57792;
    input n57793;
    input n57794;
    input n57795;
    input n57796;
    input n30717;
    input n29017;
    input n30718;
    input n29016;
    input n30719;
    input n29015;
    input n57862;
    input n57797;
    input n57733;
    input n57798;
    input n57799;
    input n57800;
    input n57801;
    input n57802;
    output DE_c;
    input n26;
    output n18;
    input n28363;
    input n30778;
    input n29013;
    input n30779;
    input n29012;
    input n57861;
    input \current[15] ;
    output n260;
    output n58520;
    output n28358;
    output n28338;
    output n15_adj_10;
    output n25961;
    input Kp_23__N_1301;
    input n58561;
    output n8_adj_11;
    input n58766;
    input n17;
    output n18_adj_12;
    input \motor_state_23__N_91[1] ;
    output \motor_state[1] ;
    input \motor_state_23__N_91[2] ;
    output \motor_state[2] ;
    input \motor_state_23__N_91[3] ;
    output \motor_state[3] ;
    input \motor_state_23__N_91[4] ;
    output \motor_state[4] ;
    input \motor_state_23__N_91[5] ;
    output \motor_state[5] ;
    input \motor_state_23__N_91[6] ;
    output \motor_state[6] ;
    input \motor_state_23__N_91[7] ;
    output \motor_state[7] ;
    input n28361;
    output n10;
    input \motor_state_23__N_91[9] ;
    output \motor_state[9] ;
    input \motor_state_23__N_91[10] ;
    output \motor_state[10] ;
    input \motor_state_23__N_91[11] ;
    output \motor_state[11] ;
    input \motor_state_23__N_91[12] ;
    output \motor_state[12] ;
    input \motor_state_23__N_91[13] ;
    output \motor_state[13] ;
    input \motor_state_23__N_91[14] ;
    output \motor_state[14] ;
    output n7_adj_13;
    input \motor_state_23__N_91[21] ;
    output \motor_state[21] ;
    input n28304;
    input \motor_state_23__N_91[17] ;
    output \motor_state[17] ;
    output n53323;
    input \motor_state_23__N_91[19] ;
    output \motor_state[19] ;
    input \motor_state_23__N_91[20] ;
    output \motor_state[20] ;
    output n25771;
    input \current[7] ;
    input \motor_state_23__N_91[22] ;
    output \motor_state[22] ;
    input \motor_state_23__N_91[23] ;
    output \motor_state[23] ;
    output n7_adj_14;
    input \motor_state_23__N_91[15] ;
    output \motor_state[15] ;
    input \motor_state_23__N_91[18] ;
    output \motor_state[18] ;
    input n58169;
    output n58405;
    output n58556;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    output n22760;
    input n52894;
    output n14;
    input n58366;
    input n66452;
    input n58711;
    output n25819;
    input n26235;
    output n26405;
    output n70252;
    input n58046;
    input n63899;
    input n63900;
    input n60683;
    output n69300;
    output n60931;
    input n63903;
    input n63902;
    output tx_o;
    output [8:0]r_Clock_Count;
    output tx_enable;
    input [31:0]baudrate;
    output n27845;
    output n58988;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_2;
    output [7:0]r_Clock_Count_adj_23;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    input n61478;
    input \r_SM_Main_2__N_3446[1] ;
    output \r_SM_Main[1] ;
    input n4939;
    output n25566;
    input n29596;
    input n29595;
    input n29591;
    input n29590;
    input n29559;
    input n29558;
    input n29557;
    output \r_Bit_Index[0] ;
    output n61043;
    input n30440;
    input n53943;
    input n30436;
    output \o_Rx_DV_N_3488[0] ;
    output n61750;
    output n61702;
    output n61734;
    output n61814;
    output n61782;
    output n61766;
    output n61798;
    output n61718;
    input n57927;
    output n27722;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n27996, n70121;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n51603, n66309, n58549, n26294, n7_c, n53195, n53787, 
        n58387, n58654, n58644, n6, n59809, n26364, n58357, n53734, 
        n51604, n26343, n58297, n25912, n6_adj_5263, n53818, n2, 
        n2_adj_5264, n53875, n14_c, n52883, n53723, n58445, n15_c, 
        n53258, n52799, n25145, Kp_23__N_872, Kp_23__N_869, n25947, 
        n26382, n58343, n52896, n53125, n58727, n8_c, n26261, 
        n58253, n52861, n52877, n58384, n58373, n58477, n6_adj_5265, 
        n53831, n58354, n58355, n53848, n58534, n6_adj_5266, n25743, 
        n1720, n10_c, n6_adj_5267, n53746, n58763, n23700, n6_adj_5268, 
        n52766, n58669, n58416, n10_adj_5269, n58381, n23704, n4, 
        n8_adj_5270, n3, n58028, n58484, n10_adj_5271, n52733, n6_adj_5272;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5273, n58501, n58025, n16, n1244, n58052, n58705, 
        n17_c, n17_adj_5274, n58120, n58186, n2_adj_5275, n58633, 
        n2_adj_5276, n26280, n2_adj_5277;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    
    wire n29670, n58259, n6_adj_5278, n53361, n7_adj_5279, n58474, 
        n52790, n58275, n26872, n25688, n2_adj_5280, n29609, n1516, 
        n58262, n58609, n12, n2_adj_5281, n58057, n58037, n26771, 
        n69296, n58741, n10_adj_5282;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    
    wire n29675, n26618, n10_adj_5283, n2_adj_5284, n58145, n14_adj_5285, 
        n25082, n58087, n58708, n12_adj_5286, n58021, n58523, n26402, 
        n58696, n26265, n1699, n1668, n58495, n2_adj_5287;
    wire [15:0]current_limit_c;   // verilog/TinyFPGA_B.v(251[22:35])
    
    wire n29678, n29679, n58699, n58071, n12_adj_5288, n29680, n58693, 
        n58604, n58242, n52569, n58481, n10_adj_5289, n2_adj_5290, 
        n2_adj_5291, n2_adj_5292, n1130, n1563, n26673, n58487, 
        n34_c, n2_adj_5293, n24, n58504, n38, n58111, n36, n32, 
        n40, n58031, n25737, n35, n58543, n10_adj_5294, n58717, 
        n14_adj_5295, n9, n26431, n53765, n6_adj_5296, n25680, n58232, 
        n58595, n10_adj_5297, n14_adj_5298, n53871, n2_adj_5299, n2_adj_5300, 
        n2_adj_5301, n58751, n36_adj_5302, n2_adj_5303, n34_adj_5304, 
        n26_c, n40_adj_5305, n53757, n38_adj_5306, n26667, n26340, 
        n52857, n42, n30, n58372, n41_c, n58769, n26794, n58739, 
        n58601, n26201, n58300, n63166, n62962;
    wire [7:0]\data_in_frame[0]_c ;   // verilog/coms.v(99[12:25])
    
    wire n25884, n58157, n58135, n10_adj_5308, n36_adj_5309, n14_adj_5310, 
        n25813, n26371;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    
    wire n42_adj_5311, n26663, n58138, n58552, n10_adj_5312, n52801, 
        n58375, n25806, Kp_23__N_767, n12_adj_5313, n58546, n53348, 
        n26427, n53891, n26875, n1655, n58636, n8_adj_5314, n26558, 
        n58333, n58197, n5, n58690, n58465, n58081, n23929, n12_adj_5317, 
        n58511, n52731, n58530, n6_adj_5318, n10_adj_5319, n26625, 
        n14_adj_5320, n58131, n58142;
    wire [7:0]\data_in_frame[3]_c ;   // verilog/coms.v(99[12:25])
    
    wire n26398, n25933, n58287, n10_adj_5321, n58468, n25915, n58507, 
        n58060, n26829;
    wire [7:0]\data_in_frame[8]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58589, n58217, n25862, n14_adj_5322, n58592, n58266, n15_adj_5323, 
        n58439, n26466, Kp_23__N_799, n58245, n58226, n58607, n58702, 
        n12_adj_5324, n58313, n58582, n25733, n26122;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire n70168, n66456, n70429, n58397, n53774, n58202, n26561, 
        n58461, n25924, n58540, n52831, n58369, n10_adj_5325, n53855, 
        n3_adj_5326, n2_adj_5327, n2_adj_5328, n2_adj_5329, n58105, 
        n2_adj_5330, n2_adj_5331, n2_adj_5332, n2_adj_5333, n58517, 
        Kp_23__N_878, n2_adj_5334;
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5335, n2_adj_5336, n27998, n51602, n66294, n2_adj_5337, 
        n14_adj_5338, n7_adj_5339;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n6_adj_5340, n2_adj_5341, n4_adj_5342, n2_adj_5343, n2_adj_5344, 
        n2_adj_5345, n2_adj_5346, n2_adj_5347, n2_adj_5348, n2_adj_5349, 
        Kp_23__N_974, n2_adj_5350, n2068, Kp_23__N_1748, n2_adj_5351, 
        n25755, n2_adj_5352, n2_adj_5353, n2_adj_5354;
    wire [23:0]n4764;
    
    wire n27736, n28000, n51601, n66286, n2_adj_5355, n2_adj_5356, 
        n58117, n28002, n51600, n66284, n2_adj_5357, n29812, n2_adj_5358, 
        n2_adj_5359, n29811, n2_adj_5360, n58256, n2_adj_5361, n2_adj_5362, 
        n58514, n2_adj_5363, n28004, n51599, n66282, n2_adj_5364, 
        n2_adj_5365, n63066, n63062, n2_adj_5366, n63064, n29809, 
        n58084, n63078, n2_adj_5367, n29808, n2_adj_5368, n63076, 
        n63082, n58223, n63088, n26337, n29807, n2_adj_5369, n29806, 
        n10_adj_5370, n2_adj_5371, n58166, n14_adj_5372, n63417, n60707, 
        n61042, n63431, n2_adj_5373, n2_adj_5374;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(246[14:26])
    
    wire n2_adj_5375, n3_adj_5376, n63549, n7_adj_5377, n28, n2_adj_5378, 
        n2_adj_5379, n2_adj_5380, n23933, n53607, n29_c, n58608;
    wire [7:0]\data_in_frame[7]_c ;   // verilog/coms.v(99[12:25])
    
    wire n63551, LED_N_3408, n52751, n8_adj_5381, n2_adj_5382, n58672, 
        n8_adj_5383;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n26414, n62972;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n58425, n62974, n58663, n8_adj_5384, n2_adj_5385, n2_adj_5386, 
        n2_adj_5387, n2_adj_5388, n2_adj_5389, n2_adj_5390, n2_adj_5391, 
        n2_adj_5392, n2_adj_5393, n2_adj_5394, n2_adj_5395, n2_adj_5396, 
        n2_adj_5397, n2_adj_5398, n2_adj_5399, n2_adj_5400, n5_adj_5401, 
        n58621, n62976, n52807, n58400, n62978, n58455, n61005, 
        n62980;
    wire [7:0]\data_in_frame[18]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58323, n6_adj_5402, n52776, n59838, n58269, n53750, n58612, 
        n10_adj_5403, n52879, n58403, n58458, n8_adj_5404, n26087, 
        n62982, n28006, n51598, n66281, n58330, n62984, n62986, 
        n52853, n58208, n60360;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n60585, n2_adj_5405, n2_adj_5406, n2_adj_5407, n2_adj_5408, 
        n2_adj_5409, n2_adj_5410, n2_adj_5411, n2_adj_5412, n58585, 
        n52410, n63156, n2_adj_5413, n2_adj_5414, n2_adj_5415, n2_adj_5416, 
        n2_adj_5417, n2_adj_5418, n2_adj_5419, n29805, n29804, n58681, 
        n63172, n63178, n58179, n60893, n63216, n28008, n51597, 
        n66256, n28010, n51596, n66255, n2_adj_5420, n62992, n58336, 
        n62994, n28012, n51595, n66254, n53861, n53829, n58211, 
        n60661, n58448, n63184, n62930, n2_adj_5421, n58745, n62998, 
        n25115, n60688, n63144, Kp_23__N_612, n28014, n51594, n66253, 
        n29803, \FRAME_MATCHER.i_31__N_2513 , n28016, n51593, n66252, 
        n28018, n51592, n66250, n2_adj_5422, n2_adj_5423, n2_adj_5424, 
        n44, n29802, n42_adj_5425, n43, n41_adj_5426, n57909, n50329, 
        n57901, n57908, n50328, n40_adj_5427, n57907, n50327, n28020, 
        n51591, n66246, n29801, n29800, n29799, n39, n50, n45, 
        n25529, n4452, \FRAME_MATCHER.i_31__N_2514 , n29798, n29797, 
        n101, n66307, n66304;
    wire [2:0]r_SM_Main_2__N_3545;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(32[16:25])
    
    wire n44525, n22192, n29796, n29795, n29794, n29793, n2_adj_5429, 
        n29792, n2_adj_5430, n57906, n50326, n28022, n51590, n66237, 
        n2_adj_5431, n57905, n50325, n2_adj_5432, n70210, n44533, 
        n57904, n50324;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    wire [2:0]n460;
    
    wire n28024, n51589, n66236, n25541, n2_adj_5433, n28026, n51588, 
        n66231, n2_adj_5434, n28028, n51587, n66224, n29791, n2_adj_5435, 
        n29790, n2_adj_5436, n2_adj_5437, n57903, n50323, n2_adj_5438, 
        n28045, n63777, n29789, n63778, n63776, n2_adj_5439, n2_adj_5440, 
        n29787, n2_adj_5441, n29786, n28030, n51586, n66221, n70222, 
        n70450, n29785, n29784, n61023, n29783, n2_adj_5442, n28032, 
        n51585, n66218, n29782, n2_adj_5443, n29781, n2_adj_5444, 
        n28034, n51584, n66217, n57902, tx_transmit_N_3416, n29780;
    wire [31:0]n133;
    
    wire n161, n29779, n2_adj_5445, n2_adj_5446, n2_adj_5447, n29778, 
        n2_adj_5448, n2_adj_5449, n29777, n2_adj_5450, n29776, n29775, 
        n70156, n70282, n68135, n29774, n70246, n29773, n29772, 
        n29771, n70150, n70288, n68139, n70240, n29770, n29769, 
        n29768, n1951, n60097, n20323, n22692, n63421, n27016, 
        n29767, n29766, n3303, \FRAME_MATCHER.i_31__N_2512 , n2060, 
        n29765, n29764, n29763, n29762, n29761, n29760, n29759, 
        n29758, n29757, n29756, n29755, n1954, n1957, n63325, 
        n29754, n29753, n60837, n57023, n29752, n29751, n29749, 
        n29748, n29747, n29746, n29745, n1955, n25514, n20328, 
        n29744, n29743, n25_c, n61073, n97, tx_active, n2049, 
        \FRAME_MATCHER.i_31__N_2507 , n29742, n771, \FRAME_MATCHER.i_31__N_2508 , 
        n2048, n25432, n29741, n5_adj_5452, n29740, n29739, n29738, 
        n27593, n60943, n25520, n27013;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n10_adj_5453;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n14_adj_5454, n25552;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n63320, n25590, n21, n20, n25526, n24_adj_5455, n25454, 
        n16_adj_5456, n17_adj_5457, n29737, n29736, n63539, n29735, 
        n9_adj_5458, n29734, n10_adj_5459, n18_c, n20_adj_5460, n15_adj_5461, 
        n16_adj_5462, n17_adj_5463, n57968, n6_adj_5464, n22691, n70526, 
        n42296, n57974, n2_adj_5465, n2_adj_5466, n2_adj_5467, n2_adj_5468, 
        n2_adj_5469, n29695, n2_adj_5470, n29694, n29693, n29692, 
        n29691, n29690, n29689, n2_adj_5471, n29597, n29688, n29687, 
        n29686, n29685, n29684, n29683, n29682, n29681, n2_adj_5472, 
        n2_adj_5473, n29956, n2_adj_5474, n2_adj_5475, n2_adj_5476, 
        n2_adj_5477, Kp_23__N_748, n24_adj_5478, n29649, n29648, n29647, 
        n2_adj_5479, n2_adj_5480, n29638, n29629, n57285, n2_adj_5482, 
        n2_adj_5483, n2_adj_5484, n2_adj_5485, n63794, n63795, n63801, 
        n63800, n29618, n29616, n29614, n29613, n29612, n2_adj_5487, 
        n63653, n63654, n2_adj_5488, n2_adj_5489, n2_adj_5490, n2_adj_5491, 
        n2_adj_5492, n2_adj_5493, n2_adj_5494, n2_adj_5495, n2_adj_5496, 
        n2_adj_5497, n2_adj_5498, n2_adj_5499, n63729, n2_adj_5500, 
        n2_adj_5501, n2_adj_5503, n2_adj_5504, n63728, n2_adj_5505, 
        n2_adj_5506, n2_adj_5508, n2_adj_5509, n2_adj_5510, n2_adj_5511, 
        n2_adj_5512, n2_adj_5513, n2_adj_5514, n2_adj_5515, n2_adj_5516, 
        n2_adj_5517, n2_adj_5518, n2_adj_5519, n63842, n2_adj_5520, 
        n2_adj_5521, n2_adj_5522, n63843, n63657, n63656, n63833, 
        n63834, n63771, n27972, n2_adj_5523, n2_adj_5524, n63770, 
        n2_adj_5525, n27974, n27976, n58909, n59553, n29148, n66400, 
        n63768, n27978, n27980, n27982, n27984, n27986, n27988, 
        n27990, n27992, n27994, n2_adj_5526, n42499, n30068, n63769, 
        n63767, n29550, n70198, n70480, n14_adj_5527, n63824, n70258, 
        n29547, n63825, n29535, n63810, n63809, n29532, n2_adj_5528, 
        n29529, n2_adj_5529, n63812, n63813, n29526, n29523, n63819, 
        n63818, n63785, n57109, n63786, n57129, n14_adj_5531;
    wire [7:0]\data_in_frame[19]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30408, n63873, n36387, n30353, n30352, n30351, n30350, 
        n30349, n30348, n30347, n30346, n30345, n30344, n30343, 
        n30342, n30341, n30340, n30339, n63872, n30338, n30337, 
        n30336, n30335, n30334, n30333, n30332, n30331, n30330, 
        n30329, n30328, n30327, n30326, n30325, n30324, n30323, 
        n30322, n17_adj_5532, n57325, n30315, n29416, n29420, n25_adj_5533, 
        n29427, n29430, n9_adj_5534, n29436, n57449, n29445, n29448, 
        n29451, n57319, n29911, n29915, n57379, n30295, n30290, 
        n29460, n29463, n29918, n29921, n29925, n29928, n29931, 
        n30275, n29934, n29937;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    
    wire n29941, n29944, n29947, n29466, n29469, n29950, n29953, 
        n29957, n29960, n29963;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    
    wire n29967, n29970, n29973, n29977, n29980, n29983, n29987, 
        n29990;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    
    wire n29993, n57277, n30000, n57339, n30007, n30010, n30013, 
        n30017, n70270, n66234, n30246, n30020;
    wire [7:0]\data_in_frame[12]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30023, n30027, n30030, n30033, n30037, n30040, n30043;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    
    wire n66436, n8_adj_5535, n30047, n30050, n30053, n30056, n30059, 
        n30062, n30065, n30069;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    
    wire n57355, n30075, n30079, n30082, n30085, n30089, n30092, 
        n30095, n30099, n30102, n30105, n30109, n30112, n30115, 
        n30119, n8_adj_5536, n57239;
    wire [7:0]\data_in_frame[17]_c ;   // verilog/coms.v(99[12:25])
    
    wire n57241, n29475, n57125, n57127, n57269, n30176, n63756, 
        n2_adj_5537, n63757, n58889, n29544, n63755, n2_adj_5538, 
        n57993, n57341, n2_adj_5539, n57303, n2_adj_5540, n2_adj_5541, 
        n70315, n70294, n66457, n28039, n63750, n63751, n63749, 
        n63732, n70300, n66439, n29419, n63650, n63651, n63897, 
        n63896, n63836, n63837, n63747, n63746, n63731, n70309, 
        \FRAME_MATCHER.i_31__N_2511 , n58004, n27276, n63735, n3472, 
        n1, n63734, n28037, n63738, n63739, n63737, n40523, n70216, 
        n70462, n14_adj_5542, n63908;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n57923, n57924, n10_adj_5543, n52835, n57925, n63909, n70306, 
        n66247, n58346, n53785, n58639, n63888, n57911, n63887, 
        n66502, n12_adj_5544, n10_adj_5545, n11, n9_adj_5546, n58065, 
        n60617, n57926, n22, n27_adj_5547, n26_adj_5548, n29_adj_5549, 
        n31, n63337, n10_adj_5550, n4_adj_5551;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n57912, n57913, n3_adj_5552, n57914, n3_adj_5553, n57915, 
        n3_adj_5554, n57916, n3_adj_5555, n57917, n3_adj_5556, n57918, 
        n3_adj_5557, n57919, n3_adj_5558, n57920, n3_adj_5559, n57921, 
        n3_adj_5560, n57922, n3_adj_5561, n3_adj_5562, n3_adj_5563, 
        n3_adj_5564, n3_adj_5565, n1_adj_5566, n1_adj_5567, n1_adj_5568, 
        n1_adj_5569, n1_adj_5570, n1_adj_5571, n86, n1_adj_5572, n28829, 
        n5_adj_5573, n28828, n26923, n28827, n1_adj_5576, n2_adj_5577, 
        n2_adj_5578, n2_adj_5579, n70303, n70297, n58229, n52743, 
        n58575, n53902, n8_adj_5580, n58731, n66310, n66289, n66312, 
        n66313, n51614, n66361, n66323, n58562, n58183, n28314, 
        n51613, n66356, n51612, n66355, n66324, n51611, n66354, 
        n51610, n66350, n8_adj_5581, n51609, n66347, n51608, n51607, 
        n51606, n51605, n58128, n52885, n25130, n26379, n25218, 
        n58093, n58090, n58598, n53066, n53743, n10_adj_5582, n25716, 
        n58068, n58154, n26463, n26274, n58657, n26493, n58310, 
        n58316, n4_adj_5583, n53833, n58015, n6_adj_5584, n53853, 
        n6_adj_5585, n28322, n25974, n20_adj_5586, n63190, n53763, 
        n8_adj_5587, n12_adj_5588, n6_adj_5589, n57986, n57983, n58012, 
        n26042, n58666, n26853, n6_adj_5590, n58419, n53720, n53921, 
        n53137, n25141, n36_adj_5592, n25996, n53737, n58272, n53706, 
        n58675, n26330, n63108, n53776, n52407, n60610, n66360, 
        n7_adj_5594, n7_adj_5595, n7_adj_5596, n6_adj_5597, n6_adj_5598, 
        n58392, n53933, n53824, n7_adj_5599, n70291, n63258, n57571, 
        n6_adj_5602, n12_adj_5603, n59012, n53963, n58678, n58435, 
        n63010, n63012, n58220, n25908, n58490, n63020, Kp_23__N_1067, 
        n58648, n63024, n52778, n60724, n58624, n63030, n63032, 
        n52737, n63038, n58432, n63044, n58096, n23886, n63132, 
        n58339, n63136, n63118, n63124, n58391, n14_adj_5606, n58714, 
        n15_adj_5607, n63206, n58378, n53795, n58627, n63224, n58451, 
        n63146, n62968, n63230, n6_adj_5608, n58176, n52723, n58034, 
        n16_adj_5609, n53770, n17_adj_5610, n58615, n53728, n58114, 
        n58429, n6_adj_5611, n25103, n59945, n58148, n60258, n14_adj_5612, 
        n15_adj_5613, n58742, n58163, n10_adj_5614, n59815, n6_adj_5616, 
        n4_adj_5617, n58526, n58160, Kp_23__N_1256, n58284, n58630, 
        n63250, n63252, n63254, n63262, n63268, n58413, n63274, 
        n58250, n16_adj_5618, n22_adj_5619, n24_adj_5620, n58733, 
        n58422, n25898, n62948, n62954, n58660, n63284, n58290, 
        n58173, n58078, n12_adj_5621, n28_adj_5622, n31_adj_5623, 
        n30_adj_5624, n34_adj_5625, n29_adj_5626, n58757, LED_N_3407, 
        n3_adj_5627, n70285, n70279, n5_adj_5628, n58214, n53918, 
        n26249, n58723, n58760, n58351, n6_adj_5630, n70501, n60186, 
        n26865, n60779, n58408, n59988, n58361, n58360, n58565, 
        n12_adj_5631, n63832, n58720, n70126, n70495, n70267, n58687, 
        n70228, n52786, n70261, n70132, n70483, n14_adj_5632, n16_adj_5633, 
        n58205, n22_adj_5634, n70264, n60912, n20_adj_5635, n24_adj_5636, 
        n70255, n10_adj_5637, n58293, n6_adj_5638, n66494, n26704, 
        n70249, n70477, n58442, n30_adj_5639, n18_adj_5640, n24_adj_5641, 
        n61386, n85, n53949, n22_adj_5642, n26_adj_5643, n60672, 
        n34_adj_5644, n32_adj_5645, n33, n58281, n31_adj_5646, n70180, 
        n70243, n70174, n70204, n70237, n70231, n70234, n58108, 
        n70225, n70219, n53789, n70213, n63851, n63852, n70207, 
        n63849, n63848, n70138, n70471, n70201, n70144, n70465, 
        n70195, n70459, n12_adj_5647, n52546, n70177, n70171, n60828, 
        n70162, n70453, n70165, n70159, n70153, n42_adj_5648, n40_adj_5649, 
        n41_adj_5650, n70147, n70447, n39_adj_5651, n38_adj_5652, 
        n37, n48, n43_adj_5653, n58363, n70141, n70135, n70129, 
        n70123, n14_adj_5654, n13, n8_adj_5655, n15_adj_5656, n58579, 
        n13_adj_5657;
    
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_22_lut  (.I0(n66309), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n51603), .O(n27996)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n29606));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29891));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[4] [5]), .I1(n58549), .I2(GND_net), 
            .I3(GND_net), .O(n26294));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[22] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_c));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n7_c), .I1(n53195), .I2(n53787), .I3(n58387), 
            .O(n58654));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1062 (.I0(n58644), .I1(\data_out_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i2_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n59809), .I1(n26364), .I2(n6), .I3(n58357), 
            .O(n53734));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29888));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_22  (.CI(n51603), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n51604));
    SB_LUT4 i3_4_lut (.I0(n26343), .I1(\data_in_frame[6] [6]), .I2(\data_in_frame[4] [6]), 
            .I3(\data_in_frame[7] [0]), .O(n58297));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25912));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1064 (.I0(n53734), .I1(n58654), .I2(\data_out_frame[21] [7]), 
            .I3(n6_adj_5263), .O(n53818));
    defparam i4_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2), .S(n57860));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5264), .S(n57859));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut (.I0(n53734), .I1(n53875), .I2(\data_out_frame[22] [1]), 
            .I3(GND_net), .O(n14_c));
    defparam i5_3_lut.LUT_INIT = 16'h6969;
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29885));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut (.I0(n58644), .I1(n52883), .I2(n53723), .I3(n58445), 
            .O(n15_c));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_c), .I1(n53258), .I2(n14_c), .I3(n52799), 
            .O(n25145));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1065 (.I0(n25912), .I1(Kp_23__N_872), .I2(Kp_23__N_869), 
            .I3(\data_in_frame[8] [4]), .O(n25947));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[25] [7]), 
            .I2(n26382), .I3(GND_net), .O(n58343));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1066 (.I0(\data_out_frame[19] [5]), .I1(n52896), 
            .I2(n53125), .I3(GND_net), .O(n26364));
    defparam i2_3_lut_adj_1066.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_out_frame[21] [7]), .I1(\data_out_frame[21] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58727));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[17] [5]), .I3(GND_net), .O(n8_c));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[18] [0]), .I1(n26261), .I2(n8_c), 
            .I3(n58253), .O(n58651));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1068 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n52861), .I3(GND_net), .O(n52877));
    defparam i2_3_lut_adj_1068.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58384));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1070 (.I0(\data_out_frame[18] [2]), .I1(n58373), 
            .I2(n58477), .I3(n6_adj_5265), .O(n53831));
    defparam i4_4_lut_adj_1070.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58354));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(n53258), .I1(n58354), .I2(GND_net), 
            .I3(GND_net), .O(n58355));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(n53848), .I1(n58534), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5266));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1074 (.I0(n53831), .I1(n25743), .I2(n58384), 
            .I3(n6_adj_5266), .O(n53723));
    defparam i4_4_lut_adj_1074.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1075 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [4]), .I3(n1720), .O(n10_c));
    defparam i4_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1076 (.I0(n58727), .I1(n26364), .I2(\data_out_frame[23] [7]), 
            .I3(n52883), .O(n6_adj_5267));
    defparam i1_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1077 (.I0(n53746), .I1(n58570), .I2(n58763), 
            .I3(n6_adj_5267), .O(n23700));
    defparam i4_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_out_frame[20] [3]), .I1(n53723), 
            .I2(GND_net), .I3(GND_net), .O(n53787));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(n25705), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5268));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1080 (.I0(\data_out_frame[17] [4]), .I1(n52766), 
            .I2(\data_out_frame[15] [3]), .I3(n6_adj_5268), .O(n53125));
    defparam i4_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_out_frame[17] [6]), .I1(n25705), 
            .I2(GND_net), .I3(GND_net), .O(n58669));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_out_frame[19] [6]), .I1(n53125), 
            .I2(GND_net), .I3(GND_net), .O(n58416));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1083 (.I0(n58416), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[22] [2]), .I3(n58669), .O(n10_adj_5269));
    defparam i4_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(n25145), .I1(n53818), .I2(GND_net), 
            .I3(GND_net), .O(n58381));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1085 (.I0(n53787), .I1(n23700), .I2(n23704), 
            .I3(n4), .O(n8_adj_5270));
    defparam i3_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_209_i3_4_lut (.I0(n58343), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5270), .I3(n58354), .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i4_4_lut_adj_1086 (.I0(n58028), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[12] [7]), .I3(n58484), .O(n10_adj_5271));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(n52733), .I1(n26261), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5272));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1088 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(n6_adj_5272), .O(n52896));
    defparam i4_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5273));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1089 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[10] [3]), 
            .I2(n58501), .I3(n58025), .O(n16));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n1244), .I1(n58052), .I2(n58705), .I3(n17_c), 
            .O(n17_adj_5274));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17_adj_5274), .I1(\data_out_frame[5] [5]), .I2(n16), 
            .I3(\data_out_frame[12] [6]), .O(n52733));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1090 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(n58120), .I3(n52733), .O(n58186));
    defparam i3_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5275));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58633));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5276));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26280));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5277));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i21273_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n22773), .I3(GND_net), .O(n29670));
    defparam i21273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1093 (.I0(\data_out_frame[21] [4]), .I1(\data_out_frame[19] [3]), 
            .I2(n58259), .I3(n6_adj_5278), .O(n53361));
    defparam i4_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1094 (.I0(\data_out_frame[21] [3]), .I1(n58186), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5279));
    defparam i2_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1095 (.I0(n7_adj_5279), .I1(n26280), .I2(n53848), 
            .I3(n58474), .O(n52790));
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1096 (.I0(\data_out_frame[14] [4]), .I1(n58275), 
            .I2(\data_out_frame[17] [0]), .I3(GND_net), .O(n26872));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1096.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25688));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5280));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n29609));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut (.I0(n1516), .I1(n58262), .I2(n25688), .I3(n58609), 
            .O(n12));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5281));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1098 (.I0(n58057), .I1(n12), .I2(\data_out_frame[14] [6]), 
            .I3(n58037), .O(n26771));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1099 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [7]), 
            .I2(n69296), .I3(n58741), .O(n10_adj_5282));
    defparam i4_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i21380_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n22773), .I3(GND_net), .O(n29675));
    defparam i21380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1100 (.I0(n26618), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5283));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_adj_1100.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5284));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1101 (.I0(n58145), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[9] [1]), .O(n14_adj_5285));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1102 (.I0(\data_out_frame[9] [3]), .I1(n14_adj_5285), 
            .I2(n10_adj_5283), .I3(\data_out_frame[11] [3]), .O(n25082));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1103 (.I0(\data_out_frame[5] [1]), .I1(n58087), 
            .I2(n58708), .I3(\data_out_frame[9] [2]), .O(n12_adj_5286));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1104 (.I0(n58021), .I1(n12_adj_5286), .I2(n58523), 
            .I3(\data_out_frame[11] [4]), .O(n26402));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1105 (.I0(\data_out_frame[11] [0]), .I1(n58052), 
            .I2(GND_net), .I3(GND_net), .O(n58696));
    defparam i1_2_lut_adj_1105.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(n25705), .I1(n26265), .I2(GND_net), 
            .I3(GND_net), .O(n1720));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58705));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(88[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58495));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5287));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23552_3_lut (.I0(current_limit_c[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n22773), .I3(GND_net), .O(n29678));
    defparam i23552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23553_3_lut (.I0(current_limit_c[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n22773), .I3(GND_net), .O(n29679));
    defparam i23553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1109 (.I0(\data_out_frame[6] [0]), .I1(n58699), 
            .I2(n58071), .I3(n58099), .O(n12_adj_5288));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i23557_3_lut (.I0(current_limit_c[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n22773), .I3(GND_net), .O(n29680));
    defparam i23557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1110 (.I0(\data_out_frame[10] [4]), .I1(n12_adj_5288), 
            .I2(\data_out_frame[13] [0]), .I3(n58495), .O(n52766));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1111 (.I0(\data_out_frame[13] [1]), .I1(n26618), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n58484));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1111.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58087));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1113 (.I0(n58087), .I1(n58693), .I2(n58604), 
            .I3(n58242), .O(n52569));
    defparam i3_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1114 (.I0(n58481), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[14] [0]), .I3(n58693), .O(n10_adj_5289));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5290));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5291));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5292));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58481));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58037));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58501));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58604));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1119 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26618));
    defparam i2_3_lut_adj_1119.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(\data_out_frame[10] [0]), .I1(n1563), 
            .I2(\data_out_frame[11] [4]), .I3(n26673), .O(n58487));
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n58604), .I1(\data_out_frame[7] [4]), .I2(n58057), 
            .I3(\data_out_frame[6] [7]), .O(n34_c));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5293));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i17_4_lut (.I0(\data_out_frame[7] [0]), .I1(n34_c), .I2(n24), 
            .I3(n58504), .O(n38));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n1130), .I1(\data_out_frame[6] [6]), .I2(n58111), 
            .I3(\data_out_frame[6] [4]), .O(n36));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[6] [1]), .I1(n38), .I2(n32), 
            .I3(\data_out_frame[4] [4]), .O(n40));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(n25676), .I1(n58031), .I2(n25737), .I3(\data_out_frame[4] [7]), 
            .O(n35));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29881));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1121 (.I0(n58543), .I1(n35), .I2(n40), .I3(n36), 
            .O(n10_adj_5294));
    defparam i2_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1122 (.I0(n58717), .I1(\data_out_frame[9] [6]), 
            .I2(n58481), .I3(\data_out_frame[9] [7]), .O(n14_adj_5295));
    defparam i6_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29872));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1123 (.I0(n9), .I1(n26431), .I2(n14_adj_5295), 
            .I3(n10_adj_5294), .O(n53765));
    defparam i1_4_lut_adj_1123.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n58052));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(n58052), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5296));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1126 (.I0(\data_out_frame[11] [0]), .I1(n25680), 
            .I2(\data_out_frame[6] [1]), .I3(n6_adj_5296), .O(n58028));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1127 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n58232));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58595));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1129 (.I0(n53765), .I1(n58487), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5297));   // verilog/coms.v(88[17:63])
    defparam i2_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29869));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1130 (.I0(n58595), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[11] [5]), .I3(n58232), .O(n14_adj_5298));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29866));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1131 (.I0(n58028), .I1(n14_adj_5298), .I2(n10_adj_5297), 
            .I3(\data_out_frame[11] [1]), .O(n53871));   // verilog/coms.v(88[17:63])
    defparam i7_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29863));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25737));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29860));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5299));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29857));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29854));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29851));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14_4_lut_adj_1133 (.I0(n25737), .I1(n52861), .I2(n53871), 
            .I3(n58751), .O(n36_adj_5302));
    defparam i14_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5303));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29848));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n29621));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29844));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29838));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[8] [6]), .I1(n1699), .I2(n58705), 
            .I3(n58232), .O(n34_adj_5304));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n52766), .I1(n36_adj_5302), .I2(n26_c), .I3(\data_out_frame[14] [3]), 
            .O(n40_adj_5305));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[8] [5]), .I1(n1720), .I2(n53757), 
            .I3(\data_out_frame[14] [1]), .O(n38_adj_5306));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1134 (.I0(n26667), .I1(n58297), .I2(n26340), 
            .I3(GND_net), .O(n26306));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[14] [6]), .I1(n40_adj_5305), 
            .I2(n34_adj_5304), .I3(n52857), .O(n42));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1135 (.I0(n58696), .I1(n38_adj_5306), .I2(n30), 
            .I3(n58372), .O(n41_c));
    defparam i19_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1136 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [3]), 
            .I2(n41_c), .I3(n42), .O(n58769));
    defparam i2_4_lut_adj_1136.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1137 (.I0(\data_out_frame[15] [0]), .I1(n58751), 
            .I2(GND_net), .I3(GND_net), .O(n58120));
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25743));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58477));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_out_frame[13] [5]), .I1(n25082), 
            .I2(GND_net), .I3(GND_net), .O(n26794));
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1141 (.I0(n26794), .I1(n58477), .I2(n25743), 
            .I3(GND_net), .O(n58739));
    defparam i2_3_lut_adj_1141.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_c));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29818));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1143 (.I0(\data_out_frame[5] [4]), .I1(n25666), 
            .I2(n17_c), .I3(n34), .O(n58601));   // verilog/coms.v(100[12:26])
    defparam i2_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1144 (.I0(n26201), .I1(n58300), .I2(\data_in_frame[5] [2]), 
            .I3(\data_in_frame[7] [4]), .O(n63166));
    defparam i1_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58242));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1146 (.I0(n63166), .I1(n62962), .I2(\data_in_frame[0]_c [6]), 
            .I3(n25884), .O(n58157));
    defparam i1_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58111));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58135));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1149 (.I0(n58242), .I1(n58601), .I2(\data_out_frame[7] [0]), 
            .I3(n58031), .O(n58708));
    defparam i3_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1150 (.I0(n58543), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5308));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1151 (.I0(n58708), .I1(\data_out_frame[6] [7]), 
            .I2(n58135), .I3(n36_adj_5309), .O(n14_adj_5310));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1152 (.I0(n25813), .I1(\data_in_frame[4] [4]), 
            .I2(n26371), .I3(GND_net), .O(n26340));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1153 (.I0(\data_out_frame[13] [3]), .I1(n14_adj_5310), 
            .I2(n10_adj_5308), .I3(\data_out_frame[8] [7]), .O(n26265));   // verilog/coms.v(88[17:28])
    defparam i7_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58262));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1155 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[8] [0]), .O(n58504));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[2] [7]), .I1(n25884), .I2(\data_in_frame[0][5] ), 
            .I3(GND_net), .O(n26201));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(\data_out_frame[4] [0]), .I1(n58504), 
            .I2(n58262), .I3(n42_adj_5311), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26673));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1158 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[7] [1]), .O(n58145));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1159 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n58071));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58717));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[4] [7]), .I1(n26663), 
            .I2(GND_net), .I3(GND_net), .O(n58138));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(\data_out_frame[8] [6]), .I1(n58071), 
            .I2(GND_net), .I3(GND_net), .O(n36_adj_5309));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1163 (.I0(n58552), .I1(n36_adj_5309), .I2(\data_out_frame[13] [4]), 
            .I3(n58717), .O(n10_adj_5312));
    defparam i4_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1164 (.I0(n58145), .I1(n10_adj_5312), .I2(n26673), 
            .I3(GND_net), .O(n52801));
    defparam i5_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_out_frame[15] [5]), .I1(n26265), 
            .I2(GND_net), .I3(GND_net), .O(n58375));
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1166 (.I0(\data_in_frame[7] [3]), .I1(n58138), 
            .I2(n25806), .I3(Kp_23__N_767), .O(n12_adj_5313));   // verilog/coms.v(74[16:69])
    defparam i5_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1167 (.I0(n26201), .I1(n12_adj_5313), .I2(\data_in_frame[0]_c [7]), 
            .I3(n58546), .O(n53348));   // verilog/coms.v(74[16:69])
    defparam i6_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26427));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26111));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_out_frame[14] [3]), .I1(n53891), 
            .I2(GND_net), .I3(GND_net), .O(n26875));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h9999;
    SB_LUT4 i3_3_lut_adj_1171 (.I0(n53848), .I1(n1655), .I2(n58636), .I3(GND_net), 
            .O(n8_adj_5314));
    defparam i3_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i53570_4_lut (.I0(n26558), .I1(n26875), .I2(n8_adj_5314), 
            .I3(n58333), .O(n69296));
    defparam i53570_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1288_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(88[17:28])
    defparam i1288_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1172 (.I0(n26558), .I1(n53848), .I2(\data_out_frame[16] [7]), 
            .I3(GND_net), .O(n58197));
    defparam i2_3_lut_adj_1172.LUT_INIT = 16'h6969;
    SB_LUT4 i26777_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_7), .O(n5));
    defparam i26777_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(n58690), .I1(n58739), .I2(GND_net), 
            .I3(GND_net), .O(n58741));
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58465));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58081));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(n26663), .I1(n58157), .I2(GND_net), 
            .I3(GND_net), .O(n23929));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1177 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[7] [5]), .I3(n26201), .O(n12_adj_5317));   // verilog/coms.v(73[16:69])
    defparam i5_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1178 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_5317), 
            .I2(n58511), .I3(\data_in_frame[5] [3]), .O(n52731));   // verilog/coms.v(73[16:69])
    defparam i6_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[2][1] ), .I1(n58530), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5318));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1180 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5319));   // verilog/coms.v(77[16:27])
    defparam i2_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1181 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(n26625), .O(n14_adj_5320));   // verilog/coms.v(77[16:27])
    defparam i6_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1182 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[0][0] ), 
            .I2(n58131), .I3(n6_adj_5318), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1183 (.I0(\data_out_frame[10] [0]), .I1(n14_adj_5320), 
            .I2(n10_adj_5319), .I3(\data_out_frame[7] [6]), .O(n58142));   // verilog/coms.v(77[16:27])
    defparam i7_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_in_frame[3]_c [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26398));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_in_frame[8] [2]), .I1(n25933), 
            .I2(GND_net), .I3(GND_net), .O(n58287));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1186 (.I0(\data_out_frame[5] [3]), .I1(n42_adj_5311), 
            .I2(\data_out_frame[12] [3]), .I3(n58081), .O(n10_adj_5321));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58468));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1188 (.I0(n25915), .I1(n58507), .I2(n58060), 
            .I3(n26398), .O(n26829));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25666));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[8]_c [5]), .I1(Kp_23__N_872), 
            .I2(GND_net), .I3(GND_net), .O(n58589));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1191 (.I0(n58217), .I1(n58589), .I2(\data_in_frame[6] [3]), 
            .I3(GND_net), .O(n25862));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1191.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1192 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[2][5] ), .I3(GND_net), .O(n14_adj_5322));
    defparam i5_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1193 (.I0(n58592), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[3][0] ), .I3(n58266), .O(n15_adj_5323));
    defparam i6_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26625));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58552));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1196 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n58439));
    defparam i2_3_lut_adj_1196.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1197 (.I0(n15_adj_5323), .I1(\data_in_frame[0] [2]), 
            .I2(n14_adj_5322), .I3(\data_in_frame[4] [6]), .O(n26466));
    defparam i8_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1198 (.I0(Kp_23__N_799), .I1(n58245), .I2(n58226), 
            .I3(\data_in_frame[6] [0]), .O(n58607));
    defparam i1_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(74[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1199 (.I0(n1563), .I1(n58702), .I2(n58021), .I3(n58439), 
            .O(n12_adj_5324));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1200 (.I0(\data_out_frame[12] [0]), .I1(n12_adj_5324), 
            .I2(\data_out_frame[14] [2]), .I3(n58498), .O(n58313));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_out_frame[14] [4]), .I1(n58313), 
            .I2(GND_net), .I3(GND_net), .O(n52857));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1202 (.I0(n58741), .I1(n58197), .I2(n2076), .I3(n69296), 
            .O(n58582));   // verilog/coms.v(88[17:28])
    defparam i2_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1203 (.I0(n53848), .I1(n58474), .I2(n25733), 
            .I3(GND_net), .O(n26122));
    defparam i2_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54667 (.I0(byte_transmit_counter[3]), 
            .I1(n70168), .I2(n66456), .I3(byte_transmit_counter[4]), .O(n70429));
    defparam byte_transmit_counter_3__bdd_4_lut_54667.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(n25915), .I1(n58397), .I2(GND_net), 
            .I3(GND_net), .O(n53774));
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n58131));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1206 (.I0(n58202), .I1(\data_out_frame[19] [0]), 
            .I2(n26122), .I3(n58582), .O(n26561));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(n52790), .I1(n53361), .I2(GND_net), 
            .I3(GND_net), .O(n58461));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1208 (.I0(n25924), .I1(n58131), .I2(\data_in_frame[6] [1]), 
            .I3(GND_net), .O(n58540));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1208.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_out_frame[21] [2]), .I1(n26561), 
            .I2(GND_net), .I3(GND_net), .O(n52831));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1210 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[23] [4]), .I3(n52883), .O(n58369));
    defparam i3_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n29641));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1211 (.I0(n58369), .I1(n52831), .I2(\data_out_frame[25] [6]), 
            .I3(n58461), .O(n10_adj_5325));
    defparam i4_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_208_i3_4_lut (.I0(n53855), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5325), .I3(\data_out_frame[25] [7]), .O(n3_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_780_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n29657));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1212 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(n58530), .I3(n58105), .O(n58217));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1213 (.I0(n58075), .I1(n58517), .I2(n26343), 
            .I3(GND_net), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1]_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58060));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1215 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25924));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1215.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_21_lut  (.I0(n66294), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n51602), .O(n27998)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29813));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5337), .S(n57858));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n70429_bdd_4_lut (.I0(n70429), .I1(n14_adj_5338), .I2(n7_adj_5339), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n70429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1216 (.I0(n25924), .I1(\data_in_frame[1][7] ), 
            .I2(n58060), .I3(n6_adj_5340), .O(Kp_23__N_869));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1217 (.I0(n25933), .I1(Kp_23__N_869), .I2(\data_in_frame[6] [2]), 
            .I3(\data_in_frame[8][3] ), .O(n4_adj_5342));   // verilog/coms.v(239[9:81])
    defparam i3_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5345), .S(n57857));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1218 (.I0(Kp_23__N_878), .I1(n58217), .I2(\data_in_frame[6] [5]), 
            .I3(GND_net), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1218.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_21  (.CI(n51602), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n51603));
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2068), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 select_780_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1219 (.I0(\data_in_frame[5] [5]), .I1(n58300), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n25755));
    defparam i1_3_lut_adj_1219.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27736), 
            .D(n4764[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_20_lut  (.I0(n66286), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n51601), .O(n28000)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_20  (.CI(n51601), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n51602));
    SB_LUT4 i1_3_lut_adj_1220 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[3]_c [4]), .I3(GND_net), .O(n25915));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(n25813), .I1(n26343), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_799));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(n25915), .I1(n25755), .I2(GND_net), 
            .I3(GND_net), .O(n58117));
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_19_lut  (.I0(n66284), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n51600), .O(n28002)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_780_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[3][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n62962));
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29812), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[2][0] ), .I1(n26371), 
            .I2(GND_net), .I3(GND_net), .O(n58105));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29811), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[3][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n58256));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_19  (.CI(n51600), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n51601));
    SB_LUT4 select_780_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1226 (.I0(\data_in_frame[3]_c [6]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58514));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1227 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58507));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[5] [2]), .I3(GND_net), .O(n58546));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1229 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58517));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1229.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n29698));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_18_lut  (.I0(n66282), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n51599), .O(n28004)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58592));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h6666;
    SB_LUT4 select_780_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1231 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1]_c [4]), 
            .I2(\data_in_frame[2][1] ), .I3(\data_in_frame[2] [7]), .O(n63066));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1232 (.I0(\data_in_frame[3][7] ), .I1(\data_in_frame[3][5] ), 
            .I2(\data_in_frame[2][3] ), .I3(\data_in_frame[4] [0]), .O(n63062));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1233 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[4] [5]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[4] [7]), .O(n63064));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29809), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1234 (.I0(n58084), .I1(n58592), .I2(n58517), 
            .I3(n63066), .O(n63078));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29808), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5368), .S(n57900));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1235 (.I0(n58546), .I1(n63064), .I2(n63062), 
            .I3(GND_net), .O(n63076));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1236 (.I0(n63076), .I1(n63078), .I2(n58507), 
            .I3(n58514), .O(n63082));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1237 (.I0(n63082), .I1(n58223), .I2(n58105), 
            .I3(n58530), .O(n63088));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1238 (.I0(n26337), .I1(n62962), .I2(n58117), 
            .I3(n63088), .O(n58245));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29807), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29806), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1239 (.I0(n58226), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5370));
    defparam i2_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5371), .S(n57856));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1240 (.I0(n58245), .I1(n25813), .I2(n58166), 
            .I3(\data_in_frame[8]_c [1]), .O(n14_adj_5372));
    defparam i6_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i47702_3_lut (.I0(Kp_23__N_974), .I1(n4_adj_5342), .I2(\data_in_frame[8][6] ), 
            .I3(GND_net), .O(n63417));
    defparam i47702_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i7_4_lut_adj_1241 (.I0(\data_in_frame[3]_c [6]), .I1(n14_adj_5372), 
            .I2(n10_adj_5370), .I3(n26343), .O(n60707));
    defparam i7_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i47715_2_lut (.I0(n61042), .I1(n26466), .I2(GND_net), .I3(GND_net), 
            .O(n63431));
    defparam i47715_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1242 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [6]), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1242.LUT_INIT = 16'ha088;
    SB_LUT4 select_780_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1243 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [4]), 
            .I2(control_mode_c[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1243.LUT_INIT = 16'ha088;
    SB_LUT4 i47832_4_lut (.I0(n3_adj_5376), .I1(n60707), .I2(n25862), 
            .I3(n63417), .O(n63549));
    defparam i47832_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n52731), .I1(n23929), .I2(n7_adj_5377), .I3(n53348), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_4_lut_adj_1244 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [3]), 
            .I2(control_mode_c[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1244.LUT_INIT = 16'ha088;
    SB_LUT4 select_780_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1245 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [1]), 
            .I2(\control_mode[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1245.LUT_INIT = 16'ha088;
    SB_LUT4 i12_4_lut_adj_1246 (.I0(n23933), .I1(n26306), .I2(n53607), 
            .I3(n25947), .O(n29_c));
    defparam i12_4_lut_adj_1246.LUT_INIT = 16'h0020;
    SB_LUT4 i47834_4_lut (.I0(n58608), .I1(n63431), .I2(n26294), .I3(\data_in_frame[7]_c [7]), 
            .O(n63551));
    defparam i47834_4_lut.LUT_INIT = 16'hfefd;
    SB_LUT4 i16_4_lut_adj_1247 (.I0(n63551), .I1(n29_c), .I2(n28), .I3(n63549), 
            .O(LED_N_3408));
    defparam i16_4_lut_adj_1247.LUT_INIT = 16'h0040;
    SB_LUT4 i3_3_lut_adj_1248 (.I0(\data_in_frame[20][4] ), .I1(\data_in_frame[20] [5]), 
            .I2(n52751), .I3(GND_net), .O(n8_adj_5381));
    defparam i3_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_adj_1249 (.I0(\data_in_frame[21][2] ), .I1(\data_in_frame[21][3] ), 
            .I2(n58672), .I3(GND_net), .O(n8_adj_5383));
    defparam i3_3_lut_adj_1249.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1250 (.I0(\data_in_frame[22] [6]), .I1(n61042), 
            .I2(n8_adj_5381), .I3(n26414), .O(n62972));
    defparam i1_4_lut_adj_1250.LUT_INIT = 16'h2112;
    SB_LUT4 i1_4_lut_adj_1251 (.I0(n62972), .I1(\data_in_frame[23] [4]), 
            .I2(n8_adj_5383), .I3(n58425), .O(n62974));
    defparam i1_4_lut_adj_1251.LUT_INIT = 16'h8228;
    SB_LUT4 i3_3_lut_adj_1252 (.I0(\data_in_frame[23] [3]), .I1(\data_in_frame[18] [5]), 
            .I2(n58663), .I3(GND_net), .O(n8_adj_5384));
    defparam i3_3_lut_adj_1252.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5385), .S(n57863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5386), .S(n57855));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5387), .S(n57854));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5388), .S(n57853));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5389), .S(n57852));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5390), .S(n57851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5391), .S(n57850));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5392), .S(n28997));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5393), .S(n57849));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5394), .S(n57848));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5395), .S(n57847));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5396), .S(n57846));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5397), .S(n57845));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5398), .S(n57844));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5399), .S(n57843));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5400), .S(n57842));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1253 (.I0(n5_adj_5401), .I1(n62974), .I2(\data_in_frame[22][5] ), 
            .I3(n58621), .O(n62976));
    defparam i1_4_lut_adj_1253.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1254 (.I0(n62976), .I1(n52807), .I2(n8_adj_5384), 
            .I3(n58400), .O(n62978));
    defparam i1_4_lut_adj_1254.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(\data_in_frame[23] [5]), .I1(n62978), 
            .I2(n58455), .I3(n61005), .O(n62980));
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[18]_c [2]), .I1(n58323), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5402));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1257 (.I0(n52776), .I1(\data_in_frame[20][3] ), 
            .I2(\data_in_frame[22][4] ), .I3(n6_adj_5402), .O(n59838));
    defparam i4_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1258 (.I0(n58269), .I1(n53750), .I2(\data_in_frame[20][0] ), 
            .I3(n58612), .O(n10_adj_5403));
    defparam i4_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1259 (.I0(n52879), .I1(n58403), .I2(n58458), 
            .I3(GND_net), .O(n8_adj_5404));
    defparam i3_3_lut_adj_1259.LUT_INIT = 16'h6969;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_18  (.CI(n51599), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n51600));
    SB_LUT4 i1_4_lut_adj_1260 (.I0(\data_in_frame[21][1] ), .I1(n59838), 
            .I2(\data_in_frame[23] [2]), .I3(n26087), .O(n62982));
    defparam i1_4_lut_adj_1260.LUT_INIT = 16'h4884;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_17_lut  (.I0(n66281), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n51598), .O(n28006)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1261 (.I0(\data_in_frame[21][5] ), .I1(n62980), 
            .I2(n58330), .I3(\data_in_frame[23] [6]), .O(n62984));
    defparam i1_4_lut_adj_1261.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1262 (.I0(\data_in_frame[22] [0]), .I1(n62982), 
            .I2(n8_adj_5404), .I3(\data_in_frame[19] [6]), .O(n62986));
    defparam i1_4_lut_adj_1262.LUT_INIT = 16'h8448;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_17  (.CI(n51598), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n51599));
    SB_LUT4 i2_3_lut_adj_1263 (.I0(n52853), .I1(n58208), .I2(\data_in_frame[23] [7]), 
            .I3(GND_net), .O(n60360));
    defparam i2_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1264 (.I0(\data_in_frame[15] [5]), .I1(n10_adj_5403), 
            .I2(\data_in_frame[22][1] ), .I3(GND_net), .O(n60585));
    defparam i5_3_lut_adj_1264.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5405), .S(n28988));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5406), .S(n57841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5407), .S(n57840));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5408), .S(n57839));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5409), .S(n57838));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5410), .S(n57837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5411), .S(n57836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5412), .S(n57835));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1265 (.I0(n58585), .I1(n52410), .I2(\data_in_frame[18] [5]), 
            .I3(\data_in_frame[22][7] ), .O(n63156));
    defparam i1_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5413), .S(n57834));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5414), .S(n57833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5415), .S(n57832));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5416), .S(n57831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5417), .S(n57830));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5418), .S(n57829));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5419), .S(n57828));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29805), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29804), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1266 (.I0(n58400), .I1(n58681), .I2(n63172), 
            .I3(n58269), .O(n63178));
    defparam i1_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1267 (.I0(n58179), .I1(n60893), .I2(\data_in_frame[17] [7]), 
            .I3(\data_in_frame[22][2] ), .O(n63216));
    defparam i1_4_lut_adj_1267.LUT_INIT = 16'h9669;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_16_lut  (.I0(n66256), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n51597), .O(n28008)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_16  (.CI(n51597), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n51598));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_15_lut  (.I0(n66255), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n51596), .O(n28010)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_15  (.CI(n51596), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n51597));
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5420), .S(n57827));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1268 (.I0(n60585), .I1(n60360), .I2(n62986), 
            .I3(n62984), .O(n62992));
    defparam i1_4_lut_adj_1268.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_adj_1269 (.I0(n58612), .I1(n62992), .I2(n58336), 
            .I3(n63216), .O(n62994));
    defparam i1_4_lut_adj_1269.LUT_INIT = 16'h8448;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_14_lut  (.I0(n66254), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n51595), .O(n28012)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1270 (.I0(n53861), .I1(n53829), .I2(n58211), 
            .I3(n63156), .O(n60661));
    defparam i1_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1271 (.I0(n58330), .I1(n58208), .I2(n58448), 
            .I3(n63178), .O(n63184));
    defparam i1_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1272 (.I0(n58323), .I1(n58621), .I2(\data_in_frame[20][1] ), 
            .I3(\data_in_frame[22][3] ), .O(n62930));
    defparam i1_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5421), .S(n57826));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1273 (.I0(n63184), .I1(n60661), .I2(n62994), 
            .I3(n58745), .O(n62998));
    defparam i1_4_lut_adj_1273.LUT_INIT = 16'h8040;
    SB_LUT4 i1_4_lut_adj_1274 (.I0(n62930), .I1(n25115), .I2(n58336), 
            .I3(\data_in_frame[19] [7]), .O(n60688));
    defparam i1_4_lut_adj_1274.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1275 (.I0(n53861), .I1(n58211), .I2(\data_in_frame[23] [0]), 
            .I3(GND_net), .O(n63144));
    defparam i1_3_lut_adj_1275.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1276 (.I0(n63144), .I1(n60688), .I2(n62998), 
            .I3(n53829), .O(Kp_23__N_612));
    defparam i1_4_lut_adj_1276.LUT_INIT = 16'h2010;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_14  (.CI(n51595), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n51596));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_13_lut  (.I0(n66253), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n51594), .O(n28014)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_13  (.CI(n51594), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n51595));
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29803), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i53608_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_612), 
            .I2(LED_N_3408), .I3(Kp_23__N_1748), .O(n27736));
    defparam i53608_4_lut.LUT_INIT = 16'hc4a0;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_12_lut  (.I0(n66252), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n51593), .O(n28016)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_12  (.CI(n51593), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n51594));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_11_lut  (.I0(n66250), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n51592), .O(n28018)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5422), .S(n57825));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5423), .S(n57824));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5424), .S(n57823));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i18_4_lut_adj_1277 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut_adj_1277.LUT_INIT = 16'hfffe;
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29802), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16_4_lut_adj_1278 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_5425));   // verilog/coms.v(157[7:23])
    defparam i16_4_lut_adj_1278.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1279 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(157[7:23])
    defparam i17_4_lut_adj_1279.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1280 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_5426));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut_adj_1280.LUT_INIT = 16'hfffe;
    SB_LUT4 add_1102_9_lut (.I0(n57901), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n50329), .O(n57909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_11  (.CI(n51592), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n51593));
    SB_LUT4 add_1102_8_lut (.I0(n57901), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n50328), .O(n57908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14_4_lut_adj_1281 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_5427));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut_adj_1281.LUT_INIT = 16'hfffe;
    SB_CARRY add_1102_8 (.CI(n50328), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n50329));
    SB_LUT4 add_1102_7_lut (.I0(n57901), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n50327), .O(n57907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_10_lut  (.I0(n66246), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n51591), .O(n28020)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29801), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29800), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29799), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_10  (.CI(n51591), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n51592));
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(157[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41_adj_5426), .I1(n43), .I2(n42_adj_5425), 
            .I3(n44), .O(n50));   // verilog/coms.v(157[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1282 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(157[7:23])
    defparam i19_4_lut_adj_1282.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40_adj_5427), 
            .O(n25529));   // verilog/coms.v(157[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28472_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25529), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i28472_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i465_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2068));   // verilog/coms.v(148[4] 304[11])
    defparam i465_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29798), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29797), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51670_3_lut (.I0(n101), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4942), 
            .I3(GND_net), .O(n66307));   // verilog/uart_tx.v(32[16:25])
    defparam i51670_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i51667_4_lut (.I0(n66307), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n66304));   // verilog/uart_tx.v(32[16:25])
    defparam i51667_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i30586_4_lut (.I0(r_SM_Main_2__N_3545[0]), .I1(n66304), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n44525));   // verilog/uart_tx.v(32[16:25])
    defparam i30586_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30587_3_lut (.I0(n44525), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n22192));   // verilog/uart_tx.v(32[16:25])
    defparam i30587_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1102_7 (.CI(n50327), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n50328));
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29796), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29795), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29794), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29793), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5429));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29792), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5430), .S(n57822));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1102_6_lut (.I0(n57901), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n50326), .O(n57906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_9_lut  (.I0(n66237), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n51590), .O(n28022)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5431), .S(n57821));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1102_6 (.CI(n50326), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n50327));
    SB_LUT4 add_1102_5_lut (.I0(n57901), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n50325), .O(n57905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_9  (.CI(n51590), .I0(n70121), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n51591));
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5432), .S(n57820));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1102_5 (.CI(n50325), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n50326));
    SB_LUT4 i30594_3_lut (.I0(n70210), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n44533));   // verilog/uart_tx.v(32[16:25])
    defparam i30594_3_lut.LUT_INIT = 16'hcbcb;
    SB_LUT4 add_1102_4_lut (.I0(n57901), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n50324), .O(n57904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i30601_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i30601_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_8_lut  (.I0(n66236), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n51589), .O(n28024)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\control_mode[0] ), .I1(n37407), .I2(GND_net), 
            .I3(GND_net), .O(n25541));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'heeee;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_8  (.CI(n51589), .I0(n70121), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n51590));
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5433), .S(n57819));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_7_lut  (.I0(n66231), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n51588), .O(n28026)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_7  (.CI(n51588), .I0(n70121), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n51589));
    SB_CARRY add_1102_4 (.CI(n50324), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n50325));
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5434), .S(n57818));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_6_lut  (.I0(n66224), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n51587), .O(n28028)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29791), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5435), .S(n57817));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29790), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5436), .S(n57734));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5437), .S(n57816));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1102_3_lut (.I0(n57901), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n50323), .O(n57903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_3_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5438), .S(n28960));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14015_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28045));   // verilog/coms.v(109[34:55])
    defparam i14015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48051_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63777));
    defparam i48051_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29789), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48052_4_lut (.I0(n63777), .I1(n28045), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63778));
    defparam i48052_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48050_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63776));
    defparam i48050_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5439), .S(n57815));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n29703));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5440), .S(n57814));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29787), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_6  (.CI(n51587), .I0(n70121), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n51588));
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5441), .S(n57813));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29786), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_5_lut  (.I0(n66221), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n51586), .O(n28030)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i2934081_i1_3_lut (.I0(n70222), .I1(n70450), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5338));
    defparam i2934081_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_5  (.CI(n51586), .I0(n70121), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n51587));
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29785), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29784), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1284 (.I0(control_mode[5]), .I1(control_mode_c[2]), 
            .I2(control_mode_c[3]), .I3(control_mode[6]), .O(n61023));   // verilog/coms.v(130[12] 305[6])
    defparam i1_4_lut_adj_1284.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1285 (.I0(control_mode[7]), .I1(n61023), .I2(control_mode_c[4]), 
            .I3(GND_net), .O(n37407));   // verilog/coms.v(130[12] 305[6])
    defparam i1_3_lut_adj_1285.LUT_INIT = 16'hfefe;
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29783), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5442));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_4_lut  (.I0(n66218), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n51585), .O(n28032)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29782), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29781), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_4  (.CI(n51585), .I0(n70121), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n51586));
    SB_CARRY add_1102_3 (.CI(n50323), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n50324));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_3_lut  (.I0(n66217), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n51584), .O(n28034)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1102_2_lut (.I0(n57901), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n57902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1102_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_3  (.CI(n51584), .I0(n70121), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n51585));
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29780), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29779), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1286 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [7]), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1286.LUT_INIT = 16'ha088;
    SB_LUT4 select_780_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29778), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5448));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29777), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29776), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i[0] ), 
            .CO(n51584));
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29775), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i52409_4_lut (.I0(n70156), .I1(n70282), .I2(byte_transmit_counter[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n68135));
    defparam i52409_4_lut.LUT_INIT = 16'h0aca;
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29774), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48157_3_lut (.I0(n70246), .I1(n68135), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i48157_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29773), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29772), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29771), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i52413_4_lut (.I0(n70150), .I1(n70288), .I2(byte_transmit_counter[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n68139));
    defparam i52413_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i48151_3_lut (.I0(n70240), .I1(n68139), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[4]));
    defparam i48151_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29770), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29769), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29768), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6624_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1951), 
            .I2(n60097), .I3(n4452), .O(n20323));   // verilog/coms.v(148[4] 304[11])
    defparam i6624_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1287 (.I0(n20323), .I1(n1951), .I2(n22692), .I3(n63421), 
            .O(n27016));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1287.LUT_INIT = 16'hbbba;
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29767), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29766), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i457_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2060));   // verilog/coms.v(148[4] 304[11])
    defparam i457_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29765), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29764), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29763), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29762), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29761), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29760), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29759), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29758), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29757), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29756), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29755), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47615_4_lut (.I0(n1951), .I1(n1954), .I2(n3303), .I3(n1957), 
            .O(n63325));   // verilog/coms.v(139[4] 141[7])
    defparam i47615_4_lut.LUT_INIT = 16'h0a02;
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29754), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29753), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1288 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1954), 
            .I2(n63325), .I3(n60837), .O(n57023));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1288.LUT_INIT = 16'hb3a0;
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29752), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29751), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n29709));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29749), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29748), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29747), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29746), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1102_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3416), .CO(n50323));
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29745), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6629_4_lut (.I0(n1955), .I1(\FRAME_MATCHER.state[3] ), .I2(n1957), 
            .I3(n25514), .O(n20328));   // verilog/coms.v(148[4] 304[11])
    defparam i6629_4_lut.LUT_INIT = 16'heccc;
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29744), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29743), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\byte_transmit_counter[0] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n25_c));   // verilog/coms.v(105[12:33])
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1290 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[3]), 
            .I2(n25_c), .I3(\byte_transmit_counter[2] ), .O(n61073));   // verilog/coms.v(105[12:33])
    defparam i2_4_lut_adj_1290.LUT_INIT = 16'h8880;
    SB_LUT4 i3_4_lut_adj_1291 (.I0(byte_transmit_counter[5]), .I1(n61073), 
            .I2(byte_transmit_counter[7]), .I3(byte_transmit_counter[6]), 
            .O(n97));   // verilog/coms.v(105[12:33])
    defparam i3_4_lut_adj_1291.LUT_INIT = 16'hfffe;
    SB_LUT4 i53661_3_lut (.I0(r_SM_Main_2__N_3545[0]), .I1(n97), .I2(tx_active), 
            .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i53661_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i446_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2049));   // verilog/coms.v(148[4] 304[11])
    defparam i446_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51722_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66217));   // verilog/coms.v(158[12:15])
    defparam i51722_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29742), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i445_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2048));   // verilog/coms.v(148[4] 304[11])
    defparam i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28471_4_lut (.I0(n8), .I1(\FRAME_MATCHER.i [31]), .I2(n25432), 
            .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i28471_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1292 (.I0(\FRAME_MATCHER.i [4]), .I1(n25529), .I2(GND_net), 
            .I3(GND_net), .O(n25432));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1292.LUT_INIT = 16'heeee;
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29741), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i28466_4_lut (.I0(n5_adj_5452), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i28466_4_lut.LUT_INIT = 16'h3332;
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29740), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29739), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29738), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51029_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66218));   // verilog/coms.v(158[12:15])
    defparam i51029_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_2_lut (.I0(n25514), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27593));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1293 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n22692));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1293.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_adj_1294 (.I0(n4452), .I1(n22692), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n27593), .O(n60943));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1294.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1295 (.I0(n25520), .I1(n1957), .I2(n1955), .I3(n60943), 
            .O(n27013));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1295.LUT_INIT = 16'hbaaa;
    SB_LUT4 i2_2_lut_adj_1296 (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5453));
    defparam i2_2_lut_adj_1296.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1297 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5454));
    defparam i6_4_lut_adj_1297.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1298 (.I0(\data_in[3] [6]), .I1(n14_adj_5454), 
            .I2(n10_adj_5453), .I3(\data_in[2] [1]), .O(n25552));
    defparam i7_4_lut_adj_1298.LUT_INIT = 16'hfffd;
    SB_LUT4 i47611_2_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n63320));
    defparam i47611_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut_adj_1299 (.I0(n25590), .I1(\data_in[2] [6]), .I2(\data_in[3] [7]), 
            .I3(n25552), .O(n21));
    defparam i8_4_lut_adj_1299.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(\data_in[3] [2]), .I1(\data_in[0] [1]), .I2(\data_in[1] [6]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i11_4_lut_adj_1300 (.I0(n21), .I1(n25526), .I2(n63320), .I3(\data_in[1] [3]), 
            .O(n24_adj_5455));
    defparam i11_4_lut_adj_1300.LUT_INIT = 16'hefff;
    SB_LUT4 i12_4_lut_adj_1301 (.I0(\data_in[0] [5]), .I1(n24_adj_5455), 
            .I2(n20), .I3(\data_in[2] [5]), .O(n1951));
    defparam i12_4_lut_adj_1301.LUT_INIT = 16'hfdff;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(\data_in[3] [0]), .I1(n25552), .I2(n25454), 
            .I3(\data_in[2] [2]), .O(n16_adj_5456));
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'hfffe;
    SB_LUT4 i50788_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66221));   // verilog/coms.v(158[12:15])
    defparam i50788_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1303 (.I0(\data_in[2] [4]), .I1(\data_in[1] [0]), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n17_adj_5457));
    defparam i7_4_lut_adj_1303.LUT_INIT = 16'hfffd;
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29737), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1304 (.I0(n17_adj_5457), .I1(\data_in[0] [6]), 
            .I2(n16_adj_5456), .I3(\data_in[1] [4]), .O(n1954));
    defparam i9_4_lut_adj_1304.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_4_lut_adj_1305 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [7]), 
            .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1305.LUT_INIT = 16'ha088;
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29736), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47822_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[1] [0]), .I2(\data_in[2] [2]), 
            .I3(\data_in[0] [3]), .O(n63539));
    defparam i47822_4_lut.LUT_INIT = 16'h8000;
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29735), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5458));
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'heeee;
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29734), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1307 (.I0(n9_adj_5458), .I1(n63539), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n25526));
    defparam i7_4_lut_adj_1307.LUT_INIT = 16'hffbf;
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n29729));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1308 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5459));
    defparam i4_4_lut_adj_1308.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1309 (.I0(\data_in[3] [4]), .I1(n10_adj_5459), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n25590));
    defparam i5_3_lut_adj_1309.LUT_INIT = 16'hdfdf;
    SB_LUT4 i7_4_lut_adj_1310 (.I0(\data_in[2] [6]), .I1(\data_in[1] [2]), 
            .I2(n25590), .I3(\data_in[3] [2]), .O(n18_c));
    defparam i7_4_lut_adj_1310.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1311 (.I0(\data_in[1] [6]), .I1(n18_c), .I2(\data_in[1] [3]), 
            .I3(\data_in[2] [0]), .O(n20_adj_5460));
    defparam i9_4_lut_adj_1311.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[2] [5]), .I1(\data_in[0] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5461));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_5461), .I1(n20_adj_5460), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [7]), .O(n25454));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 select_780_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1312 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n25454), .O(n16_adj_5462));
    defparam i6_4_lut_adj_1312.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1313 (.I0(n25526), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5463));
    defparam i7_4_lut_adj_1313.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1314 (.I0(n17_adj_5463), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5462), .I3(\data_in[3] [3]), .O(n1957));
    defparam i9_4_lut_adj_1314.LUT_INIT = 16'hfbff;
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29728));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i363_2_lut (.I0(n1954), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n1955));   // verilog/coms.v(142[4] 144[7])
    defparam i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n57968));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1316 (.I0(n57968), .I1(n1955), .I2(n1957), .I3(\FRAME_MATCHER.i_31__N_2507 ), 
            .O(n6_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1316.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1317 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [4]), 
            .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1317.LUT_INIT = 16'ha088;
    SB_LUT4 i3_4_lut_adj_1318 (.I0(n22691), .I1(n6_adj_5464), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n70526));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1318.LUT_INIT = 16'hefee;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29727));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1319 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [2]), 
            .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5436));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1319.LUT_INIT = 16'ha088;
    SB_LUT4 select_780_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29726));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29725));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29724));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29723));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29722));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29721));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29720));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i26_2_lut (.I0(n150), .I1(IntegralLimit[5]), .I2(GND_net), 
            .I3(GND_net), .O(n36515));   // verilog/TinyFPGA_B.v(248[22:35])
    defparam i26_2_lut.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29719));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29718));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50783_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66224));   // verilog/coms.v(158[12:15])
    defparam i50783_2_lut.LUT_INIT = 16'h2222;
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29717));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29716));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5434));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29715));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29714));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14352_3_lut (.I0(n42296), .I1(reset), .I2(n57974), .I3(GND_net), 
            .O(n58897));
    defparam i14352_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29713));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29712));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29708));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51256_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66231));   // verilog/coms.v(158[12:15])
    defparam i51256_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_780_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5465));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29702));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29701));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(\current_limit[2] ), .C(clk16MHz), .D(n29697));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_780_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n29695), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n29694), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n29693), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n29692), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n29691), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5303), .S(n57812));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5301), .S(n57811));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n29690), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5300), .S(n57810));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5299), .S(n57809));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n29689), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15566_3_lut (.I0(\data_in_frame[3]_c [6]), .I1(rx_data[6]), 
            .I2(n58929), .I3(GND_net), .O(n29597));   // verilog/coms.v(130[12] 305[6])
    defparam i15566_3_lut.LUT_INIT = 16'hacac;
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n29688), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n29687), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n29686), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n29685), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5293), .S(n57808));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n29684), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5292), .S(n57807));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5291), .S(n57806));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5290), .S(n57805));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n29683), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n29682), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29681), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit_c[15]), .C(clk16MHz), 
           .D(n29680));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit_c[14]), .C(clk16MHz), 
           .D(n29679));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit_c[13]), .C(clk16MHz), 
           .D(n29678));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(\current_limit[12] ), .C(clk16MHz), 
           .D(n29677));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5287), .S(n57804));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5284), .S(n57803));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(\current_limit[11] ), .C(clk16MHz), 
           .D(n29676));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29675));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(\current_limit[9] ), .C(clk16MHz), .D(n29674));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(\current_limit[8] ), .C(clk16MHz), .D(n29673));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(\current_limit[7] ), .C(clk16MHz), .D(n29671));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5281), .S(n57735));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5280), .S(n57736));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n29670));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5277), .S(n57737));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5276), .S(n57738));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(\current_limit[5] ), .C(clk16MHz), .D(n29669));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5275), .S(n57739));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(\current_limit[3] ), .C(clk16MHz), .D(n29666));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5273), .S(n57740));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5473), .S(n28940));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i20996_3_lut (.I0(n58929), .I1(rx_data[4]), .I2(\data_in_frame[3]_c [4]), 
            .I3(GND_net), .O(n29956));   // verilog/coms.v(94[13:20])
    defparam i20996_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[0][0] ), 
            .I2(\data_in_frame[2][1] ), .I3(GND_net), .O(n58075));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5474));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29655));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29654));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5475), .S(n57741));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5476), .S(n57742));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5477), .S(n57743));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29651));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[0][0] ), 
            .I2(n25806), .I3(Kp_23__N_748), .O(n24_adj_5478));   // verilog/coms.v(73[16:69])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0906;
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29650));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(\control_mode[1] ), .C(clk16MHz), .D(n29649));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode_c[2]), .C(clk16MHz), .D(n29648));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode_c[3]), .C(clk16MHz), .D(n29647));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5479), .S(n57744));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5480), .S(n57745));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode_c[4]), .C(clk16MHz), .D(n29638));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0][5] ), .I3(\data_in_frame[0]_c [7]), .O(n58223));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n29630));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29629));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_2_lut_3_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n25813));   // verilog/coms.v(99[12:25])
    defparam i11_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i53555_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[2] [7]), .I2(n7), 
            .I3(GND_net), .O(n57285));   // verilog/coms.v(94[13:20])
    defparam i53555_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5482), .S(n57746));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5483), .S(n57747));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n30552), .D(n2_adj_5484), .S(n28932));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5485), .S(n57748));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_302_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8));   // verilog/coms.v(157[7:23])
    defparam equal_302_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_301_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_8));   // verilog/coms.v(157[7:23])
    defparam equal_301_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i48068_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63794));
    defparam i48068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48069_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63795));
    defparam i48069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48075_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63801));
    defparam i48075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48074_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63800));
    defparam i48074_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29618), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(\current_limit[0] ), .C(clk16MHz), .D(n29617));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(\control_mode[0] ), .C(clk16MHz), .D(n29616));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29615));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29614), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29613), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29612), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5487), .S(n57749));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47927_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63653));
    defparam i47927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47928_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63654));
    defparam i47928_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5488), .S(n57750));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5489), .S(n57751));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5490), .S(n57752));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5491), .S(n57753));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5492), .S(n57754));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n30561), .D(n2_adj_5493), .S(n28924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5494), .S(n57755));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5495), .S(n57756));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5496), .S(n57757));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5497), .S(n57758));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5498), .S(n57759));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5499), .S(n57760));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48003_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63729));
    defparam i48003_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n30568), .D(n2_adj_5500), .S(n28917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5501), .S(n41));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5503), .S(n57761));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5504), .S(n57762));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48002_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63728));
    defparam i48002_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5505), .S(n57763));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5506), .S(n25));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5508), .S(n28911));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5509), .S(n28910));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5510), .S(n57764));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5511), .S(n57765));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5512), .S(n57766));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5513), .S(n57767));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5514), .S(n57768));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5515), .S(n57769));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5516), .S(n57770));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5517), .S(n57771));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5518), .S(n57772));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5519), .S(n57773));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48116_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63842));
    defparam i48116_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5520), .S(n57774));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5521), .S(n57775));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5522), .S(n57776));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48117_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63843));
    defparam i48117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47931_3_lut (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63657));
    defparam i47931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47930_3_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[21] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63656));
    defparam i47930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48107_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63833));
    defparam i48107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48108_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63834));
    defparam i48108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48045_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63771));
    defparam i48045_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR \FRAME_MATCHER.i_1943__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n27972), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5523), .S(n57777));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5524), .S(n57778));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48044_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63770));
    defparam i48044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1320 (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n101));
    defparam i2_3_lut_adj_1320.LUT_INIT = 16'h8080;
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5525), .S(n57779));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1943__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n27974), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n27976), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_4_lut_adj_1321 (.I0(n58909), .I1(n59553), .I2(r_SM_Main[1]), 
            .I3(n101), .O(n29148));
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'h1101;
    SB_LUT4 i51507_2_lut (.I0(\byte_transmit_counter[0] ), .I1(\data_out_frame[0][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66400));
    defparam i51507_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i48042_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63768));
    defparam i48042_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR \FRAME_MATCHER.i_1943__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n27978), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n27980), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n27982), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n27984), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n27986), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n27988), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n27990), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n27992), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n27994), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n27996), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n27998), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28000), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28002), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28004), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28006), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28008), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28010), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28012), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28014), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28016), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28018), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28020), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28022), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28024), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n28026), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n28028), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n28030), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n28032), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1943__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n28034), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5526), .S(n28893));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i39_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i21260_4_lut_4_lut (.I0(n42499), .I1(reset), .I2(\data_in_frame[23] [7]), 
            .I3(rx_data[7]), .O(n30068));
    defparam i21260_4_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_780_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48043_4_lut (.I0(n63768), .I1(n66400), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[1]), .O(n63769));
    defparam i48043_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i50945_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66294));   // verilog/coms.v(158[12:15])
    defparam i50945_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48041_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63767));
    defparam i48041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15519_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n29550));
    defparam i15519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2935287_i1_3_lut (.I0(n70198), .I1(n70480), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5527));
    defparam i2935287_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48098_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63824));
    defparam i48098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50791_2_lut (.I0(n70258), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66456));
    defparam i50791_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15516_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n29547));
    defparam i15516_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i48099_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63825));
    defparam i48099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15504_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n29535));
    defparam i15504_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i48084_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63810));
    defparam i48084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48083_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63809));
    defparam i48083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15501_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n29532));
    defparam i15501_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5528), .S(n57899));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15498_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n29529));
    defparam i15498_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5529), .S(n57898));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48086_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63812));
    defparam i48086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48087_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63813));
    defparam i48087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15495_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n29526));
    defparam i15495_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15492_3_lut_4_lut (.I0(n42499), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n29523));
    defparam i15492_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i48093_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63819));
    defparam i48093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(reset), .I1(n57974), .I2(n8), 
            .I3(GND_net), .O(n58008));
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'hfefe;
    SB_LUT4 i48092_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63818));
    defparam i48092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48059_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63785));
    defparam i48059_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF current_limit_i0_i4 (.Q(\current_limit[4] ), .C(clk16MHz), .D(n30452));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18]_c [2]), .C(clk16MHz), 
           .D(n57109));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n30441));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18][3] ), .C(clk16MHz), 
           .D(n57237));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48060_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63786));
    defparam i48060_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18][4] ), .C(clk16MHz), 
           .D(n57235));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n57233));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(reset), .I1(n57974), .I2(n8_adj_9), 
            .I3(GND_net), .O(n58010));
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18]_c [6]), .C(clk16MHz), 
           .D(n57129));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18][7] ), .C(clk16MHz), 
           .D(n57229));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29385));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29388));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i146 (.Q(\data_in_frame[18][1] ), .C(clk16MHz), 
            .E(VCC_net), .D(n57179));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n29895));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29391));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29394));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19]_c [4]), .C(clk16MHz), 
           .D(n14_adj_5531));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30408), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48147_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63873));
    defparam i48147_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n36387), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0][4] ), .C(clk16MHz), 
           .D(n29404));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30353));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30352));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30351));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30350));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30349));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30348));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30347));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30346));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30345));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30344));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30343));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30342));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30341));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30340));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30339));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48146_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63872));
    defparam i48146_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30338));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30337));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30336));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30335));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30334));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30333));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30332));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30331));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30330));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30329));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30328));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30327));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30326));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30325));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30324));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30323));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30322), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19]_c [5]), .C(clk16MHz), 
           .D(n17_adj_5532));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n29898));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n29901));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29410));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29413));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7]_c [6]), .C(clk16MHz), 
           .D(n57325));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30315), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i145 (.Q(\data_in_frame[18][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n57183));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20][0] ), .C(clk16MHz), 
           .D(n29416));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20][1] ), .C(clk16MHz), 
           .D(n29420));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n25_adj_5533));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20][3] ), .C(clk16MHz), 
           .D(n29427));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20][4] ), .C(clk16MHz), 
           .D(n29430));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n9_adj_5534));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n29436));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n57449));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0][5] ), .C(clk16MHz), 
           .D(n29442));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0]_c [6]), .C(clk16MHz), 
           .D(n29445));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0]_c [7]), .C(clk16MHz), 
           .D(n29448));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1]_c [0]), .C(clk16MHz), 
           .D(n29451));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7]_c [7]), .C(clk16MHz), 
           .D(n57319));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8]_c [0]), .C(clk16MHz), 
           .D(n29911));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8]_c [1]), .C(clk16MHz), 
           .D(n29915));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1]_c [1]), .C(clk16MHz), 
           .D(n57379));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30295), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30290), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1][2] ), .C(clk16MHz), 
           .D(n57383));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1]_c [3]), .C(clk16MHz), 
           .D(n29460));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1]_c [4]), .C(clk16MHz), 
           .D(n29463));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n29918));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8][3] ), .C(clk16MHz), 
           .D(n29921));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
           .D(n29925));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8]_c [5]), .C(clk16MHz), 
           .D(n29928));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8][6] ), .C(clk16MHz), 
           .D(n29931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30275), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8]_c [7]), .C(clk16MHz), 
           .D(n29934));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n29937));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n29941));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n29944));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n29947));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n29466));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1][6] ), .C(clk16MHz), 
           .D(n29469));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n29950));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n29953));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n29957));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9][7] ), .C(clk16MHz), 
           .D(n29960));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
           .D(n29963));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
           .D(n29967));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
           .D(n29970));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
           .D(n29973));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n29977));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
           .D(n29980));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n29983));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n29987));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n29990));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n29993));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11][2] ), .C(clk16MHz), 
           .D(n57277));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n30000));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n57339));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n30007));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n30010));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30013));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30017));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51691_2_lut (.I0(n70270), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66234));
    defparam i51691_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30246), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12]_c [1]), .C(clk16MHz), 
           .D(n30020));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12]_c [2]), .C(clk16MHz), 
           .D(n30023));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12]_c [3]), .C(clk16MHz), 
           .D(n30027));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12]_c [4]), .C(clk16MHz), 
           .D(n30030));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12]_c [5]), .C(clk16MHz), 
           .D(n30033));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12]_c [6]), .C(clk16MHz), 
           .D(n30037));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12]_c [7]), .C(clk16MHz), 
           .D(n30040));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n30043));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50979_2_lut (.I0(\data_out_frame[1][5] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n66436));
    defparam i50979_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(reset), .I1(n57974), .I2(n8_adj_5535), 
            .I3(GND_net), .O(n58011));
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30047));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n30050));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30053));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n30056));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n30059));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n30062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n30065));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n30069));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n57355));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
           .D(n30075));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
           .D(n30079));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n30082));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n30085));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n30089));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n30092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n30095));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n30099));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n30102));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n30105));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n30109));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n30112));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n30115));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n30119));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n57225));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n57223));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n57221));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n57219));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n57215));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n57211));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n57207));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n57203));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n30149));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1325 (.I0(reset), .I1(n57974), .I2(n8_adj_5536), 
            .I3(GND_net), .O(n58009));
    defparam i1_2_lut_3_lut_adj_1325.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17]_c [1]), .C(clk16MHz), 
           .D(n57239));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17]_c [2]), .C(clk16MHz), 
           .D(n57241));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17][3] ), .C(clk16MHz), 
           .D(n57199));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17][4] ), .C(clk16MHz), 
           .D(n57195));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17][5] ), .C(clk16MHz), 
           .D(n57191));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17][6] ), .C(clk16MHz), 
           .D(n30169));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n57187));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21][0] ), .C(clk16MHz), 
           .D(n57117));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1][7] ), .C(clk16MHz), 
           .D(n29475));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21][1] ), .C(clk16MHz), 
           .D(n57169));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21][2] ), .C(clk16MHz), 
           .D(n57167));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21][3] ), .C(clk16MHz), 
           .D(n57163));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21][4] ), .C(clk16MHz), 
           .D(n57159));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21][5] ), .C(clk16MHz), 
           .D(n57155));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n57125));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21][7] ), .C(clk16MHz), 
           .D(n57127));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n57269));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22][1] ), .C(clk16MHz), 
           .D(n29502));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22][2] ), .C(clk16MHz), 
           .D(n29505));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22][3] ), .C(clk16MHz), 
           .D(n29508));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22][4] ), .C(clk16MHz), 
           .D(n29511));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22][5] ), .C(clk16MHz), 
           .D(n29514));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n30176));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22][7] ), .C(clk16MHz), 
           .D(n29520));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29523));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29526));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n29529));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48030_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63756));
    defparam i48030_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5537), .S(n57897));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29532));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_306_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5536));   // verilog/coms.v(157[7:23])
    defparam equal_306_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29535));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2][0] ), .C(clk16MHz), 
           .D(n29538));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_305_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_9));   // verilog/coms.v(157[7:23])
    defparam equal_305_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i51271_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66236));   // verilog/coms.v(158[12:15])
    defparam i51271_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48031_4_lut (.I0(n63756), .I1(n66436), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63757));
    defparam i48031_4_lut.LUT_INIT = 16'haca0;
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2][1] ), .C(clk16MHz), 
           .D(n29541));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n58889), .I3(\FRAME_MATCHER.i [3]), .O(n57974));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n29544));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48029_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63755));
    defparam i48029_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29547));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5538), .S(n57896));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n29550));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n30068));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2][3] ), .C(clk16MHz), 
           .D(n29560));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_4_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[6] [3]), .O(n1244));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n58889), .I3(\FRAME_MATCHER.i [3]), .O(n57993));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'hefff;
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n57341));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5539), .S(n57895));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2][5] ), .C(clk16MHz), 
           .D(n29566));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i53556_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[2] [6]), .I2(n7), 
            .I3(GND_net), .O(n57303));   // verilog/coms.v(94[13:20])
    defparam i53556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_780_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5540));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5541), .S(n57894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5540), .S(n57893));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n57303));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54662 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[6] [4]), .I2(\data_out_frame[7] [4]), .I3(byte_transmit_counter[1]), 
            .O(n70315));
    defparam byte_transmit_counter_0__bdd_4_lut_54662.LUT_INIT = 16'he4aa;
    SB_LUT4 i51155_2_lut (.I0(n70294), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66457));
    defparam i51155_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n57285));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
           .D(n29575));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5541));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n29578));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
           .D(n29581));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14009_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28039));   // verilog/coms.v(109[34:55])
    defparam i14009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48024_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63750));
    defparam i48024_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
           .D(n29584));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5474), .S(n57892));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3]_c [4]), .C(clk16MHz), 
           .D(n29956));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5472), .S(n57891));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48025_4_lut (.I0(n63750), .I1(n28039), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63751));
    defparam i48025_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i53560_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[2] [4]), .I2(n7), 
            .I3(GND_net), .O(n57341));   // verilog/coms.v(94[13:20])
    defparam i53560_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3][5] ), .C(clk16MHz), 
           .D(n29592));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48023_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63749));
    defparam i48023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n70315_bdd_4_lut (.I0(n70315), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(byte_transmit_counter[1]), 
            .O(n63732));
    defparam n70315_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3]_c [6]), .C(clk16MHz), 
           .D(n29597));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5471), .S(n57890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5470), .S(n57889));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5469), .S(n57888));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5468), .S(n57887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5467), .S(n57886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5466), .S(n57885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5465), .S(n57884));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1327 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\data_out_frame[1][0] ), .I3(GND_net), .O(n2_adj_5538));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1327.LUT_INIT = 16'ha8a8;
    SB_LUT4 i51129_2_lut (.I0(n70300), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66439));
    defparam i51129_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15513_3_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), .I2(n7), 
            .I3(GND_net), .O(n29544));   // verilog/coms.v(130[12] 305[6])
    defparam i15513_3_lut.LUT_INIT = 16'hacac;
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3][7] ), .C(clk16MHz), 
           .D(n29600));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n29423));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29419), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47924_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63650));
    defparam i47924_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27736), 
            .D(n4764[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47925_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63651));
    defparam i47925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48171_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63897));
    defparam i48171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48170_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63896));
    defparam i48170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48110_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63836));
    defparam i48110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_780_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27736), 
            .D(n4764[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27736), 
            .D(n4764[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27736), 
            .D(n4764[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27736), 
            .D(n4764[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27736), 
            .D(n4764[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27736), 
            .D(n4764[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27736), 
            .D(n4764[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27736), 
            .D(n4764[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27736), 
            .D(n4764[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27736), 
            .D(n4764[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27736), 
            .D(n4764[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27736), 
            .D(n4764[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27736), 
            .D(n4764[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27736), 
            .D(n4764[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27736), 
            .D(n4764[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27736), 
            .D(n4764[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27736), 
            .D(n4764[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27736), 
            .D(n4764[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27736), 
            .D(n4764[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27736), 
            .D(n4764[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27736), 
            .D(n4764[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27736), 
            .D(n4764[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n70526), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i48111_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63837));
    defparam i48111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48021_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63747));
    defparam i48021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(n42296), .I1(n40525), .I2(GND_net), 
            .I3(GND_net), .O(n42499));
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h8888;
    SB_LUT4 i48020_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63746));
    defparam i48020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48005_4_lut (.I0(\byte_transmit_counter[0] ), .I1(\data_out_frame[3][4] ), 
            .I2(byte_transmit_counter[1]), .I3(\data_out_frame[0][4] ), 
            .O(n63731));
    defparam i48005_4_lut.LUT_INIT = 16'h8580;
    SB_LUT4 select_780_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54554 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(byte_transmit_counter[1]), 
            .O(n70309));
    defparam byte_transmit_counter_0__bdd_4_lut_54554.LUT_INIT = 16'he4aa;
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n27013), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2048), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2049), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20328), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n57023), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2060), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n27016), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i21420_3_lut (.I0(n28352), .I1(rx_data[6]), .I2(\data_in_frame[22] [6]), 
            .I3(GND_net), .O(n30176));   // verilog/coms.v(94[13:20])
    defparam i21420_3_lut.LUT_INIT = 16'he4e4;
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5450), .S(n57883));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5449), .S(n57882));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5448), .S(n57881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5447), .S(n57880));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5446), .S(n57879));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1329 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n58004), .I3(LED_c), .O(n27276));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1329.LUT_INIT = 16'hfe00;
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n29603));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n30680), .D(n2_adj_5445), .S(n29037));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n70309_bdd_4_lut (.I0(n70309), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(byte_transmit_counter[1]), 
            .O(n63735));
    defparam n70309_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5444), .S(n57780));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3472));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48008_4_lut (.I0(n1), .I1(\data_out_frame[3][3] ), .I2(byte_transmit_counter[1]), 
            .I3(\byte_transmit_counter[0] ), .O(n63734));
    defparam i48008_4_lut.LUT_INIT = 16'hca0a;
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5443), .S(n57781));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14007_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28037));   // verilog/coms.v(109[34:55])
    defparam i14007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48012_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63738));
    defparam i48012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48013_4_lut (.I0(n63738), .I1(n28037), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63739));
    defparam i48013_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 select_780_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5442), .S(n57782));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48011_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63737));
    defparam i48011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14322_4_lut (.I0(n40523), .I1(reset), .I2(n58889), .I3(n8_adj_5535), 
            .O(n28352));
    defparam i14322_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i11_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[22] [0]), .I2(n28352), 
            .I3(GND_net), .O(n57269));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50790_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66237));   // verilog/coms.v(158[12:15])
    defparam i50790_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_780_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5430));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15578_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n58009), 
            .I3(GND_net), .O(n29609));   // verilog/coms.v(130[12] 305[6])
    defparam i15578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 select_780_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5264));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i29412117_i1_3_lut (.I0(n70216), .I1(n70462), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5542));
    defparam i29412117_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48182_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63908));
    defparam i48182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1331 (.I0(\data_in_frame[21][7] ), .I1(n40525), 
            .I2(n28355), .I3(rx_data[7]), .O(n57127));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1331.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_1332 (.I0(\data_in_frame[21] [6]), .I1(n40525), 
            .I2(n28355), .I3(rx_data[6]), .O(n57125));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1332.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n57923));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1333 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n57924));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1333.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[18] [0]), 
            .I2(n10_adj_5543), .I3(\data_out_frame[16] [0]), .O(n52835));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1334 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n57925));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1334.LUT_INIT = 16'h5100;
    SB_LUT4 i48183_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63909));
    defparam i48183_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5429), .S(n57783));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50869_2_lut (.I0(n70306), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66247));
    defparam i50869_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5382), .S(n57878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n30686), .D(n2_adj_5380), .S(n29035));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n30687), .D(n2_adj_5379), .S(n29034));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5378), .S(n57877));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n30689), .D(n2_adj_5375), .S(n29032));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5374), .S(n57876));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n30691), .D(n2_adj_5373), .S(n29030));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5369), .S(n57875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5367), .S(n57874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5366), .S(n57873));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5365), .S(n57872));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5364), .S(n57871));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5363), .S(n57870));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5362), .S(n57869));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5361), .S(n57868));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5360), .S(n57867));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5359), .S(n57866));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5358), .S(n57865));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5357), .S(n57864));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n29403));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5356), .S(n57784));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(\current_limit[1] ), .C(clk16MHz), .D(n29401));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1335 (.I0(\data_out_frame[20] [4]), .I1(n53875), 
            .I2(\data_out_frame[22] [5]), .I3(GND_net), .O(n58346));
    defparam i1_2_lut_3_lut_adj_1335.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1336 (.I0(\data_out_frame[20] [4]), .I1(n53875), 
            .I2(\data_out_frame[20] [5]), .I3(GND_net), .O(n53785));
    defparam i1_2_lut_3_lut_adj_1336.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5355), .S(n57785));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2][5] ), .I3(\data_in_frame[0][4] ), .O(n26667));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1337 (.I0(n53787), .I1(n58346), .I2(\data_out_frame[25] [1]), 
            .I3(\data_out_frame[25] [2]), .O(n58639));
    defparam i2_3_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i48162_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63888));
    defparam i48162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1338 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n57911));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1338.LUT_INIT = 16'h5100;
    SB_LUT4 i48161_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63887));
    defparam i48161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1339 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0][0] ), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n26371));   // verilog/coms.v(76[16:42])
    defparam i1_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i51701_4_lut (.I0(\data_out_frame[6] [0]), .I1(\byte_transmit_counter[2] ), 
            .I2(\data_out_frame[7] [0]), .I3(\byte_transmit_counter[0] ), 
            .O(n66502));   // verilog/coms.v(105[12:33])
    defparam i51701_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1340 (.I0(ID[7]), .I1(\data_in_frame[0][5] ), .I2(\data_in_frame[0]_c [7]), 
            .I3(ID[5]), .O(n12_adj_5544));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1340.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1341 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0][4] ), 
            .I2(ID[2]), .I3(ID[4]), .O(n10_adj_5545));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1341.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1342 (.I0(ID[6]), .I1(\data_in_frame[0] [1]), .I2(\data_in_frame[0]_c [6]), 
            .I3(ID[1]), .O(n11));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1342.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1343 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5546));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1343.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1344 (.I0(n9_adj_5546), .I1(n11), .I2(n10_adj_5545), 
            .I3(n12_adj_5544), .O(n61042));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1344.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\data_in_frame[0]_c [6]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58266));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1346 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2][3] ), .I3(GND_net), .O(n26343));   // verilog/coms.v(78[16:43])
    defparam i1_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1347 (.I0(\data_in_frame[0]_c [6]), .I1(\data_in_frame[1]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58065));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1347.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1348 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0][4] ), 
            .I2(\data_in_frame[0][5] ), .I3(GND_net), .O(n26663));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1348.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1349 (.I0(\data_in_frame[2][5] ), .I1(\data_in_frame[0][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n58084));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1349.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1350 (.I0(\data_in_frame[0][4] ), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0]_c [6]), .I3(n58223), .O(Kp_23__N_748));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1351 (.I0(\data_in_frame[2][0] ), .I1(\data_in_frame[0][0] ), 
            .I2(Kp_23__N_748), .I3(GND_net), .O(n60617));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1352 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n57926));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1352.LUT_INIT = 16'h5100;
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5354), .S(n57786));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1353 (.I0(n25813), .I1(Kp_23__N_748), .I2(\data_in_frame[2][1] ), 
            .I3(GND_net), .O(n22));
    defparam i5_3_lut_adj_1353.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1354 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[1][2] ), .I3(\data_in_frame[1]_c [4]), .O(n27_adj_5547));
    defparam i10_4_lut_adj_1354.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut_adj_1355 (.I0(n60617), .I1(\data_in_frame[0]_c [7]), 
            .I2(\data_in_frame[1][6] ), .I3(\data_in_frame[1]_c [1]), .O(n26_adj_5548));
    defparam i9_4_lut_adj_1355.LUT_INIT = 16'h4010;
    SB_LUT4 i12_4_lut_adj_1356 (.I0(n26663), .I1(n24_adj_5478), .I2(\data_in_frame[0]_c [7]), 
            .I3(n58065), .O(n29_adj_5549));
    defparam i12_4_lut_adj_1356.LUT_INIT = 16'h0440;
    SB_LUT4 i14_4_lut_adj_1357 (.I0(n27_adj_5547), .I1(n61042), .I2(n22), 
            .I3(n26371), .O(n31));
    defparam i14_4_lut_adj_1357.LUT_INIT = 16'h0020;
    SB_LUT4 i16_4_lut_adj_1358 (.I0(n31), .I1(n29_adj_5549), .I2(n63337), 
            .I3(n26_adj_5548), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1358.LUT_INIT = 16'h0800;
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5353), .S(n57787));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51666_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66246));   // verilog/coms.v(158[12:15])
    defparam i51666_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i29_4_lut (.I0(\data_out_frame[1][0] ), .I1(n66502), .I2(byte_transmit_counter[1]), 
            .I3(\byte_transmit_counter[0] ), .O(n10_adj_5550));   // verilog/coms.v(105[12:33])
    defparam i29_4_lut.LUT_INIT = 16'hcac0;
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5352), .S(n57788));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5351), .S(n57789));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5350), .S(n57790));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5349), .S(n57791));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5348), .S(n57792));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5347), .S(n57793));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5346), .S(n57794));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5344), .S(n57795));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5343), .S(n57796));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n30717), .D(n2_adj_5341), .S(n29017));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i21471_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n4_adj_5551));   // verilog/coms.v(105[12:33])
    defparam i21471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1359 (.I0(\data_out_frame[16] [6]), .I1(n26872), 
            .I2(\data_out_frame[16] [7]), .I3(\data_out_frame[19] [2]), 
            .O(n6_adj_5278));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n30718), .D(n2_adj_5336), .S(n29016));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n30719), .D(n2_adj_5335), .S(n29015));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5334), .S(n57862));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5333), .S(n57797));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5332), .S(n57733));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5331), .S(n57798));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5330), .S(n57799));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5329), .S(n57800));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5328), .S(n57801));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5327), .S(n57802));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5326), .S(n57912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2874), .D(n3), .S(n57913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5552), .S(n57914));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5553), .S(n57915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5554), .S(n57916));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5555), .S(n57917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5556), .S(n57918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5557), .S(n57919));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5558), .S(n57920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5559), .S(n57921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5560), .S(n57922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5561), .S(n57923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5562), .S(n57924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5563), .S(n57925));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5564), .S(n57911));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2874), .D(n3_adj_5565), .S(n57926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5566), .S(n57903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5567), .S(n57904));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5568), .S(n57905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5569), .S(n57906));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5570), .S(n57907));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5571), .S(n57908));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n2874), .D(n86), .S(n57909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2874), .D(n1_adj_5572), .S(n28829));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2874), .D(n5_adj_5573), 
            .S(n28828));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2874), .D(n26923), 
            .S(n28827));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1360 (.I0(current_limit_c[14]), .I1(current_limit_c[15]), 
            .I2(n26), .I3(current_limit_c[13]), .O(n18));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i1_4_lut_adj_1360.LUT_INIT = 16'h3332;
    SB_LUT4 i11_4_lut_adj_1361 (.I0(\data_in_frame[17]_c [2]), .I1(n40525), 
            .I2(n28363), .I3(rx_data[2]), .O(n57241));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1361.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_1362 (.I0(\data_in_frame[17]_c [1]), .I1(n40525), 
            .I2(n28363), .I3(rx_data[1]), .O(n57239));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1362.LUT_INIT = 16'hca0a;
    SB_LUT4 select_780_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5424));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(clk16MHz), .E(n2874), .D(n1_adj_5576), .S(n57902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n30778), .D(n2_adj_5577), .S(n29013));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n30779), .D(n2_adj_5578), .S(n29012));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2874), .D(n2_adj_5579), .S(n57861));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_780_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5423));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54549 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n70303));
    defparam byte_transmit_counter_0__bdd_4_lut_54549.LUT_INIT = 16'he4aa;
    SB_LUT4 i50849_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66250));   // verilog/coms.v(158[12:15])
    defparam i50849_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n70303_bdd_4_lut (.I0(n70303), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n70306));
    defparam n70303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54544 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n70297));
    defparam byte_transmit_counter_0__bdd_4_lut_54544.LUT_INIT = 16'he4aa;
    SB_LUT4 n70297_bdd_4_lut (.I0(n70297), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n70300));
    defparam n70297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1363 (.I0(n4_adj_5342), .I1(n26829), 
            .I2(\data_in_frame[8] [2]), .I3(n25933), .O(n58229));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut (.I0(n52743), .I1(n58575), .I2(n52790), .I3(n53902), 
            .O(n8_adj_5580));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(n52743), .I1(n58575), .I2(n52831), 
            .I3(GND_net), .O(n58731));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 i50964_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66310));   // verilog/coms.v(158[12:15])
    defparam i50964_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50892_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66252));   // verilog/coms.v(158[12:15])
    defparam i50892_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50940_3_lut (.I0(current_limit_c[14]), .I1(n26), .I2(current_limit_c[13]), 
            .I3(GND_net), .O(n66289));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i50940_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i23543_4_lut (.I0(n18), .I1(n66289), .I2(\current[15] ), .I3(current_limit_c[15]), 
            .O(n260));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i23543_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i50968_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66312));   // verilog/coms.v(158[12:15])
    defparam i50968_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50836_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66253));   // verilog/coms.v(158[12:15])
    defparam i50836_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50972_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66313));   // verilog/coms.v(158[12:15])
    defparam i50972_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_780_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5421));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i50837_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66254));   // verilog/coms.v(158[12:15])
    defparam i50837_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_33_lut  (.I0(n66361), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n51614), .O(n27974)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_780_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5420));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i50840_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66255));   // verilog/coms.v(158[12:15])
    defparam i50840_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50987_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66323));   // verilog/coms.v(158[12:15])
    defparam i50987_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_782_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5576));   // verilog/coms.v(148[4] 304[11])
    defparam select_782_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n58562));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n58004));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1367 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [1]), .I3(\data_out_frame[20] [2]), 
            .O(n58183));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i50842_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66256));   // verilog/coms.v(158[12:15])
    defparam i50842_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[7]), .I3(GND_net), .O(n86));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[6]), .I3(GND_net), .O(n1_adj_5571));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(n8_adj_5535), .I1(n57993), .I2(GND_net), 
            .I3(GND_net), .O(n28314));
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n1_adj_5570));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1372 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[4]), .I3(GND_net), .O(n1_adj_5569));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1372.LUT_INIT = 16'h1010;
    SB_LUT4 select_782_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n1_adj_5567));   // verilog/coms.v(148[4] 304[11])
    defparam select_782_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_32_lut  (.I0(n66356), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n51613), .O(n27976)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_32  (.CI(n51613), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n51614));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_31_lut  (.I0(n66355), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n51612), .O(n27978)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i51000_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66324));   // verilog/coms.v(158[12:15])
    defparam i51000_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(byte_transmit_counter[3]), .I3(GND_net), .O(n1_adj_5568));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'h1010;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_31  (.CI(n51612), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n51613));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_30_lut  (.I0(n66354), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n51611), .O(n27980)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_30  (.CI(n51611), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n51612));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_29_lut  (.I0(n66350), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n51610), .O(n27982)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(\data_out_frame[21] [7]), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n8_adj_5581));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_29  (.CI(n51610), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n51611));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_28_lut  (.I0(n66347), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n51609), .O(n27984)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_782_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_adj_5566));   // verilog/coms.v(148[4] 304[11])
    defparam select_782_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_28  (.CI(n51609), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n51610));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_27_lut  (.I0(n66324), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n51608), .O(n27986)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_27  (.CI(n51608), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n51609));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_26_lut  (.I0(n66323), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n51607), .O(n27988)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_26  (.CI(n51607), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n51608));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_25_lut  (.I0(n66313), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n51606), .O(n27990)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_25  (.CI(n51606), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n51607));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_24_lut  (.I0(n66312), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n51605), .O(n27992)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_24  (.CI(n51605), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n51606));
    SB_LUT4 \FRAME_MATCHER.i_1943_add_4_23_lut  (.I0(n66310), .I1(n70121), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n51604), .O(n27994)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1943_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1943_add_4_23  (.CI(n51604), .I0(n70121), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n51605));
    SB_LUT4 select_780_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1375 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[12] [3]), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1375.LUT_INIT = 16'ha088;
    SB_LUT4 select_780_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i50817_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66347));   // verilog/coms.v(158[12:15])
    defparam i50817_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_780_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_304_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5535));
    defparam equal_304_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 select_780_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1376 (.I0(n23929), .I1(n23933), .I2(\data_in_frame[8]_c [1]), 
            .I3(\data_in_frame[8]_c [7]), .O(n58520));   // verilog/coms.v(88[17:28])
    defparam i1_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51032_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66350));   // verilog/coms.v(158[12:15])
    defparam i51032_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_780_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1377 (.I0(n23929), .I1(n23933), .I2(\data_in_frame[10] [0]), 
            .I3(n58128), .O(n52885));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(\data_in_frame[14] [3]), .I1(n25130), 
            .I2(n26379), .I3(GND_net), .O(n25218));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(\data_in_frame[14] [3]), .I1(n25130), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n58093));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1380 (.I0(n25862), .I1(n58090), .I2(n58598), 
            .I3(n52731), .O(n53066));
    defparam i1_3_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i28376_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n42296));
    defparam i28376_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i5_3_lut_4_lut (.I0(n25862), .I1(n58090), .I2(n53743), .I3(n10_adj_5582), 
            .O(n25130));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1381 (.I0(\data_in_frame[9] [3]), .I1(n25716), 
            .I2(n58068), .I3(n58154), .O(n26463));
    defparam i2_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(tx_active), .I1(n97), .I2(r_SM_Main_2__N_3545[0]), 
            .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n25514));
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'hfb00;
    SB_LUT4 i2_3_lut_4_lut_adj_1383 (.I0(\data_in_frame[9] [3]), .I1(n25716), 
            .I2(n26274), .I3(n58128), .O(n58598));
    defparam i2_3_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i51065_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66354));   // verilog/coms.v(158[12:15])
    defparam i51065_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1384 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(n52776), .I3(n58657), .O(n52751));
    defparam i2_3_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1385 (.I0(tx_active), .I1(n97), .I2(r_SM_Main_2__N_3545[0]), 
            .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n22691));
    defparam i1_2_lut_4_lut_adj_1385.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_4_lut_adj_1386 (.I0(n26493), .I1(n58310), .I2(\data_in_frame[13] [0]), 
            .I3(n58316), .O(n4_adj_5583));
    defparam i1_2_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1387 (.I0(n26493), .I1(n58310), .I2(\data_in_frame[13] [0]), 
            .I3(n53833), .O(n58015));
    defparam i1_2_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1388 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[19] [0]), 
            .I2(n58582), .I3(\data_out_frame[18] [6]), .O(n6_adj_5584));
    defparam i1_2_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i50895_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66281));   // verilog/coms.v(158[12:15])
    defparam i50895_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1389 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[18] [4]), 
            .I2(n53853), .I3(GND_net), .O(n6_adj_5585));
    defparam i1_2_lut_3_lut_adj_1389.LUT_INIT = 16'h6969;
    SB_LUT4 i51062_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66355));   // verilog/coms.v(158[12:15])
    defparam i51062_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1390 (.I0(\data_out_frame[16] [0]), .I1(n52801), 
            .I2(\data_out_frame[15] [5]), .I3(n26265), .O(n53848));
    defparam i1_2_lut_3_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[11][2] ), .O(n57277));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i51063_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66356));   // verilog/coms.v(158[12:15])
    defparam i51063_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_3_lut_4_lut_adj_1391 (.I0(\data_in_frame[11] [6]), .I1(n23929), 
            .I2(n26466), .I3(n25974), .O(n20_adj_5586));
    defparam i7_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1392 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12]_c [7]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n63190));
    defparam i1_2_lut_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1393 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1951), .I3(n1954), .O(n25520));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1393.LUT_INIT = 16'h4000;
    SB_LUT4 i3_3_lut_4_lut_adj_1394 (.I0(\data_out_frame[23] [0]), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[25] [3]), .I3(n53763), .O(n8_adj_5587));
    defparam i3_3_lut_4_lut_adj_1394.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1395 (.I0(\data_out_frame[14] [4]), .I1(n58313), 
            .I2(n58275), .I3(\data_out_frame[16] [5]), .O(n58202));
    defparam i1_2_lut_3_lut_4_lut_adj_1395.LUT_INIT = 16'h9669;
    SB_LUT4 select_780_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut_3_lut_4_lut (.I0(\data_out_frame[14] [4]), .I1(n58313), 
            .I2(n58275), .I3(\data_out_frame[18] [5]), .O(n12_adj_5588));
    defparam i4_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_780_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14798_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28829));   // verilog/coms.v(130[12] 305[6])
    defparam i14798_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_780_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1396 (.I0(n1951), .I1(n4452), .I2(n1954), 
            .I3(n1957), .O(n60097));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1396.LUT_INIT = 16'h2000;
    SB_LUT4 i2_2_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(\FRAME_MATCHER.i_31__N_2512 ), 
            .O(n6_adj_5589));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1951), .I1(n4452), .I2(n63421), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n60837));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 select_780_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14796_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28827));   // verilog/coms.v(130[12] 305[6])
    defparam i14796_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1397 (.I0(reset), .I1(n57993), .I2(GND_net), 
            .I3(GND_net), .O(n57986));
    defparam i1_2_lut_adj_1397.LUT_INIT = 16'heeee;
    SB_LUT4 select_780_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1398 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n57983), .O(n28358));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1398.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1399 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n57993), .O(n28322));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1399.LUT_INIT = 16'hfff7;
    SB_LUT4 i53557_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[7]_c [7]), 
            .I2(n58897), .I3(GND_net), .O(n57319));   // verilog/coms.v(94[13:20])
    defparam i53557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_780_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(n8_adj_8), .I1(n57974), .I2(GND_net), 
            .I3(GND_net), .O(n28338));
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'heeee;
    SB_LUT4 select_780_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(\data_in_frame[12]_c [1]), .I1(\data_in_frame[11] [7]), 
            .I2(n53066), .I3(\data_in_frame[9][7] ), .O(n58012));
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i15417_3_lut (.I0(\data_in_frame[0]_c [7]), .I1(rx_data[7]), 
            .I2(n58008), .I3(GND_net), .O(n29448));   // verilog/coms.v(130[12] 305[6])
    defparam i15417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 select_780_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(\data_in_frame[9] [3]), .I1(n53348), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n53743));
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'h9696;
    SB_LUT4 i15414_3_lut (.I0(\data_in_frame[0]_c [6]), .I1(rx_data[6]), 
            .I2(n58008), .I3(GND_net), .O(n29445));   // verilog/coms.v(130[12] 305[6])
    defparam i15414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 select_780_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_in_frame[10] [4]), .I1(n4_adj_5342), 
            .I2(n3_adj_5376), .I3(GND_net), .O(n26042));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n58666));
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[12]_c [3]), 
            .I2(n26853), .I3(GND_net), .O(n6_adj_5590));
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\control_mode[0] ), .I1(n37407), 
            .I2(\control_mode[1] ), .I3(GND_net), .O(n15_adj_10));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_4_lut_adj_1407 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[15] [5]), 
            .I2(n58419), .I3(\data_in_frame[17] [7]), .O(n58621));
    defparam i1_2_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1408 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n53720), .I3(GND_net), .O(n53921));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1408.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1409 (.I0(\data_in_frame[17]_c [1]), .I1(n53137), 
            .I2(\data_in_frame[19] [3]), .I3(n25141), .O(n61005));
    defparam i2_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1410 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [0]), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1410.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1411 (.I0(\data_in_frame[13] [5]), .I1(n25961), 
            .I2(n36_adj_5592), .I3(GND_net), .O(n25996));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1412 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(Kp_23__N_1301), .I3(n58561), .O(n53737));
    defparam i1_2_lut_4_lut_adj_1412.LUT_INIT = 16'h9669;
    SB_LUT4 select_780_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n58272));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i53558_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[7]_c [6]), 
            .I2(n58897), .I3(GND_net), .O(n57325));   // verilog/coms.v(94[13:20])
    defparam i53558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51684_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66361));   // verilog/coms.v(158[12:15])
    defparam i51684_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1414 (.I0(n53137), .I1(n53706), .I2(\data_in_frame[19]_c [4]), 
            .I3(n58425), .O(n58675));
    defparam i1_2_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1415 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1415.LUT_INIT = 16'ha088;
    SB_LUT4 equal_308_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_11));   // verilog/coms.v(157[7:23])
    defparam equal_308_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_3_lut_4_lut_adj_1416 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n26463), .I3(\data_in_frame[14] [0]), .O(n26330));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1417 (.I0(\data_in_frame[16] [5]), .I1(n25218), 
            .I2(\data_in_frame[18]_c [6]), .I3(\data_in_frame[20] [7]), 
            .O(n58663));
    defparam i2_3_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i25_3_lut (.I0(n28358), .I1(rx_data[5]), .I2(\data_in_frame[19]_c [5]), 
            .I3(GND_net), .O(n17_adj_5532));   // verilog/coms.v(94[13:20])
    defparam i25_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i51285_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66282));   // verilog/coms.v(158[12:15])
    defparam i51285_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut_adj_1418 (.I0(\data_in_frame[16] [5]), .I1(n25218), 
            .I2(\data_in_frame[18][0] ), .I3(n58448), .O(n63108));
    defparam i1_3_lut_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1419 (.I0(n52807), .I1(n58672), .I2(n26087), 
            .I3(GND_net), .O(n58211));
    defparam i1_2_lut_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(\data_in_frame[16] [4]), .I1(n26379), 
            .I2(\data_in_frame[16] [5]), .I3(n53776), .O(n52407));
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1421 (.I0(\data_in_frame[18][3] ), .I1(n60610), 
            .I2(\data_in_frame[20] [6]), .I3(\data_in_frame[20] [5]), .O(n58585));
    defparam i2_3_lut_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i51683_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n66360));   // verilog/uart_tx.v(32[16:25])
    defparam i51683_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1422 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n57912));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1422.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(\control_mode[0] ), .I1(n37407), 
            .I2(\control_mode[1] ), .I3(GND_net), .O(n15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n63769), .I3(n63767), .O(n7_adj_5594));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n63757), .I3(n63755), .O(n7_adj_5595));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n63751), .I3(n63749), .O(n7_adj_5596));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_3_lut_4_lut_adj_1424 (.I0(\data_in_frame[18][3] ), .I1(n60610), 
            .I2(\data_in_frame[20][4] ), .I3(\data_in_frame[20][3] ), .O(n5_adj_5401));
    defparam i1_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1425 (.I0(n26466), .I1(n58154), .I2(\data_in_frame[11] [4]), 
            .I3(\data_in_frame[9] [3]), .O(n36_adj_5592));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n40523), .I1(n3472), .I2(rx_data_ready), 
            .I3(\FRAME_MATCHER.rx_data_ready_prev ), .O(n40525));   // verilog/coms.v(156[9:50])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1426 (.I0(n26466), .I1(n26306), .I2(\data_in_frame[9] [2]), 
            .I3(n58766), .O(n6_adj_5597));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(\data_in_frame[21][2] ), .I1(\data_in_frame[21][1] ), 
            .I2(n58455), .I3(GND_net), .O(n6_adj_5598));
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1428 (.I0(\data_in_frame[21][2] ), .I1(\data_in_frame[21][1] ), 
            .I2(\data_in_frame[16] [3]), .I3(n58392), .O(n58400));
    defparam i2_3_lut_4_lut_adj_1428.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1429 (.I0(n53933), .I1(n53824), .I2(\data_in_frame[17][5] ), 
            .I3(n60893), .O(n58403));
    defparam i1_2_lut_4_lut_adj_1429.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n63739), .I3(n63737), .O(n7_adj_5599));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54539 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n70291));
    defparam byte_transmit_counter_0__bdd_4_lut_54539.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1430 (.I0(n53933), .I1(n53824), .I2(\data_in_frame[17][5] ), 
            .I3(n52407), .O(n58448));
    defparam i1_2_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n63778), .I3(n63776), .O(n7_adj_5339));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i3_3_lut_4_lut_adj_1431 (.I0(n40523), .I1(n3472), .I2(reset), 
            .I3(n161), .O(n57983));   // verilog/coms.v(156[9:50])
    defparam i3_3_lut_4_lut_adj_1431.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_4_lut_4_lut (.I0(reset), .I1(n28338), .I2(\data_in_frame[1]_c [1]), 
            .I3(rx_data[1]), .O(n57379));   // verilog/coms.v(94[13:20])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1432 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25514), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n63421));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1432.LUT_INIT = 16'hfff4;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1433 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12]_c [7]), 
            .I2(\data_in_frame[12]_c [4]), .I3(\data_in_frame[10] [5]), 
            .O(n63258));
    defparam i1_2_lut_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1057_i2_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n4764[1]));
    defparam mux_1057_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i3_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3][2] ), .I3(\data_in_frame[19] [2]), .O(n4764[2]));
    defparam mux_1057_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i4_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n4764[3]));
    defparam mux_1057_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i28_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), .I1(byte_transmit_counter[1]), 
            .I2(n10_adj_5550), .I3(n4_adj_5551), .O(n57571));   // verilog/coms.v(109[34:55])
    defparam i28_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1434 (.I0(\data_in_frame[11] [6]), .I1(n26663), 
            .I2(n58157), .I3(\data_in_frame[11] [4]), .O(n58068));
    defparam i1_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i21002_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [4]), 
            .I3(\data_in_frame[19]_c [4]), .O(n4764[4]));
    defparam i21002_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i19_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), .I2(n17), 
            .I3(encoder0_position_scaled[0]), .O(n18_adj_12));   // verilog/coms.v(130[12] 305[6])
    defparam i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_1057_i6_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3][5] ), .I3(\data_in_frame[19]_c [5]), .O(n4764[5]));
    defparam mux_1057_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i7_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3]_c [6]), .I3(\data_in_frame[19] [6]), .O(n4764[6]));
    defparam mux_1057_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_243_i2_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[1] ), .I3(encoder0_position_scaled[1]), 
            .O(\motor_state[1] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i20889_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][7] ), 
            .I3(\data_in_frame[19] [7]), .O(n4764[7]));
    defparam i20889_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i9_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][0] ), .I3(\data_in_frame[18][0] ), .O(n4764[8]));
    defparam mux_1057_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1435 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(\data_in_frame[16] [0]), .I3(\data_in_frame[16] [1]), .O(n6_adj_5602));
    defparam i1_2_lut_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1057_i10_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][1] ), .I3(\data_in_frame[18][1] ), .O(n4764[9]));
    defparam mux_1057_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i21388_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [2]), 
            .I3(\data_in_frame[18]_c [2]), .O(n4764[10]));
    defparam i21388_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_243_i3_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[2] ), .I3(encoder0_position_scaled[2]), 
            .O(\motor_state[2] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_1057_i12_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][3] ), .I3(\data_in_frame[18][3] ), .O(n4764[11]));
    defparam mux_1057_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i21236_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [4]), 
            .I3(\data_in_frame[18][4] ), .O(n4764[12]));
    defparam i21236_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i14_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[2][5] ), .I3(\data_in_frame[18] [5]), .O(n4764[13]));
    defparam mux_1057_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_243_i4_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[3] ), .I3(encoder0_position_scaled[3]), 
            .O(\motor_state[3] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i21205_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[18]_c [6]), .O(n4764[14]));
    defparam i21205_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_243_i5_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[4] ), .I3(encoder0_position_scaled[4]), 
            .O(\motor_state[4] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i21204_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[18][7] ), .O(n4764[15]));
    defparam i21204_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i17_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1]_c [0]), .I3(\data_in_frame[17] [0]), .O(n4764[16]));
    defparam mux_1057_i17_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_243_i6_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[5] ), .I3(encoder0_position_scaled[5]), 
            .O(\motor_state[5] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i21469_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[1]_c [1]), 
            .I3(\data_in_frame[17]_c [1]), .O(n4764[17]));
    defparam i21469_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i22_3_lut (.I0(n28358), .I1(rx_data[4]), .I2(\data_in_frame[19]_c [4]), 
            .I3(GND_net), .O(n14_adj_5531));   // verilog/coms.v(94[13:20])
    defparam i22_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_243_i7_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[6] ), .I3(encoder0_position_scaled[6]), 
            .O(\motor_state[6] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i21440_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[1][2] ), 
            .I3(\data_in_frame[17]_c [2]), .O(n4764[18]));
    defparam i21440_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i20_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1]_c [3]), .I3(\data_in_frame[17][3] ), .O(n4764[19]));
    defparam mux_1057_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1436 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n57913));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1436.LUT_INIT = 16'h5100;
    SB_LUT4 mux_1057_i21_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1]_c [4]), .I3(\data_in_frame[17][4] ), .O(n4764[20]));
    defparam mux_1057_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i16292_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30323));   // verilog/coms.v(130[12] 305[6])
    defparam i16292_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1057_i22_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17][5] ), .O(n4764[21]));
    defparam mux_1057_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_243_i8_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[7] ), .I3(encoder0_position_scaled[7]), 
            .O(\motor_state[7] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_1057_i23_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][6] ), .I3(\data_in_frame[17][6] ), .O(n4764[22]));
    defparam mux_1057_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1057_i24_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[1][7] ), .I3(\data_in_frame[17] [7]), .O(n4764[23]));
    defparam mux_1057_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i15388_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [0]), 
            .I3(deadband[0]), .O(n29419));
    defparam i15388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16215_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8]_c [7]), 
            .I3(PWMLimit[23]), .O(n30246));
    defparam i16215_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16322_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30353));   // verilog/coms.v(130[12] 305[6])
    defparam i16322_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16321_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30352));   // verilog/coms.v(130[12] 305[6])
    defparam i16321_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16320_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30351));   // verilog/coms.v(130[12] 305[6])
    defparam i16320_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16244_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8][6] ), 
            .I3(PWMLimit[22]), .O(n30275));
    defparam i16244_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16259_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8]_c [5]), 
            .I3(PWMLimit[21]), .O(n30290));
    defparam i16259_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16264_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n30295));
    defparam i16264_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23377_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8][3] ), 
            .I3(PWMLimit[19]), .O(n30315));
    defparam i23377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16291_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n30322));
    defparam i16291_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i22406_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8]_c [1]), 
            .I3(PWMLimit[17]), .O(n36387));
    defparam i22406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_3_lut_adj_1437 (.I0(\data_in_frame[18]_c [6]), .I1(rx_data[6]), 
            .I2(n28361), .I3(GND_net), .O(n57129));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1437.LUT_INIT = 16'hcaca;
    SB_LUT4 i16377_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[8]_c [0]), 
            .I3(PWMLimit[16]), .O(n30408));
    defparam i16377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15581_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n29612));
    defparam i15581_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15582_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][0] ), 
            .I3(\Kp[0] ), .O(n29613));
    defparam i15582_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15583_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n29614));
    defparam i15583_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i25_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), .I2(n12_adj_5603), 
            .I3(encoder0_position_scaled[8]), .O(n10));   // verilog/coms.v(130[12] 305[6])
    defparam i25_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i10_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[9] ), .I3(encoder0_position_scaled[9]), 
            .O(\motor_state[9] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15587_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n29618));
    defparam i15587_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_243_i11_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[10] ), .I3(encoder0_position_scaled[10]), 
            .O(\motor_state[10] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15650_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n29681));
    defparam i15650_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15651_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n29682));
    defparam i15651_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16319_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30350));   // verilog/coms.v(130[12] 305[6])
    defparam i16319_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15652_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n29683));
    defparam i15652_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15653_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n29684));
    defparam i15653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i50833_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66284));   // verilog/coms.v(158[12:15])
    defparam i50833_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_1438 (.I0(n66360), .I1(n59012), .I2(r_Bit_Index[0]), 
            .I3(n59553), .O(n53963));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut_adj_1438.LUT_INIT = 16'h303a;
    SB_LUT4 i15654_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n29685));
    defparam i15654_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15655_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n29686));
    defparam i15655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15656_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n29687));
    defparam i15656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i50906_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66286));   // verilog/coms.v(158[12:15])
    defparam i50906_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1439 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n57914));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1439.LUT_INIT = 16'h5100;
    SB_LUT4 i1_3_lut_adj_1440 (.I0(n58678), .I1(n58435), .I2(n60610), 
            .I3(GND_net), .O(n58336));
    defparam i1_3_lut_adj_1440.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1441 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[13] [6]), .I3(\data_in_frame[15] [7]), .O(n63010));
    defparam i1_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i15657_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n29688));
    defparam i15657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1442 (.I0(n63010), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[12]_c [5]), .I3(\data_in_frame[18][1] ), 
            .O(n63012));
    defparam i1_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i15658_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n29689));
    defparam i15658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_243_i12_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[11] ), .I3(encoder0_position_scaled[11]), 
            .O(\motor_state[11] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1443 (.I0(n58220), .I1(n25908), .I2(n26414), 
            .I3(n58490), .O(n63020));
    defparam i1_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i15659_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n29690));
    defparam i15659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1444 (.I0(Kp_23__N_1067), .I1(n63020), .I2(n58648), 
            .I3(n63012), .O(n63024));
    defparam i1_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1445 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n52778), .I3(n6_adj_5602), .O(n60724));
    defparam i4_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i15660_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n29691));
    defparam i15660_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1446 (.I0(n58624), .I1(n26330), .I2(n52778), 
            .I3(n63024), .O(n63030));
    defparam i1_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1447 (.I0(\data_in_frame[12]_c [7]), .I1(n63030), 
            .I2(n60724), .I3(\data_in_frame[15] [4]), .O(n63032));
    defparam i1_4_lut_adj_1447.LUT_INIT = 16'h9669;
    SB_LUT4 i15661_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n29692));
    defparam i15661_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1448 (.I0(n25218), .I1(n52737), .I2(n53921), 
            .I3(n63032), .O(n63038));
    defparam i1_4_lut_adj_1448.LUT_INIT = 16'h9669;
    SB_LUT4 i16318_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30349));   // verilog/coms.v(130[12] 305[6])
    defparam i16318_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1449 (.I0(n53737), .I1(n58432), .I2(n53933), 
            .I3(n63038), .O(n63044));
    defparam i1_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1450 (.I0(n58096), .I1(n53750), .I2(n58392), 
            .I3(n63044), .O(n58678));
    defparam i1_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i16317_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30348));   // verilog/coms.v(130[12] 305[6])
    defparam i16317_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15662_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n29693));
    defparam i15662_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16316_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30347));   // verilog/coms.v(130[12] 305[6])
    defparam i16316_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1451 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n57915));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1451.LUT_INIT = 16'h5100;
    SB_LUT4 i15663_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n29694));
    defparam i15663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1452 (.I0(n52751), .I1(n63108), .I2(n52410), 
            .I3(n58678), .O(n58435));
    defparam i1_4_lut_adj_1452.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1453 (.I0(n52807), .I1(n58672), .I2(GND_net), 
            .I3(GND_net), .O(n23886));
    defparam i1_2_lut_adj_1453.LUT_INIT = 16'h6666;
    SB_LUT4 i16315_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30346));   // verilog/coms.v(130[12] 305[6])
    defparam i16315_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1454 (.I0(\data_in_frame[20][3] ), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[20][4] ), .I3(\data_in_frame[20] [2]), .O(n63132));
    defparam i1_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i16314_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30345));   // verilog/coms.v(130[12] 305[6])
    defparam i16314_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_adj_1455 (.I0(n58179), .I1(n58339), .I2(n63132), 
            .I3(GND_net), .O(n63136));
    defparam i1_3_lut_adj_1455.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1456 (.I0(n23886), .I1(n58435), .I2(n58585), 
            .I3(n63136), .O(n58745));
    defparam i1_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i15664_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[9][7] ), 
            .I3(PWMLimit[15]), .O(n29695));
    defparam i15664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1457 (.I0(n53737), .I1(n25996), .I2(\data_in_frame[18][3] ), 
            .I3(\data_in_frame[19] [7]), .O(n63118));
    defparam i1_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1458 (.I0(n61005), .I1(n52407), .I2(n63118), 
            .I3(n58663), .O(n63124));
    defparam i1_4_lut_adj_1458.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1459 (.I0(n58403), .I1(n58745), .I2(n58675), 
            .I3(n63124), .O(n53829));
    defparam i1_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 mux_243_i13_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[12] ), .I3(encoder0_position_scaled[12]), 
            .O(\motor_state[12] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16313_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30344));   // verilog/coms.v(130[12] 305[6])
    defparam i16313_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1460 (.I0(n52853), .I1(\data_in_frame[21][5] ), 
            .I2(n58458), .I3(n6_adj_5598), .O(n53861));
    defparam i4_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i16312_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30343));   // verilog/coms.v(130[12] 305[6])
    defparam i16312_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15703_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n29734));
    defparam i15703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1461 (.I0(\data_in_frame[20][1] ), .I1(n58419), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[20][0] ), .O(n58179));
    defparam i3_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(\data_in_frame[21][7] ), .I1(\data_in_frame[21] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58458));
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n57901));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_adj_1463 (.I0(n58093), .I1(n58391), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n52410));
    defparam i2_3_lut_adj_1463.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1464 (.I0(\data_in_frame[18][3] ), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58220));
    defparam i1_2_lut_adj_1464.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1465 (.I0(n61005), .I1(\data_in_frame[21][5] ), 
            .I2(\data_in_frame[21] [6]), .I3(GND_net), .O(n58208));
    defparam i2_3_lut_adj_1465.LUT_INIT = 16'h6969;
    SB_LUT4 i15704_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n29735));
    defparam i15704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1466 (.I0(n60893), .I1(\data_in_frame[19]_c [5]), 
            .I2(n53706), .I3(GND_net), .O(n52853));
    defparam i2_3_lut_adj_1466.LUT_INIT = 16'h6969;
    SB_LUT4 mux_243_i14_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[13] ), .I3(encoder0_position_scaled[13]), 
            .O(\motor_state[13] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15705_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n29736));
    defparam i15705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16311_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30342));   // verilog/coms.v(130[12] 305[6])
    defparam i16311_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1467 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n40523));
    defparam i2_3_lut_adj_1467.LUT_INIT = 16'h1010;
    SB_LUT4 i16310_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30341));   // verilog/coms.v(130[12] 305[6])
    defparam i16310_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16309_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30340));   // verilog/coms.v(130[12] 305[6])
    defparam i16309_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1468 (.I0(n53137), .I1(n53706), .I2(\data_in_frame[19]_c [4]), 
            .I3(GND_net), .O(n52879));
    defparam i2_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 mux_243_i15_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[14] ), .I3(encoder0_position_scaled[14]), 
            .O(\motor_state[14] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 equal_300_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_13));   // verilog/coms.v(157[7:23])
    defparam equal_300_i7_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_in_frame[21][4] ), .I1(n58675), 
            .I2(GND_net), .I3(GND_net), .O(n58330));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1470 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[20] [6]), 
            .I2(\data_in_frame[16] [2]), .I3(GND_net), .O(n14_adj_5606));
    defparam i5_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1471 (.I0(n58714), .I1(\data_in_frame[21][0] ), 
            .I2(n58392), .I3(n58657), .O(n15_adj_5607));
    defparam i6_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1472 (.I0(n15_adj_5607), .I1(\data_in_frame[18] [5]), 
            .I2(n14_adj_5606), .I3(\data_in_frame[18][4] ), .O(n26087));
    defparam i8_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i15706_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n29737));
    defparam i15706_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16308_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30339));   // verilog/coms.v(130[12] 305[6])
    defparam i16308_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15707_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n29738));
    defparam i15707_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1473 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[12]_c [6]), .I3(GND_net), .O(n58648));
    defparam i2_3_lut_adj_1473.LUT_INIT = 16'h9696;
    SB_LUT4 i15708_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n29739));
    defparam i15708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_adj_1474 (.I0(n58648), .I1(\data_in_frame[13] [2]), 
            .I2(\data_in_frame[12]_c [7]), .I3(GND_net), .O(n63206));
    defparam i1_3_lut_adj_1474.LUT_INIT = 16'h9696;
    SB_LUT4 i15709_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n29740));
    defparam i15709_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16307_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30338));   // verilog/coms.v(130[12] 305[6])
    defparam i16307_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_243_i22_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[21] ), .I3(encoder0_position_scaled[21]), 
            .O(\motor_state[21] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16306_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30337));   // verilog/coms.v(130[12] 305[6])
    defparam i16306_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1475 (.I0(n26042), .I1(n58378), .I2(n25862), 
            .I3(n63206), .O(n53795));
    defparam i1_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1476 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(n58627), .I3(\data_in_frame[13] [1]), .O(n53933));
    defparam i1_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1477 (.I0(\data_in_frame[15] [3]), .I1(n53795), 
            .I2(\data_in_frame[17][4] ), .I3(GND_net), .O(n60893));
    defparam i1_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1478 (.I0(\data_in_frame[18]_c [2]), .I1(n28304), 
            .I2(n28361), .I3(rx_data[2]), .O(n57109));
    defparam i12_4_lut_adj_1478.LUT_INIT = 16'h3a0a;
    SB_LUT4 i16305_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30336));   // verilog/coms.v(130[12] 305[6])
    defparam i16305_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15710_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n29741));
    defparam i15710_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1479 (.I0(n58253), .I1(n10_adj_5269), .I2(\data_out_frame[20] [0]), 
            .I3(n58381), .O(n4));
    defparam i1_2_lut_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i15711_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n29742));
    defparam i15711_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1480 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[17][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n63224));
    defparam i1_2_lut_adj_1480.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1481 (.I0(n58451), .I1(n53795), .I2(n53921), 
            .I3(n63224), .O(n58681));
    defparam i1_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i15712_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n29743));
    defparam i15712_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_243_i18_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[17] ), .I3(encoder0_position_scaled[17]), 
            .O(\motor_state[17] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_3_lut_adj_1482 (.I0(n58681), .I1(n53737), .I2(n25996), 
            .I3(GND_net), .O(n53706));
    defparam i1_3_lut_adj_1482.LUT_INIT = 16'h6969;
    SB_LUT4 i16304_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30335));   // verilog/coms.v(130[12] 305[6])
    defparam i16304_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1483 (.I0(n53824), .I1(\data_in_frame[17][6] ), 
            .I2(n53737), .I3(GND_net), .O(n58612));
    defparam i2_3_lut_adj_1483.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(n58403), .I1(n53706), .I2(GND_net), 
            .I3(GND_net), .O(n53750));
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h9999;
    SB_LUT4 i15713_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n29744));
    defparam i15713_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15714_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n29745));
    defparam i15714_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1485 (.I0(\data_in_frame[21][7] ), .I1(\data_in_frame[19]_c [5]), 
            .I2(\data_in_frame[19] [7]), .I3(GND_net), .O(n58269));
    defparam i2_3_lut_adj_1485.LUT_INIT = 16'h9696;
    SB_LUT4 i15715_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n29746));
    defparam i15715_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n63146));
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'h6666;
    SB_LUT4 i16303_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30334));   // verilog/coms.v(130[12] 305[6])
    defparam i16303_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1487 (.I0(Kp_23__N_974), .I1(n53323), .I2(n63146), 
            .I3(\data_in_frame[8][6] ), .O(n58378));
    defparam i1_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i16302_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30333));   // verilog/coms.v(130[12] 305[6])
    defparam i16302_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16301_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30332));   // verilog/coms.v(130[12] 305[6])
    defparam i16301_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1488 (.I0(n25947), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[13] [3]), .O(n62968));
    defparam i1_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i16300_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30331));   // verilog/coms.v(130[12] 305[6])
    defparam i16300_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_780_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1489 (.I0(\data_in_frame[15] [4]), .I1(n58378), 
            .I2(n58561), .I3(n62968), .O(n53824));
    defparam i1_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(\data_in_frame[17][6] ), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n63230));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 i16299_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30330));   // verilog/coms.v(130[12] 305[6])
    defparam i16299_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_780_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1491 (.I0(n25996), .I1(n53824), .I2(n63230), 
            .I3(\data_in_frame[17] [7]), .O(n58096));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1491.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_in_frame[20] [2]), .I1(Kp_23__N_1301), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5608));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1493 (.I0(\data_in_frame[18][0] ), .I1(\data_in_frame[13] [4]), 
            .I2(n58096), .I3(n6_adj_5608), .O(n58323));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i15716_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n29747));
    defparam i15716_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(n25961), .I1(n36_adj_5592), .I2(GND_net), 
            .I3(GND_net), .O(n58176));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 mux_243_i20_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[19] ), .I3(encoder0_position_scaled[19]), 
            .O(\motor_state[19] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1495 (.I0(n25862), .I1(n53323), .I2(n4_adj_5342), 
            .I3(n63190), .O(n58627));
    defparam i1_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i16298_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30329));   // verilog/coms.v(130[12] 305[6])
    defparam i16298_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(Kp_23__N_1301), .I1(n58561), .I2(GND_net), 
            .I3(GND_net), .O(n52723));
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h9999;
    SB_LUT4 i20894_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n29748));
    defparam i20894_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_adj_1497 (.I0(\data_in_frame[14] [7]), .I1(n36_adj_5592), 
            .I2(n58015), .I3(GND_net), .O(n58451));
    defparam i1_3_lut_adj_1497.LUT_INIT = 16'h6969;
    SB_LUT4 i16297_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30328));   // verilog/coms.v(130[12] 305[6])
    defparam i16297_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15718_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n29749));
    defparam i15718_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1498 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58490));
    defparam i1_2_lut_adj_1498.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1499 (.I0(n58034), .I1(n26042), .I2(\data_in_frame[17]_c [2]), 
            .I3(n58490), .O(n16_adj_5609));
    defparam i6_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i15720_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n29751));
    defparam i15720_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut_adj_1500 (.I0(n53770), .I1(n58627), .I2(n58176), 
            .I3(n53833), .O(n17_adj_5610));
    defparam i7_4_lut_adj_1500.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1501 (.I0(n17_adj_5610), .I1(n58451), .I2(n16_adj_5609), 
            .I3(n52723), .O(n53137));
    defparam i9_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\data_in_frame[17]_c [1]), .I1(n53137), 
            .I2(GND_net), .I3(GND_net), .O(n58432));
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h6666;
    SB_LUT4 i15721_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][5] ), 
            .I3(\Kp[13] ), .O(n29752));
    defparam i15721_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15722_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n29753));
    defparam i15722_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1503 (.I0(\data_in_frame[21][4] ), .I1(n52807), 
            .I2(\data_in_frame[21][3] ), .I3(GND_net), .O(n58455));
    defparam i2_3_lut_adj_1503.LUT_INIT = 16'h9696;
    SB_LUT4 i16296_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30327));   // verilog/coms.v(130[12] 305[6])
    defparam i16296_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1504 (.I0(\data_in_frame[13] [7]), .I1(n58615), 
            .I2(n53728), .I3(\data_in_frame[11] [5]), .O(n58391));
    defparam i3_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(n26379), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58114));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1506 (.I0(\data_in_frame[14] [3]), .I1(n58429), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5611));
    defparam i1_2_lut_adj_1506.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1507 (.I0(n52778), .I1(n25130), .I2(n58114), 
            .I3(n6_adj_5611), .O(n52737));
    defparam i4_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i16295_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30326));   // verilog/coms.v(130[12] 305[6])
    defparam i16295_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_243_i21_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[20] ), .I3(encoder0_position_scaled[20]), 
            .O(\motor_state[20] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15723_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][3] ), 
            .I3(\Kp[11] ), .O(n29754));
    defparam i15723_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i21379_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n29755));
    defparam i21379_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(n53776), .I1(n58391), .I2(GND_net), 
            .I3(GND_net), .O(n58392));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h6666;
    SB_LUT4 i47626_3_lut_4_lut (.I0(n26343), .I1(\data_in_frame[0][5] ), 
            .I2(\data_in_frame[0]_c [6]), .I3(\data_in_frame[2] [7]), .O(n63337));
    defparam i47626_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i2_3_lut_adj_1509 (.I0(\data_in_frame[18][7] ), .I1(n52737), 
            .I2(\data_in_frame[19] [1]), .I3(GND_net), .O(n52807));
    defparam i2_3_lut_adj_1509.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1510 (.I0(n25103), .I1(n53066), .I2(n52731), 
            .I3(GND_net), .O(n59945));
    defparam i1_3_lut_adj_1510.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1511 (.I0(n7_adj_5377), .I1(n59945), .I2(n58598), 
            .I3(n58148), .O(n53323));
    defparam i1_4_lut_adj_1511.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1512 (.I0(n53323), .I1(n26463), .I2(n60258), 
            .I3(\data_in_frame[16] [0]), .O(n58419));
    defparam i3_4_lut_adj_1512.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1513 (.I0(\data_in_frame[15] [5]), .I1(n58419), 
            .I2(\data_in_frame[17] [7]), .I3(GND_net), .O(n25115));
    defparam i2_3_lut_adj_1513.LUT_INIT = 16'h9696;
    SB_LUT4 i16294_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30325));   // verilog/coms.v(130[12] 305[6])
    defparam i16294_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1514 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2][5] ), 
            .I2(\data_in_frame[0][4] ), .I3(GND_net), .O(n25806));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1514.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1515 (.I0(\data_in_frame[14] [1]), .I1(n58607), 
            .I2(n25771), .I3(n6_adj_5597), .O(n58615));
    defparam i4_4_lut_adj_1515.LUT_INIT = 16'h9669;
    SB_LUT4 i16293_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30324));   // verilog/coms.v(130[12] 305[6])
    defparam i16293_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_780_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_adj_1516 (.I0(\data_in_frame[16] [1]), .I1(n25961), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n14_adj_5612));
    defparam i5_3_lut_adj_1516.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1517 (.I0(n58615), .I1(\data_in_frame[16] [2]), 
            .I2(n53743), .I3(n58272), .O(n15_adj_5613));
    defparam i6_4_lut_adj_1517.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1518 (.I0(n15_adj_5613), .I1(n26294), .I2(n14_adj_5612), 
            .I3(n53728), .O(n60610));
    defparam i8_4_lut_adj_1518.LUT_INIT = 16'h9669;
    SB_LUT4 i15598_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29629));   // verilog/coms.v(130[12] 305[6])
    defparam i15598_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15725_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][1] ), 
            .I3(\Kp[9] ), .O(n29756));
    defparam i15725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1519 (.I0(\data_out_frame[20] [3]), .I1(n53723), 
            .I2(n58346), .I3(\data_out_frame[24] [7]), .O(n58742));
    defparam i1_2_lut_3_lut_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i15_2_lut (.I0(\data_in_frame[18][4] ), .I1(\data_in_frame[18]_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26414));   // verilog/coms.v(99[12:25])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15726_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[2][0] ), 
            .I3(\Kp[8] ), .O(n29757));
    defparam i15726_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1520 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(n58163), .I3(\data_in_frame[12]_c [6]), .O(n10_adj_5614));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1521 (.I0(n25947), .I1(n10_adj_5614), .I2(n4_adj_5342), 
            .I3(GND_net), .O(n58034));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_adj_1521.LUT_INIT = 16'h9696;
    SB_LUT4 mux_243_i23_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[22] ), .I3(encoder0_position_scaled[22]), 
            .O(\motor_state[22] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i24_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[23] ), .I3(encoder0_position_scaled[23]), 
            .O(\motor_state[23] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15727_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][7] ), 
            .I3(\Kp[7] ), .O(n29758));
    defparam i15727_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i26778_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), .I2(n5), 
            .I3(encoder0_position_scaled[16]), .O(n7_adj_14));   // verilog/coms.v(130[12] 305[6])
    defparam i26778_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i20888_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [6]), 
            .I3(\Kp[6] ), .O(n29759));
    defparam i20888_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1522 (.I0(\data_in_frame[12]_c [4]), .I1(n59815), 
            .I2(GND_net), .I3(GND_net), .O(n58624));
    defparam i1_2_lut_adj_1522.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1523 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5616));
    defparam i1_2_lut_adj_1523.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1524 (.I0(\data_in_frame[17] [0]), .I1(n58624), 
            .I2(n58310), .I3(n6_adj_5616), .O(n58429));
    defparam i4_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1525 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[12]_c [5]), 
            .I2(n58034), .I3(n6_adj_5590), .O(n25141));
    defparam i4_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i15729_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][5] ), 
            .I3(\Kp[5] ), .O(n29760));
    defparam i15729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_in_frame[17]_c [1]), .I1(n25141), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5617));
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1527 (.I0(\data_in_frame[19] [2]), .I1(n58429), 
            .I2(n4_adj_5617), .I3(n58526), .O(n58425));
    defparam i1_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1528 (.I0(n58253), .I1(n10_adj_5269), .I2(\data_out_frame[20] [0]), 
            .I3(n52835), .O(n58387));
    defparam i1_2_lut_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i21003_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3]_c [4]), 
            .I3(\Kp[4] ), .O(n29761));
    defparam i21003_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1529 (.I0(n26306), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58154));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1529.LUT_INIT = 16'h6666;
    SB_LUT4 i15731_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [3]), 
            .I3(\Kp[3] ), .O(n29762));
    defparam i15731_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1530 (.I0(n26463), .I1(n58160), .I2(Kp_23__N_1256), 
            .I3(GND_net), .O(n60258));
    defparam i2_3_lut_adj_1530.LUT_INIT = 16'h9696;
    SB_LUT4 i15732_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3][2] ), 
            .I3(\Kp[2] ), .O(n29763));
    defparam i15732_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15733_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n29764));
    defparam i15733_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1531 (.I0(n58272), .I1(n58316), .I2(n25974), 
            .I3(\data_in_frame[13] [1]), .O(n53833));
    defparam i1_4_lut_adj_1531.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1532 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n25771));
    defparam i2_3_lut_adj_1532.LUT_INIT = 16'h9696;
    SB_LUT4 i15734_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n29765));
    defparam i15734_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15735_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n29766));
    defparam i15735_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1533 (.I0(\data_in_frame[8]_c [7]), .I1(n58666), 
            .I2(n58549), .I3(n58284), .O(n25961));
    defparam i3_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 i15736_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n29767));
    defparam i15736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14362_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_13), 
            .I2(reset), .I3(n57974), .O(n7));
    defparam i14362_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1534 (.I0(\data_in_frame[15] [6]), .I1(Kp_23__N_1301), 
            .I2(GND_net), .I3(GND_net), .O(n58339));
    defparam i1_2_lut_adj_1534.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1535 (.I0(\data_in_frame[11] [5]), .I1(n58015), 
            .I2(n26294), .I3(n53743), .O(Kp_23__N_1256));
    defparam i3_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58148));
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1537 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25974));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'h6666;
    SB_LUT4 i23096_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n29768));
    defparam i23096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15738_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n29769));
    defparam i15738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1538 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n57916));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1538.LUT_INIT = 16'h5100;
    SB_LUT4 i23196_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11][2] ), 
            .I3(IntegralLimit[18]), .O(n29770));
    defparam i23196_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15740_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n29771));
    defparam i15740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1539 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58630));
    defparam i1_2_lut_adj_1539.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(n26493), .I1(n59815), .I2(GND_net), 
            .I3(GND_net), .O(n53770));
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1541 (.I0(\data_in_frame[12]_c [4]), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58163));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1541.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1542 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[12]_c [1]), 
            .O(n63250));
    defparam i1_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i15741_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n29772));
    defparam i15741_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15742_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [7]), 
            .I3(IntegralLimit[15]), .O(n29773));
    defparam i15742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_1057_i1_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), 
            .I2(\data_in_frame[3][0] ), .I3(\data_in_frame[19] [0]), .O(n4764[0]));
    defparam mux_1057_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_4_lut_adj_1543 (.I0(\data_in_frame[12]_c [6]), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[11][2] ), .I3(\data_in_frame[12] [0]), .O(n63252));
    defparam i1_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1544 (.I0(n63250), .I1(\data_in_frame[12]_c [5]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n63254));
    defparam i1_3_lut_adj_1544.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1545 (.I0(n58148), .I1(n63258), .I2(n63254), 
            .I3(n63252), .O(n63262));
    defparam i1_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1546 (.I0(n26294), .I1(n58287), .I2(n63262), 
            .I3(n58666), .O(n63268));
    defparam i1_4_lut_adj_1546.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1547 (.I0(n58068), .I1(n58413), .I2(n53348), 
            .I3(n63268), .O(n63274));
    defparam i1_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_LUT4 i15781_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n29812));
    defparam i15781_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1548 (.I0(n58090), .I1(n53770), .I2(n58250), 
            .I3(n63274), .O(n53720));
    defparam i1_4_lut_adj_1548.LUT_INIT = 16'h9669;
    SB_LUT4 i15780_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n29811));
    defparam i15780_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1549 (.I0(\data_in_frame[12]_c [5]), .I1(n26042), 
            .I2(GND_net), .I3(GND_net), .O(n58310));
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1550 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n57917));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1550.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1551 (.I0(\data_in_frame[13] [2]), .I1(n53720), 
            .I2(GND_net), .I3(GND_net), .O(n58316));
    defparam i1_2_lut_adj_1551.LUT_INIT = 16'h6666;
    SB_LUT4 i15778_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n29809));
    defparam i15778_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_4_lut_adj_1552 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[15] [7]), 
            .I2(\data_in_frame[13] [7]), .I3(n4_adj_5583), .O(n58160));
    defparam i2_4_lut_adj_1552.LUT_INIT = 16'h9669;
    SB_LUT4 i43216_2_lut_3_lut (.I0(n3472), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n58889));
    defparam i43216_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i3_2_lut_adj_1553 (.I0(n26330), .I1(n58160), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_5618));   // verilog/coms.v(88[17:63])
    defparam i3_2_lut_adj_1553.LUT_INIT = 16'h6666;
    SB_LUT4 mux_243_i16_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[15] ), .I3(encoder0_position_scaled[15]), 
            .O(\motor_state[15] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15777_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n29808));
    defparam i15777_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_4_lut_adj_1554 (.I0(n58630), .I1(\data_in_frame[13] [5]), 
            .I2(n25716), .I3(\data_in_frame[13] [3]), .O(n22_adj_5619));   // verilog/coms.v(88[17:63])
    defparam i9_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1555 (.I0(Kp_23__N_1256), .I1(n22_adj_5619), .I2(n16_adj_5618), 
            .I3(n58339), .O(n24_adj_5620));   // verilog/coms.v(88[17:63])
    defparam i11_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1556 (.I0(n60258), .I1(n24_adj_5620), .I2(n20_adj_5586), 
            .I3(n25961), .O(n52776));   // verilog/coms.v(88[17:63])
    defparam i12_4_lut_adj_1556.LUT_INIT = 16'h9669;
    SB_LUT4 mux_243_i19_3_lut_4_lut (.I0(\control_mode[1] ), .I1(n25541), 
            .I2(\motor_state_23__N_91[18] ), .I3(encoder0_position_scaled[18]), 
            .O(\motor_state[18] ));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15776_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n29807));
    defparam i15776_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(n26330), .I1(n53776), .I2(GND_net), 
            .I3(GND_net), .O(n58657));
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i54355_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n59012));
    defparam i54355_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i2_3_lut_adj_1558 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[6] [1]), .I3(GND_net), .O(n58733));
    defparam i2_3_lut_adj_1558.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1559 (.I0(n53348), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58422));
    defparam i1_2_lut_adj_1559.LUT_INIT = 16'h6666;
    SB_LUT4 i15753_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n29784));
    defparam i15753_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i22526_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n29783));
    defparam i22526_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15751_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n29782));
    defparam i15751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15750_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n29781));
    defparam i15750_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_780_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5579));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15749_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n29780));
    defparam i15749_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1560 (.I0(n25862), .I1(n25947), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1067));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1560.LUT_INIT = 16'h6666;
    SB_LUT4 i15748_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [1]), 
            .I3(IntegralLimit[9]), .O(n29779));
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1561 (.I0(n58169), .I1(n25898), .I2(Kp_23__N_974), 
            .I3(n26466), .O(n62948));
    defparam i1_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1562 (.I0(Kp_23__N_1067), .I1(n26294), .I2(n58229), 
            .I3(n62948), .O(n62954));
    defparam i1_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1563 (.I0(n58520), .I1(n53774), .I2(n53728), 
            .I3(n62954), .O(n25103));
    defparam i1_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(\data_in_frame[9] [0]), .I1(n25103), 
            .I2(GND_net), .I3(GND_net), .O(n58090));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25716));
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [0]), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5578));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1567 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n57918));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1567.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(\data_in_frame[11] [7]), .I1(n53066), 
            .I2(GND_net), .I3(GND_net), .O(n58405));
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26274));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1570 (.I0(n26274), .I1(\data_in_frame[12]_c [2]), 
            .I2(n26853), .I3(n58012), .O(n10_adj_5582));
    defparam i4_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5577));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1571 (.I0(n26829), .I1(\data_in_frame[8] [2]), 
            .I2(n25933), .I3(GND_net), .O(n3_adj_5376));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1571.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1572 (.I0(\data_in_frame[9][7] ), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58128));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1572.LUT_INIT = 16'h6666;
    SB_LUT4 i15747_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [2]), 
            .I3(IntegralLimit[10]), .O(n29778));
    defparam i15747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1573 (.I0(\data_in_frame[8]_c [1]), .I1(\data_in_frame[7]_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58660));
    defparam i1_2_lut_adj_1573.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1574 (.I0(\data_in_frame[12]_c [2]), .I1(n52885), 
            .I2(\data_in_frame[12]_c [3]), .I3(GND_net), .O(n58250));
    defparam i2_3_lut_adj_1574.LUT_INIT = 16'h9696;
    SB_LUT4 i15746_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [3]), 
            .I3(IntegralLimit[11]), .O(n29777));
    defparam i15746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1575 (.I0(n25755), .I1(n58660), .I2(\data_in_frame[7]_c [6]), 
            .I3(\data_in_frame[10] [2]), .O(n63284));
    defparam i1_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i15775_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n29806));
    defparam i15775_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(n58608), .I1(n58397), .I2(n25898), 
            .I3(n63284), .O(n59815));
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1577 (.I0(n59815), .I1(n58250), .I2(\data_in_frame[14] [4]), 
            .I3(GND_net), .O(n26379));
    defparam i2_3_lut_adj_1577.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1578 (.I0(\data_in_frame[8]_c [0]), .I1(\data_in_frame[7]_c [7]), 
            .I2(n58290), .I3(\data_in_frame[1] [5]), .O(n58556));
    defparam i3_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i15774_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n29805));
    defparam i15774_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1579 (.I0(n58166), .I1(n58556), .I2(n26398), 
            .I3(GND_net), .O(n25898));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1579.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1580 (.I0(n25898), .I1(n52731), .I2(GND_net), 
            .I3(GND_net), .O(n58413));
    defparam i1_2_lut_adj_1580.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(\data_in_frame[10] [1]), .I1(n26829), 
            .I2(n58413), .I3(\data_in_frame[9][7] ), .O(n26853));
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(\data_in_frame[12]_c [3]), .I1(n26853), 
            .I2(GND_net), .I3(GND_net), .O(n58173));
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1583 (.I0(n58507), .I1(n58540), .I2(\data_in_frame[10] [3]), 
            .I3(n58078), .O(n12_adj_5621));   // verilog/coms.v(79[16:43])
    defparam i5_4_lut_adj_1583.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1584 (.I0(\data_in_frame[8] [2]), .I1(n12_adj_5621), 
            .I2(n58660), .I3(\data_in_frame[5] [5]), .O(n26493));   // verilog/coms.v(79[16:43])
    defparam i6_4_lut_adj_1584.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1585 (.I0(\data_in_frame[14] [5]), .I1(n26493), 
            .I2(n58173), .I3(\data_in_frame[12]_c [4]), .O(n52778));
    defparam i3_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15773_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n29804));
    defparam i15773_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_4_lut_adj_1586 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[1]_c [3]), .I3(n58060), .O(n58511));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(\data_in_frame[16] [6]), .I1(n26379), 
            .I2(GND_net), .I3(GND_net), .O(n58526));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1588 (.I0(\data_in_frame[18][7] ), .I1(\data_in_frame[18]_c [6]), 
            .I2(GND_net), .I3(GND_net), .O(n25908));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1588.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1589 (.I0(n25908), .I1(n58526), .I2(n52778), 
            .I3(GND_net), .O(n58714));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_adj_1589.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1590 (.I0(\data_in_frame[5] [0]), .I1(n58733), 
            .I2(n58245), .I3(\data_in_frame[11] [6]), .O(n28_adj_5622));
    defparam i10_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1591 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n58530));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1591.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_1592 (.I0(n58157), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[6] [2]), .I3(\data_in_frame[9] [5]), .O(n31_adj_5623));
    defparam i13_4_lut_adj_1592.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1593 (.I0(n25103), .I1(n58589), .I2(n58766), 
            .I3(n58297), .O(n30_adj_5624));
    defparam i12_4_lut_adj_1593.LUT_INIT = 16'h6996;
    SB_LUT4 i13942_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3472), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n27972));   // verilog/coms.v(158[12:15])
    defparam i13942_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i15772_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n29803));
    defparam i15772_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut_adj_1594 (.I0(n31_adj_5623), .I1(\data_in_frame[6] [0]), 
            .I2(n28_adj_5622), .I3(\data_in_frame[6] [5]), .O(n34_adj_5625));
    defparam i16_4_lut_adj_1594.LUT_INIT = 16'h6996;
    SB_LUT4 i15771_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n29802));
    defparam i15771_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_4_lut_adj_1595 (.I0(n52885), .I1(n58012), .I2(n58422), 
            .I3(\data_in_frame[7] [1]), .O(n29_adj_5626));
    defparam i11_4_lut_adj_1595.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(\data_in_frame[14] [2]), .I1(n29_adj_5626), 
            .I2(n34_adj_5625), .I3(n30_adj_5624), .O(n53776));
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'h9669;
    SB_LUT4 i15770_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n29801));
    defparam i15770_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1597 (.I0(\data_in_frame[19] [0]), .I1(n53776), 
            .I2(n58714), .I3(n58093), .O(n58672));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1597.LUT_INIT = 16'h9669;
    SB_LUT4 i15754_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n29785));
    defparam i15754_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1598 (.I0(n58078), .I1(\data_in_frame[5] [5]), 
            .I2(n25915), .I3(GND_net), .O(n58290));
    defparam i2_3_lut_adj_1598.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1599 (.I0(n26337), .I1(n58138), .I2(n26667), 
            .I3(\data_in_frame[7] [1]), .O(n58549));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i15755_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n29786));
    defparam i15755_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15756_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n29787));
    defparam i15756_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15758_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n29789));
    defparam i15758_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15759_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n29790));
    defparam i15759_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15760_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n29791));
    defparam i15760_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15761_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n29792));
    defparam i15761_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15762_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n29793));
    defparam i15762_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15763_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n29794));
    defparam i15763_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_780_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5521));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1600 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n25529), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_5452));
    defparam i1_3_lut_4_lut_adj_1600.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_4_lut_adj_1601 (.I0(n25705), .I1(n10_c), .I2(n26261), 
            .I3(\data_out_frame[21] [6]), .O(n58757));
    defparam i1_2_lut_4_lut_adj_1601.LUT_INIT = 16'h6996;
    SB_LUT4 i22410_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n29795));
    defparam i22410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15765_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n29796));
    defparam i15765_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15766_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n29797));
    defparam i15766_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_780_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15767_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n29798));
    defparam i15767_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15768_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n29799));
    defparam i15768_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [0]), 
            .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'ha088;
    SB_LUT4 i15769_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n29800));
    defparam i15769_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_780_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5518));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15745_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [4]), 
            .I3(IntegralLimit[12]), .O(n29776));
    defparam i15745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_780_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5516));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5515));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15743_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [6]), 
            .I3(IntegralLimit[14]), .O(n29774));
    defparam i15743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i22941_3_lut_4_lut (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(\data_in_frame[12]_c [5]), 
            .I3(IntegralLimit[13]), .O(n29775));
    defparam i22941_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_780_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n70291_bdd_4_lut (.I0(n70291), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n70294));
    defparam n70291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i43256_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_13), 
            .I2(n57974), .I3(reset), .O(n58929));   // verilog/coms.v(157[7:23])
    defparam i43256_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 select_780_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5512));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1603 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [6]), 
            .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5509));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1603.LUT_INIT = 16'ha088;
    SB_LUT4 select_780_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5508));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [4]), 
            .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1605 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5589), .I3(n57968), .O(n26923));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1605.LUT_INIT = 16'haaa8;
    SB_LUT4 select_780_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5504));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1606 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n57919));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1606.LUT_INIT = 16'h5100;
    SB_LUT4 i2_3_lut_3_lut (.I0(LED_N_3408), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(reset), .I3(GND_net), .O(n22760));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_4_lut_adj_1607 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [0]), 
            .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'ha088;
    SB_LUT4 i1_3_lut_4_lut_adj_1608 (.I0(\data_in_frame[18][3] ), .I1(\data_in_frame[18] [5]), 
            .I2(\data_in_frame[21][3] ), .I3(\data_in_frame[23] [1]), .O(n63172));
    defparam i1_3_lut_4_lut_adj_1608.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i28280_2_lut (.I0(LED_c), .I1(LED_N_3408), .I2(GND_net), .I3(GND_net), 
            .O(LED_N_3407));   // verilog/coms.v(253[15] 255[9])
    defparam i28280_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 select_780_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14797_4_lut (.I0(n2874), .I1(LED_N_3407), .I2(n27276), .I3(\FRAME_MATCHER.i_31__N_2513 ), 
            .O(n28828));   // verilog/coms.v(130[12] 305[6])
    defparam i14797_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 select_780_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5497));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_1651_Select_0_i3_3_lut (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n3_adj_5627));   // verilog/coms.v(148[4] 304[11])
    defparam select_1651_Select_0_i3_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_780_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5496));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(LED_c), .I1(n3_adj_5627), .I2(Kp_23__N_1748), 
            .I3(Kp_23__N_612), .O(n5_adj_5573));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'hfcec;
    SB_LUT4 select_780_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5494));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1610 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [0]), 
            .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1610.LUT_INIT = 16'ha088;
    SB_LUT4 select_1653_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5572));   // verilog/coms.v(148[4] 304[11])
    defparam select_1653_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_780_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5492));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1611 (.I0(n25915), .I1(n58397), .I2(\data_in_frame[8]_c [0]), 
            .I3(GND_net), .O(n53607));
    defparam i1_2_lut_3_lut_adj_1611.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_150_i2_4_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_150_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1612 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n57920));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1612.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1613 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[3][5] ), .I3(GND_net), .O(n58166));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1613.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5489));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54534 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n70285));
    defparam byte_transmit_counter_0__bdd_4_lut_54534.LUT_INIT = 16'he4aa;
    SB_LUT4 select_780_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5488));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5487));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n70285_bdd_4_lut (.I0(n70285), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n70288));
    defparam n70285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1614 (.I0(\data_in_frame[5] [0]), .I1(n25813), 
            .I2(n26343), .I3(GND_net), .O(n26337));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1614.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1615 (.I0(\data_in_frame[1]_c [4]), .I1(n58256), 
            .I2(n58540), .I3(\data_in_frame[5] [7]), .O(n25933));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1615.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1616 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n57921));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1616.LUT_INIT = 16'h5100;
    SB_LUT4 i1_3_lut_4_lut_adj_1617 (.I0(\data_in_frame[1]_c [1]), .I1(\data_in_frame[0]_c [6]), 
            .I2(\data_in_frame[1]_c [0]), .I3(\data_in_frame[3][2] ), .O(n58300));   // verilog/coms.v(73[16:27])
    defparam i1_3_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1618 (.I0(\data_in_frame[1]_c [4]), .I1(n58256), 
            .I2(\data_in_frame[5] [6]), .I3(n58607), .O(n58397));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1618.LUT_INIT = 16'h9669;
    SB_LUT4 i11_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(\data_in_frame[20] [7]), 
            .I3(rx_data[7]), .O(n57449));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i15405_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29436));
    defparam i15405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(\data_in_frame[20] [5]), 
            .I3(rx_data[5]), .O(n9_adj_5534));
    defparam i17_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1619 (.I0(\data_in_frame[2][0] ), .I1(\data_in_frame[3]_c [6]), 
            .I2(\data_in_frame[4] [1]), .I3(GND_net), .O(n6_adj_5340));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1619.LUT_INIT = 16'h9696;
    SB_LUT4 i15399_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(rx_data[4]), 
            .I3(\data_in_frame[20][4] ), .O(n29430));
    defparam i15399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15396_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(rx_data[3]), 
            .I3(\data_in_frame[20][3] ), .O(n29427));
    defparam i15396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(\data_in_frame[20] [2]), 
            .I3(rx_data[2]), .O(n25_adj_5533));
    defparam i33_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i15389_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(rx_data[1]), 
            .I3(\data_in_frame[20][1] ), .O(n29420));
    defparam i15389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54529 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n70279));
    defparam byte_transmit_counter_0__bdd_4_lut_54529.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1620 (.I0(\data_out_frame[25] [6]), .I1(n26382), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5628));
    defparam i1_2_lut_adj_1620.LUT_INIT = 16'h6666;
    SB_LUT4 i15385_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57983), .I2(rx_data[0]), 
            .I3(\data_in_frame[20][0] ), .O(n29416));
    defparam i15385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_780_Select_223_i3_4_lut (.I0(n5_adj_5628), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\data_out_frame[25] [5]), .I3(n53902), .O(n3_adj_5565));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_223_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(n52894), .I3(GND_net), .O(n58702));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1622 (.I0(\data_out_frame[7] [5]), .I1(n58468), 
            .I2(\data_out_frame[12] [1]), .I3(\data_out_frame[7] [4]), .O(n14));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1622.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1623 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n58021));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1623.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_222_i3_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5580), .I3(n58214), 
            .O(n3_adj_5564));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_780_Select_221_i3_4_lut (.I0(n53918), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58731), .I3(\data_out_frame[25] [4]), .O(n3_adj_5563));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_221_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_3_lut_adj_1624 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[10] [2]), .I3(GND_net), .O(n42_adj_5311));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1624.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1625 (.I0(\data_out_frame[25] [3]), .I1(n53763), 
            .I2(GND_net), .I3(GND_net), .O(n53918));
    defparam i1_2_lut_adj_1625.LUT_INIT = 16'h6666;
    SB_LUT4 i15444_3_lut_4_lut (.I0(n28338), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[1][7] ), .O(n29475));
    defparam i15444_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n70279_bdd_4_lut (.I0(n70279), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n70282));
    defparam n70279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1626 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n26558));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1626.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1627 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[14] [5]), 
            .O(n58333));
    defparam i2_3_lut_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1628 (.I0(\data_out_frame[7] [5]), .I1(n58468), 
            .I2(n10_adj_5321), .I3(\data_out_frame[5] [7]), .O(n26249));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1628.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1629 (.I0(\data_out_frame[16] [5]), .I1(n58690), 
            .I2(n58739), .I3(GND_net), .O(n58636));
    defparam i1_2_lut_3_lut_adj_1629.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1630 (.I0(\data_out_frame[10] [1]), .I1(n58142), 
            .I2(\data_out_frame[7] [7]), .I3(n52894), .O(n53891));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1630.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_220_i3_4_lut (.I0(n58723), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5587), .I3(\data_out_frame[22] [6]), .O(n3_adj_5562));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_220_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i23458_3_lut (.I0(\control_mode[0] ), .I1(\data_in_frame[1]_c [0]), 
            .I2(n22773), .I3(GND_net), .O(n29616));
    defparam i23458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15438_3_lut_4_lut (.I0(n28338), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[1][6] ), .O(n29469));
    defparam i15438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_780_Select_219_i3_4_lut (.I0(n58639), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58760), .I3(\data_out_frame[24] [7]), .O(n3_adj_5561));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_219_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_4_lut_adj_1631 (.I0(\data_in_frame[1]_c [0]), .I1(\data_in_frame[1][2] ), 
            .I2(\data_in_frame[1]_c [1]), .I3(n58511), .O(n25884));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_4_lut_adj_1631.LUT_INIT = 16'h6996;
    SB_LUT4 i15435_3_lut_4_lut (.I0(n28338), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29466));
    defparam i15435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1632 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[8] [5]), 
            .I2(n25680), .I3(n58071), .O(n58543));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1632.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1633 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n25680));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1633.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1634 (.I0(\data_in_frame[7]_c [6]), .I1(n25915), 
            .I2(n25755), .I3(GND_net), .O(n23933));
    defparam i1_2_lut_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 i15432_3_lut_4_lut (.I0(n28338), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[1]_c [4]), .O(n29463));
    defparam i15432_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15429_3_lut_4_lut (.I0(n28338), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[1]_c [3]), .O(n29460));
    defparam i15429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1635 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(n58601), .I3(GND_net), .O(n58031));
    defparam i1_2_lut_3_lut_adj_1635.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_4_lut (.I0(\data_out_frame[18] [1]), .I1(n58690), .I2(n58739), 
            .I3(n58373), .O(n58534));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'ha55a;
    SB_LUT4 i2_2_lut_adj_1636 (.I0(n58351), .I1(\data_out_frame[25] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5630));
    defparam i2_2_lut_adj_1636.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n70501));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i15420_3_lut_4_lut (.I0(n28338), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[1]_c [0]), .O(n29451));
    defparam i15420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15903_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[7]), 
            .I3(\data_in_frame[8]_c [7]), .O(n29934));
    defparam i15903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_780_Select_218_i3_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5630), .I3(n60186), 
            .O(n3_adj_5560));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i15900_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[6]), 
            .I3(\data_in_frame[8][6] ), .O(n29931));
    defparam i15900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15897_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[5]), 
            .I3(\data_in_frame[8]_c [5]), .O(n29928));
    defparam i15897_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15894_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n29925));
    defparam i15894_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15890_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[3]), 
            .I3(\data_in_frame[8][3] ), .O(n29921));
    defparam i15890_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15887_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n29918));
    defparam i15887_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15884_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[1]), 
            .I3(\data_in_frame[8]_c [1]), .O(n29915));
    defparam i15884_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1637 (.I0(n26865), .I1(n60779), .I2(\data_out_frame[23] [1]), 
            .I3(GND_net), .O(n58408));
    defparam i2_3_lut_adj_1637.LUT_INIT = 16'h6969;
    SB_LUT4 i15880_3_lut_4_lut (.I0(n8), .I1(n57986), .I2(rx_data[0]), 
            .I3(\data_in_frame[8]_c [0]), .O(n29911));
    defparam i15880_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1638 (.I0(\data_out_frame[15] [0]), .I1(n58751), 
            .I2(n58769), .I3(\data_out_frame[15] [1]), .O(n58690));
    defparam i2_3_lut_4_lut_adj_1638.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_3_lut (.I0(reset), .I1(Kp_23__N_612), .I2(Kp_23__N_1748), 
            .I3(GND_net), .O(n22773));   // verilog/coms.v(130[12] 305[6])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i3_4_lut_adj_1639 (.I0(n59988), .I1(n58644), .I2(n58366), 
            .I3(n58361), .O(n60779));
    defparam i3_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1640 (.I0(n25705), .I1(n10_c), .I2(n26261), 
            .I3(\data_out_frame[19] [3]), .O(n58570));
    defparam i1_2_lut_4_lut_adj_1640.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1641 (.I0(\data_out_frame[16] [4]), .I1(n58360), 
            .I2(GND_net), .I3(GND_net), .O(n58361));
    defparam i1_2_lut_adj_1641.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1642 (.I0(n26561), .I1(n25733), .I2(n26280), 
            .I3(GND_net), .O(n58565));
    defparam i2_3_lut_adj_1642.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1643 (.I0(n58183), .I1(n58565), .I2(n58361), 
            .I3(n60779), .O(n12_adj_5631));
    defparam i5_4_lut_adj_1643.LUT_INIT = 16'h6996;
    SB_LUT4 i8_2_lut_3_lut (.I0(n58142), .I1(\data_out_frame[4] [1]), .I2(\data_out_frame[6] [2]), 
            .I3(GND_net), .O(n30));
    defparam i8_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15929_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[7]), 
            .I3(\data_in_frame[9][7] ), .O(n29960));
    defparam i15929_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15926_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29957));
    defparam i15926_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15922_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29953));
    defparam i15922_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_780_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n70501_bdd_4_lut (.I0(n70501), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n63832));
    defparam n70501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15919_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29950));
    defparam i15919_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1644 (.I0(n53875), .I1(n12_adj_5631), .I2(n58720), 
            .I3(\data_out_frame[20] [6]), .O(n60186));
    defparam i6_4_lut_adj_1644.LUT_INIT = 16'h9669;
    SB_LUT4 i15916_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29947));
    defparam i15916_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15913_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29944));
    defparam i15913_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [0]), 
            .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5484));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'ha088;
    SB_LUT4 i15910_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29941));
    defparam i15910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_780_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n70126), .I2(n66452), .I3(byte_transmit_counter[4]), .O(n70495));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i15906_3_lut_4_lut (.I0(n8_adj_8), .I1(n57986), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29937));
    defparam i15906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[13] [1]), .I1(n26618), .I2(\data_out_frame[10] [5]), 
            .I3(n58081), .O(n26_c));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5482));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15956_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n29987));
    defparam i15956_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15952_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n29983));
    defparam i15952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15949_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n29980));
    defparam i15949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15946_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n29977));
    defparam i15946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15942_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n29973));
    defparam i15942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15939_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n29970));
    defparam i15939_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15936_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n29967));
    defparam i15936_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15932_3_lut_4_lut (.I0(n8_adj_11), .I1(n57986), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29963));
    defparam i15932_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54524 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n70267));
    defparam byte_transmit_counter_0__bdd_4_lut_54524.LUT_INIT = 16'he4aa;
    SB_LUT4 i15982_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n30013));
    defparam i15982_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15979_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n30010));
    defparam i15979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15976_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n30007));
    defparam i15976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1646 (.I0(n52743), .I1(n58565), .I2(n58408), 
            .I3(n53831), .O(n58723));
    defparam i3_4_lut_adj_1646.LUT_INIT = 16'h9669;
    SB_LUT4 i53559_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(\data_in_frame[11] [4]), 
            .I3(rx_data[4]), .O(n57339));
    defparam i53559_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i15969_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n30000));
    defparam i15969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n70267_bdd_4_lut (.I0(n70267), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n70270));
    defparam n70267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1647 (.I0(n59809), .I1(n58723), .I2(n60186), 
            .I3(n53785), .O(n58760));
    defparam i3_4_lut_adj_1647.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1648 (.I0(\data_out_frame[10] [1]), .I1(n58142), 
            .I2(\data_out_frame[7] [7]), .I3(n26249), .O(n58275));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1648.LUT_INIT = 16'h6996;
    SB_LUT4 i15962_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n29993));
    defparam i15962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15959_3_lut_4_lut (.I0(n28322), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n29990));
    defparam i15959_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1649 (.I0(\data_out_frame[16] [0]), .I1(n52801), 
            .I2(n58687), .I3(GND_net), .O(n6_adj_5265));
    defparam i1_2_lut_3_lut_adj_1649.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1650 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n1516), .I3(n26249), .O(n58751));
    defparam i1_2_lut_4_lut_adj_1650.LUT_INIT = 16'h6996;
    SB_LUT4 n70495_bdd_4_lut (.I0(n70495), .I1(n70228), .I2(n57571), .I3(byte_transmit_counter[4]), 
            .O(tx_data[0]));
    defparam n70495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1651 (.I0(n52786), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n53902));
    defparam i1_2_lut_adj_1651.LUT_INIT = 16'h6666;
    SB_LUT4 i16009_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[7]), 
            .I3(\data_in_frame[12]_c [7]), .O(n30040));
    defparam i16009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16006_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[6]), 
            .I3(\data_in_frame[12]_c [6]), .O(n30037));
    defparam i16006_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n63887), .I2(n63888), .I3(\byte_transmit_counter[2] ), 
            .O(n70261));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i16002_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[5]), 
            .I3(\data_in_frame[12]_c [5]), .O(n30033));
    defparam i16002_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1652 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[5] [4]), .O(n9));
    defparam i1_2_lut_4_lut_adj_1652.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1653 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1]_c [1]), 
            .I2(\data_in_frame[0]_c [7]), .I3(\data_in_frame[3] [3]), .O(n58078));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i15999_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[4]), 
            .I3(\data_in_frame[12]_c [4]), .O(n30030));
    defparam i15999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1654 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1]_c [1]), 
            .I2(n58511), .I3(GND_net), .O(Kp_23__N_767));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_adj_1654.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(\data_out_frame[12] [4]), .I1(n1516), 
            .I2(n26249), .I3(GND_net), .O(n1655));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'h9696;
    SB_LUT4 i11_3_lut_4_lut_adj_1656 (.I0(n26618), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [5]), .I3(n58711), .O(n32));
    defparam i11_3_lut_4_lut_adj_1656.LUT_INIT = 16'h6996;
    SB_LUT4 i15996_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[3]), 
            .I3(\data_in_frame[12]_c [3]), .O(n30027));
    defparam i15996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54702 (.I0(byte_transmit_counter[3]), 
            .I1(n70132), .I2(n66247), .I3(byte_transmit_counter[4]), .O(n70483));
    defparam byte_transmit_counter_3__bdd_4_lut_54702.LUT_INIT = 16'he4aa;
    SB_LUT4 i15992_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[2]), 
            .I3(\data_in_frame[12]_c [2]), .O(n30023));
    defparam i15992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15989_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[1]), 
            .I3(\data_in_frame[12]_c [1]), .O(n30020));
    defparam i15989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1657 (.I0(\data_out_frame[12] [4]), .I1(n1516), 
            .I2(n58739), .I3(n58197), .O(n14_adj_5632));   // verilog/coms.v(78[16:43])
    defparam i5_3_lut_4_lut_adj_1657.LUT_INIT = 16'h6996;
    SB_LUT4 i15986_3_lut_4_lut (.I0(n8_adj_5536), .I1(n57986), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n30017));
    defparam i15986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_2_lut_adj_1658 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[21] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5633));
    defparam i3_2_lut_adj_1658.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1659 (.I0(n25819), .I1(n58205), .I2(n58562), 
            .I3(\data_out_frame[16] [5]), .O(n22_adj_5634));
    defparam i9_4_lut_adj_1659.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[4] [5]), .I1(n58284), .I2(\data_in_frame[8]_c [7]), 
            .I3(GND_net), .O(n7_adj_5377));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 n70261_bdd_4_lut (.I0(n70261), .I1(n63909), .I2(n63908), .I3(\byte_transmit_counter[2] ), 
            .O(n70264));
    defparam n70261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16034_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n30065));
    defparam i16034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_adj_1660 (.I0(n60912), .I1(n58408), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n20_adj_5635));
    defparam i7_3_lut_adj_1660.LUT_INIT = 16'h6969;
    SB_LUT4 i11_4_lut_adj_1661 (.I0(n26427), .I1(n22_adj_5634), .I2(n16_adj_5633), 
            .I3(n58687), .O(n24_adj_5636));
    defparam i11_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i16031_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n30062));
    defparam i16031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54515 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n70255));
    defparam byte_transmit_counter_0__bdd_4_lut_54515.LUT_INIT = 16'he4aa;
    SB_LUT4 i16028_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n30059));
    defparam i16028_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1662 (.I0(\data_in_frame[4] [5]), .I1(n58284), 
            .I2(n53348), .I3(GND_net), .O(n53728));
    defparam i1_2_lut_3_lut_adj_1662.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1663 (.I0(\data_out_frame[22] [7]), .I1(n24_adj_5636), 
            .I2(n20_adj_5635), .I3(\data_out_frame[23] [2]), .O(n53763));
    defparam i12_4_lut_adj_1663.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1664 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n58057));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1664.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1665 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n25676));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1665.LUT_INIT = 16'h9696;
    SB_LUT4 i16025_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n30056));
    defparam i16025_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1666 (.I0(n58742), .I1(n53763), .I2(n53902), 
            .I3(n58760), .O(n10_adj_5637));
    defparam i4_4_lut_adj_1666.LUT_INIT = 16'h6996;
    SB_LUT4 i16022_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n30053));
    defparam i16022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1667 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n26340), .I3(Kp_23__N_878), .O(n58284));   // verilog/coms.v(80[16:43])
    defparam i2_3_lut_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 i16019_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n30050));
    defparam i16019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n70255_bdd_4_lut (.I0(n70255), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n70258));
    defparam n70255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16016_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n30047));
    defparam i16016_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1668 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n58733), .I3(n25912), .O(n58226));   // verilog/coms.v(80[16:43])
    defparam i2_3_lut_4_lut_adj_1668.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1669 (.I0(\data_out_frame[8] [5]), .I1(n25680), 
            .I2(\data_out_frame[10] [7]), .I3(n10_adj_5271), .O(n26261));   // verilog/coms.v(78[16:43])
    defparam i5_3_lut_4_lut_adj_1669.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_217_i3_4_lut (.I0(n58293), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5637), .I3(n58731), .O(n3_adj_5559));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i16012_3_lut_4_lut (.I0(n8_adj_9), .I1(n57986), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n30043));
    defparam i16012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16061_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n30092));
    defparam i16061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16058_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n30089));
    defparam i16058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16054_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n30085));
    defparam i16054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16051_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n30082));
    defparam i16051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1670 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n26865));
    defparam i1_2_lut_3_lut_adj_1670.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1671 (.I0(\data_out_frame[8] [5]), .I1(n25680), 
            .I2(n58071), .I3(GND_net), .O(n26431));   // verilog/coms.v(78[16:43])
    defparam i2_2_lut_3_lut_adj_1671.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1672 (.I0(\data_out_frame[25] [0]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5638));
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1673 (.I0(n58346), .I1(\data_out_frame[22] [4]), 
            .I2(n52835), .I3(n6_adj_5638), .O(n58351));
    defparam i4_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 i51173_2_lut (.I0(displacement[8]), .I1(\control_mode[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n66494));
    defparam i51173_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i26_4_lut (.I0(encoder1_position_scaled[8]), .I1(n66494), .I2(n15), 
            .I3(n37407), .O(n12_adj_5603));
    defparam i26_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16048_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n30079));
    defparam i16048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16044_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n30075));
    defparam i16044_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1674 (.I0(\data_out_frame[7] [2]), .I1(n58552), 
            .I2(n10_adj_5289), .I3(\data_out_frame[11] [6]), .O(n26704));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n57355));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_780_Select_216_i3_3_lut (.I0(n58293), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58351), .I3(GND_net), .O(n3_adj_5558));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_216_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_3_lut_adj_1675 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n58693));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1675.LUT_INIT = 16'h9696;
    SB_LUT4 i16038_3_lut_4_lut (.I0(n28314), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n30069));
    defparam i16038_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1676 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[5] [6]), .O(n58699));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1677 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58575));
    defparam i1_2_lut_adj_1677.LUT_INIT = 16'h6666;
    SB_LUT4 i16088_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n30119));
    defparam i16088_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16084_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n30115));
    defparam i16084_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1678 (.I0(n52801), .I1(\data_out_frame[13] [5]), 
            .I2(n25082), .I3(GND_net), .O(n53757));
    defparam i1_2_lut_3_lut_adj_1678.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1679 (.I0(\data_out_frame[16] [4]), .I1(n26235), 
            .I2(n58202), .I3(n6_adj_5585), .O(n59988));
    defparam i4_4_lut_adj_1679.LUT_INIT = 16'h6996;
    SB_LUT4 n70483_bdd_4_lut (.I0(n70483), .I1(n14_adj_5542), .I2(n7_adj_5599), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n70483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1680 (.I0(\data_out_frame[21] [0]), .I1(n59988), 
            .I2(GND_net), .I3(GND_net), .O(n52743));
    defparam i1_2_lut_adj_1680.LUT_INIT = 16'h9999;
    SB_LUT4 i16081_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n30112));
    defparam i16081_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16078_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n30109));
    defparam i16078_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16074_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n30105));
    defparam i16074_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16071_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n30102));
    defparam i16071_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54505 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n70249));
    defparam byte_transmit_counter_0__bdd_4_lut_54505.LUT_INIT = 16'he4aa;
    SB_LUT4 i16068_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n30099));
    defparam i16068_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1681 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n58523));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1681.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1682 (.I0(\data_out_frame[16] [3]), .I1(n26111), 
            .I2(n10_adj_5282), .I3(\data_out_frame[19] [1]), .O(n58474));
    defparam i5_3_lut_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1683 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[22] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58720));
    defparam i1_2_lut_adj_1683.LUT_INIT = 16'h6666;
    SB_LUT4 i16064_3_lut_4_lut (.I0(n42296), .I1(n57986), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n30095));
    defparam i16064_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1684 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n58609));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1684.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1685 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58214));
    defparam i1_2_lut_adj_1685.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1686 (.I0(\data_out_frame[18] [5]), .I1(n60912), 
            .I2(n53891), .I3(n26405), .O(n58360));
    defparam i3_4_lut_adj_1686.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54707 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n70477));
    defparam byte_transmit_counter_0__bdd_4_lut_54707.LUT_INIT = 16'he4aa;
    SB_LUT4 n70249_bdd_4_lut (.I0(n70249), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n70252));
    defparam n70249_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1687 (.I0(n52831), .I1(\data_out_frame[21] [1]), 
            .I2(n58360), .I3(n6_adj_5584), .O(n52786));
    defparam i4_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1688 (.I0(\data_out_frame[25] [6]), .I1(n58442), 
            .I2(n58639), .I3(n58214), .O(n30_adj_5639));
    defparam i11_4_lut_adj_1688.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1689 (.I0(\data_out_frame[20] [1]), .I1(n58757), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5640));
    defparam i4_2_lut_adj_1689.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1690 (.I0(n58654), .I1(n52883), .I2(n58346), 
            .I3(n52786), .O(n24_adj_5641));
    defparam i10_4_lut_adj_1690.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1691 (.I0(tx_active), .I1(r_SM_Main[1]), .I2(n61386), 
            .I3(n85), .O(n53949));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut_adj_1691.LUT_INIT = 16'h3aba;
    SB_LUT4 i8_4_lut_adj_1692 (.I0(n58720), .I1(n53746), .I2(n52743), 
            .I3(n58355), .O(n22_adj_5642));
    defparam i8_4_lut_adj_1692.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1693 (.I0(n58461), .I1(n24_adj_5641), .I2(n18_adj_5640), 
            .I3(\data_out_frame[21] [7]), .O(n26_adj_5643));
    defparam i12_4_lut_adj_1693.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1694 (.I0(\data_out_frame[20] [5]), .I1(n26_adj_5643), 
            .I2(n22_adj_5642), .I3(n59809), .O(n60672));
    defparam i13_4_lut_adj_1694.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1695 (.I0(\data_out_frame[25] [3]), .I1(n30_adj_5639), 
            .I2(n26382), .I3(n58343), .O(n34_adj_5644));
    defparam i15_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1696 (.I0(\data_out_frame[23] [7]), .I1(n58575), 
            .I2(\data_out_frame[24] [6]), .I3(n58369), .O(n32_adj_5645));
    defparam i13_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 i27113_3_lut (.I0(control_mode_c[4]), .I1(\data_in_frame[1]_c [4]), 
            .I2(n22773), .I3(GND_net), .O(n29638));
    defparam i27113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1697 (.I0(\data_out_frame[23] [0]), .I1(n53855), 
            .I2(\data_out_frame[24] [5]), .I3(\data_out_frame[23] [5]), 
            .O(n33));
    defparam i14_4_lut_adj_1697.LUT_INIT = 16'h6996;
    SB_LUT4 i51672_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n66309));   // verilog/coms.v(158[12:15])
    defparam i51672_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_1698 (.I0(\data_out_frame[23] [1]), .I1(n58742), 
            .I2(n60672), .I3(n58281), .O(n31_adj_5646));
    defparam i12_4_lut_adj_1698.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_1699 (.I0(n31_adj_5646), .I1(n33), .I2(n32_adj_5645), 
            .I3(n34_adj_5644), .O(n58293));
    defparam i18_4_lut_adj_1699.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(n70180), .I2(n63832), .I3(byte_transmit_counter[3]), .O(n70243));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70243_bdd_4_lut (.I0(n70243), .I1(n63735), .I2(n63734), .I3(byte_transmit_counter[3]), 
            .O(n70246));
    defparam n70243_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_54495 (.I0(\byte_transmit_counter[2] ), 
            .I1(n70174), .I2(n70204), .I3(byte_transmit_counter[3]), .O(n70237));
    defparam byte_transmit_counter_2__bdd_4_lut_54495.LUT_INIT = 16'he4aa;
    SB_LUT4 n70237_bdd_4_lut (.I0(n70237), .I1(n63732), .I2(n63731), .I3(byte_transmit_counter[3]), 
            .O(n70240));
    defparam n70237_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54510 (.I0(byte_transmit_counter[1]), 
            .I1(n63746), .I2(n63747), .I3(\byte_transmit_counter[2] ), 
            .O(n70231));
    defparam byte_transmit_counter_1__bdd_4_lut_54510.LUT_INIT = 16'he4aa;
    SB_LUT4 n70231_bdd_4_lut (.I0(n70231), .I1(n63837), .I2(n63836), .I3(\byte_transmit_counter[2] ), 
            .O(n70234));
    defparam n70231_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1700 (.I0(n52766), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[17] [2]), 
            .O(n58259));
    defparam i2_3_lut_4_lut_adj_1700.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_215_i3_4_lut (.I0(n58108), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58293), .I3(\data_out_frame[25] [0]), .O(n3_adj_5557));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_215_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 n70477_bdd_4_lut (.I0(n70477), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n70480));
    defparam n70477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1701 (.I0(\data_out_frame[24] [5]), .I1(n23704), 
            .I2(GND_net), .I3(GND_net), .O(n58108));
    defparam i1_2_lut_adj_1701.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54486 (.I0(byte_transmit_counter[1]), 
            .I1(n63896), .I2(n63897), .I3(\byte_transmit_counter[2] ), 
            .O(n70225));
    defparam byte_transmit_counter_1__bdd_4_lut_54486.LUT_INIT = 16'he4aa;
    SB_LUT4 n70225_bdd_4_lut (.I0(n70225), .I1(n63651), .I2(n63650), .I3(\byte_transmit_counter[2] ), 
            .O(n70228));
    defparam n70225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54500 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n70219));
    defparam byte_transmit_counter_0__bdd_4_lut_54500.LUT_INIT = 16'he4aa;
    SB_LUT4 n70219_bdd_4_lut (.I0(n70219), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n70222));
    defparam n70219_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_780_Select_214_i3_4_lut (.I0(n53789), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58108), .I3(\data_out_frame[24] [4]), .O(n3_adj_5556));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_214_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54476 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n70213));
    defparam byte_transmit_counter_0__bdd_4_lut_54476.LUT_INIT = 16'he4aa;
    SB_LUT4 n70213_bdd_4_lut (.I0(n70213), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n70216));
    defparam n70213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1702 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58442));
    defparam i1_2_lut_adj_1702.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1703 (.I0(\data_out_frame[22] [3]), .I1(n58387), 
            .I2(GND_net), .I3(GND_net), .O(n53789));
    defparam i1_2_lut_adj_1703.LUT_INIT = 16'h6666;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(n63851), 
            .I2(n63852), .I3(r_Bit_Index[1]), .O(n70207));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70207_bdd_4_lut (.I0(n70207), .I1(n63849), .I2(n63848), .I3(r_Bit_Index[1]), 
            .O(n70210));
    defparam n70207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54692 (.I0(byte_transmit_counter[3]), 
            .I1(n70138), .I2(n66439), .I3(byte_transmit_counter[4]), .O(n70471));
    defparam byte_transmit_counter_3__bdd_4_lut_54692.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1704 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[8] [3]), .O(n58025));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1704.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5480));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54471 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n70201));
    defparam byte_transmit_counter_0__bdd_4_lut_54471.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1705 (.I0(\data_out_frame[19] [3]), .I1(n26771), 
            .I2(n58259), .I3(n58186), .O(n53855));
    defparam i1_2_lut_4_lut_adj_1705.LUT_INIT = 16'h6996;
    SB_LUT4 n70201_bdd_4_lut (.I0(n70201), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n70204));
    defparam n70201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n70471_bdd_4_lut (.I0(n70471), .I1(n70264), .I2(n7_adj_5596), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n70471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54682 (.I0(byte_transmit_counter[3]), 
            .I1(n70144), .I2(n66457), .I3(byte_transmit_counter[4]), .O(n70465));
    defparam byte_transmit_counter_3__bdd_4_lut_54682.LUT_INIT = 16'he4aa;
    SB_LUT4 n70465_bdd_4_lut (.I0(n70465), .I1(n70234), .I2(n7_adj_5595), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n70465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54462 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n70195));
    defparam byte_transmit_counter_0__bdd_4_lut_54462.LUT_INIT = 16'he4aa;
    SB_LUT4 n70195_bdd_4_lut (.I0(n70195), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n70198));
    defparam n70195_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_780_Select_213_i3_4_lut (.I0(n53789), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58442), .I3(n53818), .O(n3_adj_5555));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_213_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_3_lut_adj_1706 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(n52801), .I3(GND_net), .O(n58253));
    defparam i1_2_lut_3_lut_adj_1706.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5479));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i21004_3_lut (.I0(control_mode_c[3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n22773), .I3(GND_net), .O(n29647));
    defparam i21004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20997_3_lut (.I0(control_mode_c[2]), .I1(\data_in_frame[1][2] ), 
            .I2(n22773), .I3(GND_net), .O(n29648));
    defparam i20997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21468_3_lut (.I0(\control_mode[1] ), .I1(\data_in_frame[1]_c [1]), 
            .I2(n22773), .I3(GND_net), .O(n29649));
    defparam i21468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_780_Select_212_i3_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n58381), .I3(\data_out_frame[24] [3]), 
            .O(n3_adj_5554));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_212_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1707 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58281));
    defparam i1_2_lut_adj_1707.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54687 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n70459));
    defparam byte_transmit_counter_0__bdd_4_lut_54687.LUT_INIT = 16'he4aa;
    SB_LUT4 select_780_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1708 (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[19] [6]), 
            .I2(n53125), .I3(GND_net), .O(n53746));
    defparam i1_2_lut_3_lut_adj_1708.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_780_Select_211_i3_4_lut (.I0(n23700), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58281), .I3(n25145), .O(n3_adj_5553));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_211_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_4_lut_adj_1709 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(n58651), .I3(n53757), .O(n53258));
    defparam i2_3_lut_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 n70459_bdd_4_lut (.I0(n70459), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n70462));
    defparam n70459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1710 (.I0(n58445), .I1(n53855), .I2(\data_out_frame[24] [1]), 
            .I3(\data_out_frame[23] [6]), .O(n12_adj_5647));
    defparam i5_4_lut_adj_1710.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_210_i3_4_lut (.I0(n53361), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5647), .I3(n8_adj_5581), .O(n3_adj_5552));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1711 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n57922));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1711.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1712 (.I0(n53746), .I1(n58757), .I2(GND_net), 
            .I3(GND_net), .O(n58445));
    defparam i1_2_lut_adj_1712.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1713 (.I0(n52546), .I1(\data_out_frame[18] [3]), 
            .I2(n53831), .I3(GND_net), .O(n53875));
    defparam i2_3_lut_adj_1713.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1714 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[11] [5]), 
            .I2(n52569), .I3(n26402), .O(n58373));
    defparam i1_2_lut_4_lut_adj_1714.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54457 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n70177));
    defparam byte_transmit_counter_0__bdd_4_lut_54457.LUT_INIT = 16'he4aa;
    SB_LUT4 n70177_bdd_4_lut (.I0(n70177), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n70180));
    defparam n70177_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1715 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[13] [7]), .I3(n52861), .O(n58687));
    defparam i1_2_lut_4_lut_adj_1715.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54443 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n70171));
    defparam byte_transmit_counter_0__bdd_4_lut_54443.LUT_INIT = 16'he4aa;
    SB_LUT4 n70171_bdd_4_lut (.I0(n70171), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n70174));
    defparam n70171_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1716 (.I0(\data_out_frame[23] [5]), .I1(n52790), 
            .I2(n53361), .I3(GND_net), .O(n26382));
    defparam i1_2_lut_3_lut_adj_1716.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1717 (.I0(n58562), .I1(n53195), .I2(n58183), 
            .I3(GND_net), .O(n58644));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1717.LUT_INIT = 16'h9696;
    SB_LUT4 select_780_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1718 (.I0(n58313), .I1(\data_out_frame[16] [3]), 
            .I2(n60912), .I3(GND_net), .O(n60828));
    defparam i2_3_lut_adj_1718.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54677 (.I0(byte_transmit_counter[3]), 
            .I1(n70162), .I2(n66234), .I3(byte_transmit_counter[4]), .O(n70453));
    defparam byte_transmit_counter_3__bdd_4_lut_54677.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54481 (.I0(byte_transmit_counter[1]), 
            .I1(n63872), .I2(n63873), .I3(\byte_transmit_counter[2] ), 
            .O(n70165));
    defparam byte_transmit_counter_1__bdd_4_lut_54481.LUT_INIT = 16'he4aa;
    SB_LUT4 n70165_bdd_4_lut (.I0(n70165), .I1(n63786), .I2(n63785), .I3(\byte_transmit_counter[2] ), 
            .O(n70168));
    defparam n70165_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54434 (.I0(byte_transmit_counter[1]), 
            .I1(n63818), .I2(n63819), .I3(\byte_transmit_counter[2] ), 
            .O(n70159));
    defparam byte_transmit_counter_1__bdd_4_lut_54434.LUT_INIT = 16'he4aa;
    SB_LUT4 n70159_bdd_4_lut (.I0(n70159), .I1(n63813), .I2(n63812), .I3(\byte_transmit_counter[2] ), 
            .O(n70162));
    defparam n70159_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54429 (.I0(byte_transmit_counter[1]), 
            .I1(n63809), .I2(n63810), .I3(\byte_transmit_counter[2] ), 
            .O(n70153));
    defparam byte_transmit_counter_1__bdd_4_lut_54429.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1719 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(n58355), .I3(n53723), .O(n23704));
    defparam i2_3_lut_4_lut_adj_1719.LUT_INIT = 16'h9669;
    SB_LUT4 n70153_bdd_4_lut (.I0(n70153), .I1(n63825), .I2(n63824), .I3(\byte_transmit_counter[2] ), 
            .O(n70156));
    defparam n70153_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i17_4_lut_adj_1720 (.I0(n58465), .I1(n58595), .I2(\data_out_frame[12] [0]), 
            .I3(n58135), .O(n42_adj_5648));   // verilog/coms.v(88[17:63])
    defparam i17_4_lut_adj_1720.LUT_INIT = 16'h6996;
    SB_LUT4 n70453_bdd_4_lut (.I0(n70453), .I1(n14_adj_5527), .I2(n7_adj_5594), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n70453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15_4_lut_adj_1721 (.I0(\data_out_frame[5] [2]), .I1(n58702), 
            .I2(n53871), .I3(n58468), .O(n40_adj_5649));   // verilog/coms.v(88[17:63])
    defparam i15_4_lut_adj_1721.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_1722 (.I0(n58046), .I1(n1244), .I2(n1668), .I3(\data_out_frame[13] [7]), 
            .O(n41_adj_5650));   // verilog/coms.v(88[17:63])
    defparam i16_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54424 (.I0(byte_transmit_counter[1]), 
            .I1(n63770), .I2(n63771), .I3(\byte_transmit_counter[2] ), 
            .O(n70147));
    defparam byte_transmit_counter_1__bdd_4_lut_54424.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54672 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n70447));
    defparam byte_transmit_counter_0__bdd_4_lut_54672.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1723 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n58099));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1723.LUT_INIT = 16'h9696;
    SB_LUT4 n70147_bdd_4_lut (.I0(n70147), .I1(n63834), .I2(n63833), .I3(\byte_transmit_counter[2] ), 
            .O(n70150));
    defparam n70147_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n24));   // verilog/coms.v(100[12:26])
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut_adj_1724 (.I0(\data_out_frame[4] [0]), .I1(n1668), 
            .I2(n58025), .I3(\data_out_frame[5] [4]), .O(n39_adj_5651));   // verilog/coms.v(88[17:63])
    defparam i14_4_lut_adj_1724.LUT_INIT = 16'h6996;
    SB_LUT4 i13_3_lut (.I0(n53765), .I1(\data_out_frame[14] [1]), .I2(n58609), 
            .I3(GND_net), .O(n38_adj_5652));   // verilog/coms.v(88[17:63])
    defparam i13_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i12_2_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/coms.v(88[17:63])
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i23_4_lut (.I0(n39_adj_5651), .I1(n41_adj_5650), .I2(n40_adj_5649), 
            .I3(n42_adj_5648), .O(n48));   // verilog/coms.v(88[17:63])
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1725 (.I0(n52569), .I1(n58487), .I2(n58696), 
            .I3(n58262), .O(n43_adj_5653));   // verilog/coms.v(88[17:63])
    defparam i18_4_lut_adj_1725.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1726 (.I0(n43_adj_5653), .I1(n48), .I2(n37), 
            .I3(n38_adj_5652), .O(n60912));   // verilog/coms.v(88[17:63])
    defparam i24_4_lut_adj_1726.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1727 (.I0(n60912), .I1(n26704), .I2(n26402), 
            .I3(n1699), .O(n58363));
    defparam i3_4_lut_adj_1727.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54419 (.I0(byte_transmit_counter[1]), 
            .I1(n63656), .I2(n63657), .I3(\byte_transmit_counter[2] ), 
            .O(n70141));
    defparam byte_transmit_counter_1__bdd_4_lut_54419.LUT_INIT = 16'he4aa;
    SB_LUT4 n70447_bdd_4_lut (.I0(n70447), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n70450));
    defparam n70447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1728 (.I0(\data_out_frame[11] [5]), .I1(n52569), 
            .I2(n26402), .I3(GND_net), .O(n58372));
    defparam i1_2_lut_3_lut_adj_1728.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1729 (.I0(\data_out_frame[11] [5]), .I1(n52569), 
            .I2(n26794), .I3(n26704), .O(n52861));
    defparam i2_3_lut_4_lut_adj_1729.LUT_INIT = 16'h6996;
    SB_LUT4 n70141_bdd_4_lut (.I0(n70141), .I1(n63843), .I2(n63842), .I3(\byte_transmit_counter[2] ), 
            .O(n70144));
    defparam n70141_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1730 (.I0(n52877), .I1(n58363), .I2(n26111), 
            .I3(GND_net), .O(n52546));
    defparam i2_3_lut_adj_1730.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1731 (.I0(\data_out_frame[16] [2]), .I1(n58363), 
            .I2(n60828), .I3(GND_net), .O(n53853));
    defparam i2_3_lut_adj_1731.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54414 (.I0(byte_transmit_counter[1]), 
            .I1(n63728), .I2(n63729), .I3(\byte_transmit_counter[2] ), 
            .O(n70135));
    defparam byte_transmit_counter_1__bdd_4_lut_54414.LUT_INIT = 16'he4aa;
    SB_LUT4 n70135_bdd_4_lut (.I0(n70135), .I1(n63654), .I2(n63653), .I3(\byte_transmit_counter[2] ), 
            .O(n70138));
    defparam n70135_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54409 (.I0(byte_transmit_counter[1]), 
            .I1(n63800), .I2(n63801), .I3(\byte_transmit_counter[2] ), 
            .O(n70129));
    defparam byte_transmit_counter_1__bdd_4_lut_54409.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1732 (.I0(\data_out_frame[16] [6]), .I1(n26872), 
            .I2(n26771), .I3(GND_net), .O(n25733));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1732.LUT_INIT = 16'h9696;
    SB_LUT4 n70129_bdd_4_lut (.I0(n70129), .I1(n63795), .I2(n63794), .I3(\byte_transmit_counter[2] ), 
            .O(n70132));
    defparam n70129_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1733 (.I0(\data_out_frame[18] [4]), .I1(n53853), 
            .I2(GND_net), .I3(GND_net), .O(n58357));
    defparam i1_2_lut_adj_1733.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1734 (.I0(n53853), .I1(n52546), .I2(n25819), 
            .I3(GND_net), .O(n59809));
    defparam i2_3_lut_adj_1734.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1735 (.I0(n58534), .I1(n25082), .I2(\data_out_frame[13] [5]), 
            .I3(n58669), .O(n10_adj_5543));
    defparam i4_4_lut_adj_1735.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1736 (.I0(n26771), .I1(n58259), .I2(n58186), 
            .I3(GND_net), .O(n58763));
    defparam i1_2_lut_3_lut_adj_1736.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1737 (.I0(n26771), .I1(n58259), .I2(n52896), 
            .I3(\data_out_frame[19] [4]), .O(n52883));
    defparam i1_3_lut_4_lut_adj_1737.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54404 (.I0(byte_transmit_counter[1]), 
            .I1(n63899), .I2(n63900), .I3(\byte_transmit_counter[2] ), 
            .O(n70123));
    defparam byte_transmit_counter_1__bdd_4_lut_54404.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_adj_1738 (.I0(\data_out_frame[18] [0]), .I1(n10_adj_5543), 
            .I2(\data_out_frame[16] [0]), .I3(GND_net), .O(n52799));
    defparam i5_3_lut_adj_1738.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1739 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26405));
    defparam i1_2_lut_adj_1739.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1740 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25819));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1740.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1741 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[17] [5]), .I3(n69296), .O(n14_adj_5654));
    defparam i6_4_lut_adj_1741.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1742 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[17] [7]), .I3(\data_out_frame[17] [1]), 
            .O(n13));
    defparam i5_4_lut_adj_1742.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1743 (.I0(\data_out_frame[17] [6]), .I1(n26872), 
            .I2(n13), .I3(n14_adj_5654), .O(n8_adj_5655));
    defparam i3_4_lut_adj_1743.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1744 (.I0(\data_out_frame[20] [4]), .I1(n53875), 
            .I2(\data_out_frame[20] [5]), .I3(\data_out_frame[20] [6]), 
            .O(n6_adj_5263));
    defparam i1_2_lut_4_lut_adj_1744.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1745 (.I0(n58333), .I1(n26427), .I2(\data_out_frame[19] [6]), 
            .I3(n58633), .O(n15_adj_5656));
    defparam i6_4_lut_adj_1745.LUT_INIT = 16'h6996;
    SB_LUT4 i53574_4_lut (.I0(n52801), .I1(n60683), .I2(n8_adj_5655), 
            .I3(n58375), .O(n69300));
    defparam i53574_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1746 (.I0(n15_adj_5656), .I1(n58769), .I2(n14_adj_5632), 
            .I3(n58636), .O(n60931));
    defparam i8_4_lut_adj_1746.LUT_INIT = 16'h6996;
    SB_LUT4 select_780_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_780_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1747 (.I0(n58078), .I1(\data_in_frame[5] [5]), 
            .I2(n25915), .I3(n58607), .O(n58608));
    defparam i1_2_lut_4_lut_adj_1747.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1748 (.I0(\data_out_frame[19] [0]), .I1(n58582), 
            .I2(\data_out_frame[18] [6]), .I3(GND_net), .O(n58579));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1748.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1749 (.I0(n26280), .I1(n26122), .I2(\data_out_frame[17] [0]), 
            .I3(n26771), .O(n58205));
    defparam i3_4_lut_adj_1749.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1750 (.I0(n58205), .I1(n58579), .I2(\data_out_frame[16] [6]), 
            .I3(n58366), .O(n13_adj_5657));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1750.LUT_INIT = 16'h6996;
    SB_LUT4 n70123_bdd_4_lut (.I0(n70123), .I1(n63903), .I2(n63902), .I3(\byte_transmit_counter[2] ), 
            .O(n70126));
    defparam n70123_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i54395_1_lut (.I0(n3472), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70121));   // verilog/coms.v(148[4] 304[11])
    defparam i54395_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1751 (.I0(n13_adj_5657), .I1(n60828), .I2(n12_adj_5588), 
            .I3(n26875), .O(n53195));   // verilog/coms.v(88[17:28])
    defparam i7_4_lut_adj_1751.LUT_INIT = 16'h9669;
    uart_tx tx (.n462(n460[1]), .n59012(n59012), .r_Bit_Index({r_Bit_Index}), 
            .clk16MHz(clk16MHz), .n29148(n29148), .n461(n460[2]), .n44533(n44533), 
            .tx_o(tx_o), .tx_data({tx_data}), .n22192(n22192), .r_SM_Main({r_SM_Main}), 
            .GND_net(GND_net), .n85(n85), .n53949(n53949), .tx_active(tx_active), 
            .\r_SM_Main_2__N_3536[1] (\r_SM_Main_2__N_3536[1] ), .n59553(n59553), 
            .n58909(n58909), .r_Clock_Count({r_Clock_Count}), .n53963(n53963), 
            .VCC_net(VCC_net), .n63848(n63848), .n63849(n63849), .n63852(n63852), 
            .n63851(n63851), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n61386(n61386), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n29(n29), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .n23(n23), .n4942(n4942), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .baudrate({baudrate}), .VCC_net(VCC_net), 
            .n27845(n27845), .clk16MHz(clk16MHz), .n58988(n58988), .\r_SM_Main[2] (\r_SM_Main[2] ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .r_Clock_Count({r_Clock_Count_adj_23}), 
            .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), 
            .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n29(n29), .n23(n23), .n61478(n61478), .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), 
            .n27(n27), .\r_SM_Main[1] (\r_SM_Main[1] ), .n4939(n4939), 
            .n25566(n25566), .n29596(n29596), .rx_data({rx_data}), .n29595(n29595), 
            .n29591(n29591), .n29590(n29590), .n29559(n29559), .n29558(n29558), 
            .n29557(n29557), .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n61043(n61043), 
            .n30440(n30440), .n53943(n53943), .rx_data_ready(rx_data_ready), 
            .n30436(n30436), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n61750(n61750), .n61702(n61702), .n61734(n61734), .n61814(n61814), 
            .n61782(n61782), .n61766(n61766), .n61798(n61798), .n61718(n61718), 
            .n57927(n57927), .n27722(n27722)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n462, n59012, r_Bit_Index, clk16MHz, n29148, n461, 
            n44533, tx_o, tx_data, n22192, r_SM_Main, GND_net, n85, 
            n53949, tx_active, \r_SM_Main_2__N_3536[1] , n59553, n58909, 
            r_Clock_Count, n53963, VCC_net, n63848, n63849, n63852, 
            n63851, \r_SM_Main_2__N_3545[0] , n61386, \o_Rx_DV_N_3488[24] , 
            n27, n29, \o_Rx_DV_N_3488[12] , n23, n4942, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input n462;
    input n59012;
    output [2:0]r_Bit_Index;
    input clk16MHz;
    input n29148;
    input n461;
    input n44533;
    output tx_o;
    input [7:0]tx_data;
    input n22192;
    output [2:0]r_SM_Main;
    input GND_net;
    output n85;
    input n53949;
    output tx_active;
    input \r_SM_Main_2__N_3536[1] ;
    output n59553;
    output n58909;
    output [8:0]r_Clock_Count;
    input n53963;
    input VCC_net;
    output n63848;
    output n63849;
    output n63852;
    output n63851;
    input \r_SM_Main_2__N_3545[0] ;
    output n61386;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    input n29;
    input \o_Rx_DV_N_3488[12] ;
    input n23;
    input n4942;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n40063, n25022;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n3, n70506;
    wire [8:0]n41;
    
    wire n40035, n51704, n51703, n51702, n51701, n51700, n51699, 
        n51698, n51697, n14, n15, n61380;
    
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n59012), 
            .D(n462), .R(n29148));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n59012), 
            .D(n461), .R(n29148));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n40063), .D(n44533));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n22192), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40063));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_2_lut (.I0(n85), .I1(r_SM_Main[1]), .I2(GND_net), .I3(GND_net), 
            .O(n3));   // verilog/uart_tx.v(32[16:25])
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n53949));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n70506));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i43118_rep_31_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n59553));
    defparam i43118_rep_31_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i43236_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n58909));
    defparam i43236_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR r_Clock_Count_1954__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n40063), .D(n41[0]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n40063), .D(n41[1]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n40063), .D(n41[2]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n40063), .D(n41[3]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n40063), .D(n41[4]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n40063), .D(n41[5]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n40063), .D(n41[6]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n40063), .D(n41[7]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1954__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n40063), .D(n41[8]), .R(n40035));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n53963));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i48122_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63848));
    defparam i48122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48123_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63849));
    defparam i48123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48126_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63852));
    defparam i48126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48125_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63851));
    defparam i48125_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25022), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_1954_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n51704), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1954_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n51703), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_9 (.CI(n51703), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n51704));
    SB_LUT4 r_Clock_Count_1954_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n51702), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_8 (.CI(n51702), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n51703));
    SB_LUT4 r_Clock_Count_1954_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n51701), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_7 (.CI(n51701), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n51702));
    SB_LUT4 r_Clock_Count_1954_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n51700), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_6 (.CI(n51700), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n51701));
    SB_LUT4 r_Clock_Count_1954_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n51699), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_5 (.CI(n51699), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n51700));
    SB_LUT4 r_Clock_Count_1954_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n51698), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_4 (.CI(n51698), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n51699));
    SB_LUT4 r_Clock_Count_1954_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n51697), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_3 (.CI(n51697), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n51698));
    SB_LUT4 r_Clock_Count_1954_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1954_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1954_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n51697));
    SB_LUT4 i1_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n61386));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h3130;
    SB_LUT4 i54322_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n40035));
    defparam i54322_4_lut.LUT_INIT = 16'h1113;
    SB_LUT4 i2_3_lut_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n25022));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4942), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n40063), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n70506));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4942), 
            .I3(r_SM_Main[0]), .O(n61380));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n61380), .O(n85));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'h0100;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, baudrate, VCC_net, n27845, clk16MHz, n58988, 
            \r_SM_Main[2] , r_Rx_Data, RX_N_2, r_Clock_Count, \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[4] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , 
            n29, n23, n61478, \r_SM_Main_2__N_3446[1] , n27, \r_SM_Main[1] , 
            n4939, n25566, n29596, rx_data, n29595, n29591, n29590, 
            n29559, n29558, n29557, \r_Bit_Index[0] , n61043, n30440, 
            n53943, rx_data_ready, n30436, \o_Rx_DV_N_3488[0] , n61750, 
            n61702, n61734, n61814, n61782, n61766, n61798, n61718, 
            n57927, n27722) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [31:0]baudrate;
    input VCC_net;
    output n27845;
    input clk16MHz;
    output n58988;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_2;
    output [7:0]r_Clock_Count;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    input n61478;
    input \r_SM_Main_2__N_3446[1] ;
    output n27;
    output \r_SM_Main[1] ;
    input n4939;
    output n25566;
    input n29596;
    output [7:0]rx_data;
    input n29595;
    input n29591;
    input n29590;
    input n29559;
    input n29558;
    input n29557;
    output \r_Bit_Index[0] ;
    output n61043;
    input n30440;
    input n53943;
    output rx_data_ready;
    input n30436;
    output \o_Rx_DV_N_3488[0] ;
    output n61750;
    output n61702;
    output n61734;
    output n61814;
    output n61782;
    output n61766;
    output n61798;
    output n61718;
    input n57927;
    output n27722;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n8367;
    
    wire n2940, n2977, n51490, n58877, n63559, n62822, n42418, 
        n61930, n59605, n60615, n66329, n63557, n61984, n66330;
    wire [23:0]n8107;
    
    wire n1702, n858;
    wire [23:0]n294;
    
    wire n63322, n58832, n51424, n2607, n1459, n51425, n58834, 
        n803, n59595, n44, n46;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n51330, n58836, n62914, n62918, n62920, n62770, n62916, 
        n25654;
    wire [23:0]n8081;
    
    wire n1552, n1879, n51329, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire r_Rx_Data_R, n51491, n1553, n1742, n51328;
    wire [23:0]n8289;
    
    wire n2608, n1460, n51423, n2941, n2867, n51489, n2609, n1011, 
        n51422, n1554, n1602, n51327, n1555, n51326, n61850, n61842, 
        n61846, n61848, n63296, n63298, n61844, n63575, n2942, 
        n2754, n51488, n63601, n63475, n63635, n63639, n1556, 
        n51325, n1557, n51324, n2610, n856, n51421, n1558, n51323, 
        n2611, n698, n51420, n2943, n2638, n51487, n2612, n51419, 
        n1559, n51322, n2944, n2519, n51486, n61356, n538, n59078, 
        n1560, n51321, n2945, n2397, n51485;
    wire [23:0]n8263;
    
    wire n2476, n51418, n2477, n51417, n2946, n2272, n51484, n3066;
    wire [23:0]n8393;
    
    wire n3171, n2947, n2144, n51483;
    wire [23:0]n8055;
    
    wire n1408, n51320, n2948, n2013, n51482, n2478, n51416, n2479, 
        n51415, n1409, n51319, n1410, n51318, n2949, n51481, n3065, 
        n3170, n1411, n51317, n3064, n3169, n2480, n51414, n3063, 
        n3168, n2481, n51413, n3062, n3167, n1412, n51316, n2950, 
        n51480, n1413, n51315, n2951, n51479, n1414, n51314, n2482, 
        n51412, n1415, n51313, n61346, n59108, n2483, n51411, 
        n3061, n3166, n62404, n3_adj_4993, n2484, n51410;
    wire [23:0]n8419;
    
    wire n3151, n3186, n51536, n3152, n3082, n51535, n2485, n51409, 
        n2486, n51408, n62408, n5, n62412, n8, n57703, n63517, 
        n63621, n2, n2487, n51407, n3153, n3188, n51534, n3154, 
        n3084, n51533, n3155, n51532, n2952, n51478, n2488, n51406, 
        n11608, n2953, n51477, n2489, n51405;
    wire [23:0]n8029;
    
    wire n1261, n51307, n1262, n51306, n2490, n51404, n3156, n51531, 
        n2954, n51476, n1263, n51305, n2491, n51403, n2955, n51475, 
        n61354, n59082, n3157, n51530, n2956, n51474, n3158, n51529;
    wire [23:0]n8237;
    
    wire n2353, n51402, n2354, n51401, n3159, n51528, n2957, n51473, 
        n1264, n51304, n1265, n51303, n2355, n51400, n1266, n51302, 
        n61362, n59066, n3160, n51527, n1267, n51301, n2356, n51399;
    wire [23:0]n8341;
    
    wire n2827, n51472, n2828, n51471, n2829, n51470, n3161, n51526, 
        n3060, n3165, n66373, n66379, n61344, n59112, n3162, n51525;
    wire [23:0]n8003;
    
    wire n1111, n51300, n1112, n51299, n66370, n66376, n2830, 
        n51469, n3_adj_4994, n3163, n51524, n3059, n3164, n2831, 
        n51468, n1113, n51298, n51523, n2357, n51398, n2358, n51397, 
        n3058, n2359, n51396, n51522, n2832, n51467, n2360, n51395, 
        n1114, n51297, n1115, n51296, n2361, n51394, n2833, n51466, 
        n2834, n51465, n2362, n51393, n1116, n51295, n51521, n51520, 
        n61342, n59116, n51519, n51518, n3057, n3056, n3055, n2835, 
        n51464, n2836, n51463, n51517, n3054, n3053, n3052, n2837, 
        n51462, n51516, n50455, n50454, n61330, n2838, n51461, 
        n50453, n61418, n3051, n2363, n51392, n3172, n51515, n2364, 
        n51391, n2839, n51460, n2365, n51390, n50452;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n2840, n51459, n2366, n51389, n2367, n51388, n50451, 
        n61416, n50450, n61414, n61366, n51514, n59058, n61352, 
        n59086, n2841, n51458;
    wire [23:0]n8211;
    
    wire n2227, n51387, n2228, n51386, n2842, n51457, n2229, n51385, 
        n3050, n2230, n51384, n3049, n3048, n50449, n3046, n51513, 
        n50448, n61412, n63523, n2843, n51456, n50447, n61410, 
        n804, n20834, n20836, n3047, n51512, n2939, n2844, n51455, 
        n2231, n51383, n39, n50446, n61328, n19, n35, n33, n37, 
        n2232, n51382, n35_adj_4995, n27_adj_4996, n50445, n61408, 
        n29_adj_4997, n23_adj_4998, n21, n23_adj_4999, n25, n2845, 
        n51454, n51511, n2233, n51381, n2234, n51380, n11, n13, 
        n21_adj_5000, n61360, n59070, n50444, n17, n25_adj_5001, 
        n2728;
    wire [23:0]n8315;
    
    wire n2938, n37_adj_5002, n15, n41, n35_adj_5003, n39_adj_5004, 
        n23_adj_5005, n25_adj_5006, n27_adj_5007, n2235, n51379, n50443, 
        n29_adj_5008, n27_adj_5009, n50442, n2713, n51453, n51510, 
        n2236, n51378, n2714, n51452, n31, n45, n2237, n51377, 
        n29_adj_5010, n959, n59555, n44_adj_5011, n46_adj_5012, n31_adj_5013, 
        n37_adj_5014, n50441, n69211, n1831, n61348, n1977, n41_adj_5015, 
        n39_adj_5016, n35_adj_5017, n2716, n41_adj_5018, n2717, n39_adj_5019, 
        n37_adj_5020, n29_adj_5021, n2715, n43, n17_adj_5022, n2727, 
        n19_adj_5023, n2726, n21_adj_5024, n2725, n23_adj_5025, n39_adj_5026, 
        n31_adj_5027, n2724, n25_adj_5028, n2720, n33_adj_5029, n2719, 
        n35_adj_5030, n41_adj_5031, n23_adj_5032, n2718, n37_adj_5033, 
        n2723, n27_adj_5034, n63577, n25_adj_5035, n2238, n51376, 
        n33_adj_5036, n1699, n1700, n67155, n33_adj_5037, n7, n45_adj_5038, 
        n9, n2722, n29_adj_5039, n17_adj_5040, n19_adj_5041, n2721, 
        n31_adj_5042, n66902, n2729, n67806, n68371, n68367, n66904, 
        n2730, n14, n68817, n68818, n1693;
    wire [23:0]n8133;
    
    wire n1966;
    wire [23:0]n8159;
    
    wire n2098;
    wire [23:0]n8185;
    
    wire n2596, n34, n62724, n62726, n51451, n21_adj_5043, n2239, 
        n51375, n51509, n43_adj_5044, n11_adj_5045, n22, n40, n66897, 
        n20, n66895, n68391, n13_adj_5046, n15_adj_5047, n68714, 
        n27_adj_5048, n66622, n66640, n16, n66560, n18, n26, n16_adj_5049, 
        n66918, n69127, n69128, n8_adj_5050, n69021, n68665, n68965, 
        n68964, n68967, n24, n3274, n2601, n37_adj_5051, n2598, 
        n43_adj_5052, n2599, n41_adj_5053, n2600, n39_adj_5054, n70507, 
        n2240, n51374, n66656, n67540, n67534, n2604, n31_adj_5055, 
        n2603, n33_adj_5056, n2602, n35_adj_5057, n68861, n2606, 
        n27_adj_5058, n2605, n29_adj_5059, n51508, n50440, n68247, 
        n69076, n61350, n59090, n12, n19_adj_5060, n21_adj_5061, 
        n23_adj_5062, n48, n4, n25_adj_5063, n68787, n17_adj_5064, 
        n66990, n66983, n68697, n16_adj_5065, n68823, n51450, n68788, 
        n66602, n10, n50439, n51449, n30, n66608, n69139, n68824, 
        n66986, n67823, n22_adj_5066, n68389, n68707, n51507, n20_adj_5067, 
        n28, n18_adj_5068, n66967, n69125, n68746, n69256, n69126, 
        n69023, n67834, n68821, n68962, n69145, n69257, n6;
    wire [7:0]n1;
    
    wire n27766, n29073, n68789, n68790, n2597, n69146, n50438, 
        n51373, n2099, n51372, n66564, n13_adj_5075, n50437, n68401, 
        n68744, n50436, n15_adj_5076, n69201, n66569, n68982, n17_adj_5077, 
        n40_adj_5078, n61294, n3253, n19_adj_5079, n21_adj_5080, n33_adj_5081, 
        n63545, n62814, n63543, n62768, n66808, n63499, n61988, 
        n63617, n67724, n68984, n61664, n62772, n61302, n60390, 
        n33_adj_5082, n68331, n68329, n63563, n66813, n61692, n63483, 
        n63629, n66729, n69304, n37_adj_5083, n10_adj_5084, n68807, 
        n68808, n31_adj_5085, n44_adj_5086, n2100, n51371, n35_adj_5087, 
        n25_adj_5088, n27_adj_5089, n18_adj_5090, n36, n21_adj_5091, 
        n66802, n16_adj_5092, n66800, n69133, n68724, n14_adj_5093, 
        n22_adj_5094, n6_adj_5095, n12_adj_5096, n66822, n69131, n69132, 
        n23_adj_5097, n69015, n9_adj_5098, n1694, n51448, n68625, 
        n13_adj_5099, n69250, n15_adj_5100, n17_adj_5101, n68973, 
        n29_adj_5102, n69272, n69273, n69269, n2101, n51370, n25593, 
        n11_adj_5103, n19_adj_5104, n66680, n15_adj_5105, n17_adj_5106, 
        n19_adj_5107, n31_adj_5108, n66738, n67674, n67586, n68309, 
        n68281, n68277, n66682, n2102, n51369, n51506, n51447, 
        n6_adj_5109, n68795, n68305, n2103, n51368, n66742, n50435, 
        n50434, n8_adj_5110, n68801, n68802, n14_adj_5111, n32, 
        n68796, n66675, n16_adj_5112, n34_adj_5113, n12_adj_5114, 
        n66673, n69137, n66731, n14_adj_5115, n66722, n69135, n68730, 
        n10_adj_5116, n68803, n68804, n66753, n67654, n12_adj_5117, 
        n20_adj_5118, n26_adj_5119, n1832, n2104, n51367, n68736, 
        n68611, n69252, n8_adj_5120, n68797, n68798, n66692, n67566, 
        n68395, n69276, n10_adj_5121, n68399, n69277, n69265, n68734, 
        n68584, n68397, n50433, n51505, n51446, n2105, n51366, 
        n69254, n51504, n68791, n69274, n69275, n69267, n51445, 
        n69070, n69071, n2106, n51365, n51444, n2107, n51364, 
        n50432, n2108, n51363, n61364, n25651, n51503, n51443, 
        n63599, n2109, n51362, n1967, n20844, n11422, n960, n25639, 
        n2110, n51442, n51361, n62774, n61358, n1695, n43_adj_5122, 
        n1696, n41_adj_5123, n1697, n39_adj_5124, n1698, n37_adj_5125, 
        n59102, n1701, n32_adj_5126, n68574, n68575, n68014, n68685, 
        n67828, n25642, n68871, n68872, n48_adj_5127, n62800, n62802, 
        n62790, n25618, n1841, n1835, n39_adj_5128, n1836, n37_adj_5129, 
        n1833, n43_adj_5130, n1834, n41_adj_5131, n1837, n1838, 
        n1839, n31_adj_5132, n33_adj_5133, n35_adj_5134, n1840, n29_adj_5135, 
        n67137, n32_adj_5136, n40_adj_5137, n28_adj_5138, n68572, 
        n68573, n67131, n30_adj_5139, n67129, n69028, n67833, n69210, 
        n42_adj_5140, n20846, n51360, n51502, n42_adj_5141, n51441, 
        n1968, n51359, n1969, n51358, n1970, n51357, n51440, n51501, 
        n51439, n1971, n51356, n1972, n51355, n1973, n51354, n51438, 
        n1974, n51353, n69259, n1975, n51352, n25645, n61852, 
        n63605, n48_adj_5142, n962, n51500, n51437, n1976, n51351, 
        n51499, n51436, n51350, n51498, n51349, n59074, n51348, 
        n51347, n51435, n51497, n51346, n51434, n4_adj_5143, n51345, 
        n51496, n51344, n51433, n51343, n48_adj_5144, n63391, n48_adj_5145, 
        n62828, n61320, n61318, n62818, n51342, n39_adj_5146, n45_adj_5147, 
        n51432, n43_adj_5148, n41_adj_5149, n51341, n29_adj_5150, 
        n31_adj_5151, n21_adj_5152, n23_adj_5153, n42420, n51696, 
        n51695, n51694, n25_adj_5154, n27_adj_5155, n51431, n51340, 
        n33_adj_5156, n35_adj_5157, n51693, n51339, n51430, n59099, 
        n51338, n51337, n51429, n51495, n51428, n51494, n51336, 
        n37_adj_5158, n19_adj_5159, n67029, n51335, n51427, n67023, 
        n68753, n18_adj_5160, n51334, n51692, n51333, n51493, n51426, 
        n51332, n68543, n68544, n67025, n67892, n24_adj_5161, n26_adj_5162, 
        n59062, n67873, n51691, n51331, n51690, n22_adj_5163, n30_adj_5164, 
        n20_adj_5165, n67019, n69060, n69061, n51492, n68854, n67894, 
        n68701, n67871, n68703, n41_adj_5166, n39_adj_5167, n37_adj_5168, 
        n66733, n35_adj_5169, n48_adj_5170, n29_adj_5171, n31_adj_5172, 
        n33_adj_5173, n23_adj_5174, n25_adj_5175, n27_adj_5176, n21_adj_5177, 
        n67051, n67047, n20_adj_5178, n26_adj_5179, n28_adj_5180, 
        n43_adj_5181, n24_adj_5182, n32_adj_5183, n22_adj_5184, n67045, 
        n69058, n62012, n69059, n68856, n62820, n66858, n68757, 
        n67049, n69123, n67865, n69208, n69209, n69188, n67773, 
        n43_adj_5185, n62730, n68351, n62728, n68349, n43_adj_5186, 
        n39_adj_5187, n41_adj_5188, n37_adj_5189, n25_adj_5190, n14_adj_5191, 
        n37_adj_5192, n66878, n27_adj_5193, n16_adj_5194, n29_adj_5195, 
        n41_adj_5196, n31_adj_5197, n33_adj_5198, n35_adj_5199, n23_adj_5200, 
        n67078, n67074, n22_adj_5201, n28_adj_5202, n30_adj_5203, 
        n39_adj_5204, n26_adj_5205, n34_adj_5206, n24_adj_5207, n67072, 
        n69056, n69057, n68858, n68759, n67076, n68953, n67859, 
        n69026, n69027, n45_adj_5208, n39_adj_5209, n43_adj_5210, 
        n63361, n62710, n41_adj_5211, n18_adj_5212, n66848, n34_adj_5213, 
        n20_adj_5214, n68580, n68581, n67173, n68032, n36_adj_5215, 
        n38_adj_5216, n67817, n68677, n41_adj_5217, n961, n40_adj_5218, 
        n43_adj_5219, n28_adj_5220, n61870, n67107, n30_adj_5221, 
        n37_adj_5222, n35_adj_5223, n41_adj_5224, n39_adj_5225, n29_adj_5226, 
        n31_adj_5227, n33_adj_5228, n27_adj_5229, n67096, n30_adj_5230, 
        n38_adj_5231, n59093, n26_adj_5232, n68566, n68567, n67090, 
        n62700, n61890, n28_adj_5233, n67088, n69054, n62816, n67849, 
        n69220, n69221, n69156, n48_adj_5234, n62824, n62832, n38_adj_5235, 
        n62830, n25627, n40_adj_5236, n42_adj_5237, n67186, n69030, 
        n66393, n69031, n805, n59119, n42_adj_5238, n68588, n68589, 
        n48_adj_5239, n25603, n36_adj_5240, n38_adj_5241, n40_adj_5242, 
        n67179, n69050, n69051, n68880, n66862, n32_adj_5243, n68578, 
        n68579, n67165, n68026, n34_adj_5244, n68683, n37_adj_5245, 
        n35_adj_5246, n41_adj_5247, n67821, n39_adj_5248, n29_adj_5249, 
        n68875, n68876, n31_adj_5250, n33_adj_5251, n27_adj_5252, 
        n67117, n38_adj_5253, n26_adj_5254, n68570, n68571, n67109, 
        n69052, n67837, n69218, n69219, n69160, n66243, n66240, 
        n66301, n66298, n66295, n61432, n61438, n46_adj_5255, n12_adj_5256, 
        n48_adj_5257, n68813, n25597, n61996, n63603, n38_adj_5258, 
        n68814, n14_adj_5259, n15_adj_5260, n66850, n68811, n68718, 
        n24_adj_5261, n42_adj_5262, n68592, n68593, n69129, n69130, 
        n69017, n68651, n69181, n68971, n69258, n63569, n61282, 
        n61608, n61626, n63631, n61864, n61866;
    
    SB_LUT4 add_2797_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n51490), 
            .O(n8367[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i43206_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n58877));
    defparam i43206_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(n63559), .I1(n62822), .I2(baudrate[16]), .I3(n42418), 
            .O(n61930));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i51714_3_lut (.I0(n59605), .I1(n60615), .I2(baudrate[2]), 
            .I3(GND_net), .O(n66329));   // verilog/uart_rx.v(119[33:55])
    defparam i51714_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i51591_4_lut (.I0(n58877), .I1(n61930), .I2(n63557), .I3(n61984), 
            .O(n66330));   // verilog/uart_rx.v(119[33:55])
    defparam i51591_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 add_2787_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8107[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i427_4_lut (.I0(n66330), .I1(n66329), .I2(n294[21]), 
            .I3(n63322), .O(n58832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_CARRY add_2794_8 (.CI(n51424), .I0(n2607), .I1(n1459), .CO(n51425));
    SB_LUT4 div_37_i534_3_lut (.I0(n58832), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n58834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i5589_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n59595), .I3(n44), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i5589_4_lut.LUT_INIT = 16'hb3a0;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27845), 
            .D(n479[1]), .R(n58988));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2787_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n51330));
    SB_LUT4 div_37_i639_4_lut (.I0(n58834), .I1(n294[19]), .I2(n46), .I3(baudrate[4]), 
            .O(n58836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 i1_2_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n62914));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_968 (.I0(n62918), .I1(n62920), .I2(n62770), .I3(n62916), 
            .O(n25654));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'hfffe;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27845), 
            .D(n479[2]), .R(n58988));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2786_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n51329), 
            .O(n8081[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2797_20 (.CI(n51490), .I0(n2940), .I1(n2977), .CO(n51491));
    SB_LUT4 add_2786_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n51328), 
            .O(n8081[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n51423), 
            .O(n8289[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_7 (.CI(n51423), .I0(n2608), .I1(n1460), .CO(n51424));
    SB_LUT4 add_2797_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n51489), 
            .O(n8367[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_19 (.CI(n51489), .I0(n2941), .I1(n2867), .CO(n51490));
    SB_CARRY add_2786_10 (.CI(n51328), .I0(n1553), .I1(n1742), .CO(n51329));
    SB_LUT4 add_2794_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n51422), 
            .O(n8289[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2786_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n51327), 
            .O(n8081[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_9 (.CI(n51327), .I0(n1554), .I1(n1602), .CO(n51328));
    SB_LUT4 add_2786_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n51326), 
            .O(n8081[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_8 (.CI(n51326), .I0(n1555), .I1(n1459), .CO(n51327));
    SB_LUT4 i1_2_lut_adj_969 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n61850));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_970 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n61842));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_971 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n61846));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_972 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n61848));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'heeee;
    SB_LUT4 i47587_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n63296));
    defparam i47587_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_973 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n63298));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'heeee;
    SB_LUT4 i47858_4_lut (.I0(n61848), .I1(n61844), .I2(n61846), .I3(n61842), 
            .O(n63575));
    defparam i47858_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2797_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n51488), 
            .O(n8367[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47918_4_lut (.I0(n63601), .I1(n63475), .I2(n58877), .I3(baudrate[4]), 
            .O(n63635));
    defparam i47918_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53594_4_lut (.I0(n63575), .I1(n63298), .I2(n63635), .I3(n63296), 
            .O(n63639));
    defparam i53594_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY add_2794_6 (.CI(n51422), .I0(n2609), .I1(n1011), .CO(n51423));
    SB_LUT4 add_2786_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n51325), 
            .O(n8081[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_7 (.CI(n51325), .I0(n1556), .I1(n1460), .CO(n51326));
    SB_LUT4 add_2786_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n51324), 
            .O(n8081[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_6 (.CI(n51324), .I0(n1557), .I1(n1011), .CO(n51325));
    SB_CARRY add_2797_18 (.CI(n51488), .I0(n2942), .I1(n2754), .CO(n51489));
    SB_LUT4 add_2794_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n51421), 
            .O(n8289[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2786_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n51323), 
            .O(n8081[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_5 (.CI(n51421), .I0(n2610), .I1(n856), .CO(n51422));
    SB_LUT4 add_2794_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n51420), 
            .O(n8289[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_4 (.CI(n51420), .I0(n2611), .I1(n698), .CO(n51421));
    SB_LUT4 add_2797_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n51487), 
            .O(n8367[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_17 (.CI(n51487), .I0(n2943), .I1(n2638), .CO(n51488));
    SB_LUT4 add_2794_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n51419), 
            .O(n8289[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_5 (.CI(n51323), .I0(n1558), .I1(n856), .CO(n51324));
    SB_CARRY add_2794_3 (.CI(n51419), .I0(n2612), .I1(n858), .CO(n51420));
    SB_LUT4 add_2786_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n51322), 
            .O(n8081[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n51486), 
            .O(n8367[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_16 (.CI(n51486), .I0(n2944), .I1(n2519), .CO(n51487));
    SB_LUT4 add_2794_2_lut (.I0(n59078), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61356)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2794_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51419));
    SB_CARRY add_2786_4 (.CI(n51322), .I0(n1559), .I1(n698), .CO(n51323));
    SB_LUT4 add_2786_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n51321), 
            .O(n8081[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n51485), 
            .O(n8367[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n51418), 
            .O(n8263[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n51417), 
            .O(n8263[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_15 (.CI(n51485), .I0(n2945), .I1(n2397), .CO(n51486));
    SB_LUT4 add_2797_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n51484), 
            .O(n8367[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_3 (.CI(n51321), .I0(n1560), .I1(n858), .CO(n51322));
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8393[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2786_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8081[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_14 (.CI(n51484), .I0(n2946), .I1(n2272), .CO(n51485));
    SB_LUT4 add_2797_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n51483), 
            .O(n8367[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_13 (.CI(n51483), .I0(n2947), .I1(n2144), .CO(n51484));
    SB_CARRY add_2793_17 (.CI(n51417), .I0(n2477), .I1(n2638), .CO(n51418));
    SB_CARRY add_2786_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51321));
    SB_LUT4 add_2785_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n51320), 
            .O(n8055[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n51482), 
            .O(n8367[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n51416), 
            .O(n8263[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_16 (.CI(n51416), .I0(n2478), .I1(n2519), .CO(n51417));
    SB_CARRY add_2797_12 (.CI(n51482), .I0(n2948), .I1(n2013), .CO(n51483));
    SB_LUT4 add_2793_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n51415), 
            .O(n8263[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_15 (.CI(n51415), .I0(n2479), .I1(n2397), .CO(n51416));
    SB_LUT4 add_2785_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n51319), 
            .O(n8055[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_9 (.CI(n51319), .I0(n1409), .I1(n1602), .CO(n51320));
    SB_LUT4 add_2785_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n51318), 
            .O(n8055[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_8 (.CI(n51318), .I0(n1410), .I1(n1459), .CO(n51319));
    SB_LUT4 add_2797_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n51481), 
            .O(n8367[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8393[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2785_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n51317), 
            .O(n8055[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8393[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2793_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n51414), 
            .O(n8263[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8393[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2785_7 (.CI(n51317), .I0(n1411), .I1(n1460), .CO(n51318));
    SB_CARRY add_2797_11 (.CI(n51481), .I0(n2949), .I1(n1879), .CO(n51482));
    SB_CARRY add_2793_14 (.CI(n51414), .I0(n2480), .I1(n2272), .CO(n51415));
    SB_LUT4 add_2793_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n51413), 
            .O(n8263[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8393[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2785_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n51316), 
            .O(n8055[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_6 (.CI(n51316), .I0(n1412), .I1(n1011), .CO(n51317));
    SB_LUT4 add_2797_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n51480), 
            .O(n8367[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2785_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n51315), 
            .O(n8055[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_10 (.CI(n51480), .I0(n2950), .I1(n1742), .CO(n51481));
    SB_CARRY add_2793_13 (.CI(n51413), .I0(n2481), .I1(n2144), .CO(n51414));
    SB_CARRY add_2785_5 (.CI(n51315), .I0(n1413), .I1(n856), .CO(n51316));
    SB_LUT4 add_2797_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n51479), 
            .O(n8367[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2785_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n51314), 
            .O(n8055[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n51412), 
            .O(n8263[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_4 (.CI(n51314), .I0(n1414), .I1(n698), .CO(n51315));
    SB_LUT4 add_2785_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n51313), 
            .O(n8055[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_12 (.CI(n51412), .I0(n2482), .I1(n2013), .CO(n51413));
    SB_CARRY add_2785_3 (.CI(n51313), .I0(n1415), .I1(n858), .CO(n51314));
    SB_LUT4 add_2785_2_lut (.I0(n59108), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61346)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2785_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2793_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n51411), 
            .O(n8263[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2785_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51313));
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8393[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2797_9 (.CI(n51479), .I0(n2951), .I1(n1602), .CO(n51480));
    SB_LUT4 i1_4_lut_adj_974 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n62404));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_974.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_268_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4993));   // verilog/uart_rx.v(69[17:62])
    defparam equal_268_i3_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2793_11 (.CI(n51411), .I0(n2483), .I1(n1879), .CO(n51412));
    SB_LUT4 add_2793_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n51410), 
            .O(n8263[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_10 (.CI(n51410), .I0(n2484), .I1(n1742), .CO(n51411));
    SB_LUT4 add_2799_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n51536), 
            .O(n8419[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n51535), 
            .O(n8419[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n51409), 
            .O(n8263[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_9 (.CI(n51409), .I0(n2485), .I1(n1602), .CO(n51410));
    SB_LUT4 add_2793_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n51408), 
            .O(n8263[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_975 (.I0(r_Clock_Count[3]), .I1(n3_adj_4993), .I2(\o_Rx_DV_N_3488[4] ), 
            .I3(n62404), .O(n62408));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_975.LUT_INIT = 16'hffde;
    SB_LUT4 equal_268_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_268_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_976 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n62408), .O(n62412));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_976.LUT_INIT = 16'hffde;
    SB_CARRY add_2793_8 (.CI(n51408), .I0(n2486), .I1(n1459), .CO(n51409));
    SB_LUT4 equal_268_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(69[17:62])
    defparam equal_268_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_977 (.I0(r_Clock_Count[6]), .I1(n8), .I2(n62412), 
            .I3(\o_Rx_DV_N_3488[7] ), .O(n57703));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_977.LUT_INIT = 16'hfdfe;
    SB_LUT4 i47800_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n57703), .I2(GND_net), 
            .I3(GND_net), .O(n63517));
    defparam i47800_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47904_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n63517), .O(n63621));
    defparam i47904_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n61478), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 add_2793_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n51407), 
            .O(n8263[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_24 (.CI(n51535), .I0(n3152), .I1(n3082), .CO(n51536));
    SB_LUT4 add_2799_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n51534), 
            .O(n8419[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_23 (.CI(n51534), .I0(n3153), .I1(n3188), .CO(n51535));
    SB_LUT4 add_2799_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n51533), 
            .O(n8419[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_22 (.CI(n51533), .I0(n3154), .I1(n3084), .CO(n51534));
    SB_LUT4 add_2799_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n51532), 
            .O(n8419[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_7 (.CI(n51407), .I0(n2487), .I1(n1460), .CO(n51408));
    SB_LUT4 add_2797_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n51478), 
            .O(n8367[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_21 (.CI(n51532), .I0(n3155), .I1(n2977), .CO(n51533));
    SB_CARRY add_2797_8 (.CI(n51478), .I0(n2952), .I1(n1459), .CO(n51479));
    SB_LUT4 add_2793_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n51406), 
            .O(n8263[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n63621), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n11608));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n11608), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_2797_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n51477), 
            .O(n8367[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_6 (.CI(n51406), .I0(n2488), .I1(n1011), .CO(n51407));
    SB_LUT4 add_2793_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n51405), 
            .O(n8263[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_7 (.CI(n51477), .I0(n2953), .I1(n1460), .CO(n51478));
    SB_LUT4 add_2784_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n51307), 
            .O(n8029[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_5 (.CI(n51405), .I0(n2489), .I1(n856), .CO(n51406));
    SB_LUT4 add_2784_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n51306), 
            .O(n8029[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_8 (.CI(n51306), .I0(n1262), .I1(n1459), .CO(n51307));
    SB_LUT4 add_2793_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n51404), 
            .O(n8263[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n51531), 
            .O(n8419[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n51476), 
            .O(n8367[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2784_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n51305), 
            .O(n8029[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_4 (.CI(n51404), .I0(n2490), .I1(n698), .CO(n51405));
    SB_CARRY add_2797_6 (.CI(n51476), .I0(n2954), .I1(n1011), .CO(n51477));
    SB_LUT4 add_2793_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n51403), 
            .O(n8263[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_3 (.CI(n51403), .I0(n2491), .I1(n858), .CO(n51404));
    SB_CARRY add_2784_7 (.CI(n51305), .I0(n1263), .I1(n1460), .CO(n51306));
    SB_CARRY add_2799_20 (.CI(n51531), .I0(n3156), .I1(n2867), .CO(n51532));
    SB_LUT4 add_2797_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n51475), 
            .O(n8367[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_2_lut (.I0(n59082), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61354)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2797_5 (.CI(n51475), .I0(n2955), .I1(n856), .CO(n51476));
    SB_LUT4 add_2799_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n51530), 
            .O(n8419[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_19 (.CI(n51530), .I0(n3157), .I1(n2754), .CO(n51531));
    SB_CARRY add_2793_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51403));
    SB_LUT4 add_2797_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n51474), 
            .O(n8367[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n51529), 
            .O(n8419[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n51402), 
            .O(n8237[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_18 (.CI(n51529), .I0(n3158), .I1(n2638), .CO(n51530));
    SB_LUT4 add_2792_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n51401), 
            .O(n8237[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n51528), 
            .O(n8419[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_4 (.CI(n51474), .I0(n2956), .I1(n698), .CO(n51475));
    SB_LUT4 add_2797_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n51473), 
            .O(n8367[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2784_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n51304), 
            .O(n8029[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_6 (.CI(n51304), .I0(n1264), .I1(n1011), .CO(n51305));
    SB_LUT4 add_2784_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n51303), 
            .O(n8029[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_5 (.CI(n51303), .I0(n1265), .I1(n856), .CO(n51304));
    SB_CARRY add_2797_3 (.CI(n51473), .I0(n2957), .I1(n858), .CO(n51474));
    SB_CARRY add_2792_16 (.CI(n51401), .I0(n2354), .I1(n2519), .CO(n51402));
    SB_LUT4 add_2792_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n51400), 
            .O(n8237[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2784_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n51302), 
            .O(n8029[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_4 (.CI(n51302), .I0(n1266), .I1(n698), .CO(n51303));
    SB_CARRY add_2792_15 (.CI(n51400), .I0(n2355), .I1(n2397), .CO(n51401));
    SB_CARRY add_2799_17 (.CI(n51528), .I0(n3159), .I1(n2519), .CO(n51529));
    SB_LUT4 add_2797_2_lut (.I0(n59066), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61362)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2797_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51473));
    SB_LUT4 add_2799_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n51527), 
            .O(n8419[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2784_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n51301), 
            .O(n8029[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_3 (.CI(n51301), .I0(n1267), .I1(n858), .CO(n51302));
    SB_LUT4 add_2792_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n51399), 
            .O(n8237[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2796_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n51472), 
            .O(n8341[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_16 (.CI(n51527), .I0(n3160), .I1(n2397), .CO(n51528));
    SB_LUT4 add_2796_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n51471), 
            .O(n8341[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_20 (.CI(n51471), .I0(n2828), .I1(n2977), .CO(n51472));
    SB_LUT4 add_2796_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n51470), 
            .O(n8341[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n51526), 
            .O(n8419[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8393[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51521_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4939), .I3(\o_Rx_DV_N_3488[8] ), .O(n66373));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51521_4_lut.LUT_INIT = 16'hfffd;
    SB_CARRY add_2799_15 (.CI(n51526), .I0(n3161), .I1(n2272), .CO(n51527));
    SB_LUT4 i51597_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n57703), 
            .I3(r_SM_Main[0]), .O(n66379));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51597_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 add_2784_2_lut (.I0(n59112), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61344)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2784_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2799_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n51525), 
            .O(n8419[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2784_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51301));
    SB_CARRY add_2796_19 (.CI(n51470), .I0(n2829), .I1(n2867), .CO(n51471));
    SB_LUT4 add_2783_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n51300), 
            .O(n8003[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2783_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n51299), 
            .O(n8003[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51518_4_lut (.I0(n66373), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n66370));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51518_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51524_4_lut (.I0(n66379), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n66376));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51524_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY add_2799_14 (.CI(n51525), .I0(n3162), .I1(n2144), .CO(n51526));
    SB_LUT4 add_2796_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n51469), 
            .O(n8341[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n66376), .I1(n66370), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_4994));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 add_2799_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n51524), 
            .O(n8419[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_13 (.CI(n51524), .I0(n3163), .I1(n2013), .CO(n51525));
    SB_CARRY add_2796_18 (.CI(n51469), .I0(n2830), .I1(n2754), .CO(n51470));
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8393[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2796_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n51468), 
            .O(n8341[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_14 (.CI(n51399), .I0(n2356), .I1(n2272), .CO(n51400));
    SB_CARRY add_2783_7 (.CI(n51299), .I0(n1112), .I1(n1460), .CO(n51300));
    SB_LUT4 add_2783_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n51298), 
            .O(n8003[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n51523), 
            .O(n8419[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n51398), 
            .O(n8237[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_12 (.CI(n51523), .I0(n3164), .I1(n1879), .CO(n51524));
    SB_CARRY add_2796_17 (.CI(n51468), .I0(n2831), .I1(n2638), .CO(n51469));
    SB_CARRY add_2792_13 (.CI(n51398), .I0(n2357), .I1(n2144), .CO(n51399));
    SB_CARRY add_2783_6 (.CI(n51298), .I0(n1113), .I1(n1011), .CO(n51299));
    SB_LUT4 add_2792_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n51397), 
            .O(n8237[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8393[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2792_12 (.CI(n51397), .I0(n2358), .I1(n2013), .CO(n51398));
    SB_LUT4 add_2792_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n51396), 
            .O(n8237[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_11 (.CI(n51396), .I0(n2359), .I1(n1879), .CO(n51397));
    SB_LUT4 add_2799_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n51522), 
            .O(n8419[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2796_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n51467), 
            .O(n8341[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n51395), 
            .O(n8237[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2783_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n51297), 
            .O(n8003[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_5 (.CI(n51297), .I0(n1114), .I1(n856), .CO(n51298));
    SB_CARRY add_2796_16 (.CI(n51467), .I0(n2832), .I1(n2519), .CO(n51468));
    SB_CARRY add_2792_10 (.CI(n51395), .I0(n2360), .I1(n1742), .CO(n51396));
    SB_LUT4 add_2783_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n51296), 
            .O(n8003[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_4 (.CI(n51296), .I0(n1115), .I1(n698), .CO(n51297));
    SB_LUT4 add_2792_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n51394), 
            .O(n8237[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2796_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n51466), 
            .O(n8341[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_15 (.CI(n51466), .I0(n2833), .I1(n2397), .CO(n51467));
    SB_LUT4 add_2796_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n51465), 
            .O(n8341[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_11 (.CI(n51522), .I0(n3165), .I1(n1742), .CO(n51523));
    SB_CARRY add_2796_14 (.CI(n51465), .I0(n2834), .I1(n2272), .CO(n51466));
    SB_CARRY add_2792_9 (.CI(n51394), .I0(n2361), .I1(n1602), .CO(n51395));
    SB_LUT4 add_2792_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n51393), 
            .O(n8237[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2783_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n51295), 
            .O(n8003[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n51521), 
            .O(n8419[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2783_3 (.CI(n51295), .I0(n1116), .I1(n858), .CO(n51296));
    SB_CARRY add_2799_10 (.CI(n51521), .I0(n3166), .I1(n1602), .CO(n51522));
    SB_LUT4 add_2799_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n51520), 
            .O(n8419[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_9 (.CI(n51520), .I0(n3167), .I1(n1459), .CO(n51521));
    SB_LUT4 add_2783_2_lut (.I0(n59116), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61342)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2783_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2799_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n51519), 
            .O(n8419[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_8 (.CI(n51519), .I0(n3168), .I1(n1460), .CO(n51520));
    SB_LUT4 add_2799_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n51518), 
            .O(n8419[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8393[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8393[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2783_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51295));
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8393[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2796_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n51464), 
            .O(n8341[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47885_1_lut (.I0(n63601), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59066));
    defparam i47885_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2796_13 (.CI(n51464), .I0(n2835), .I1(n2144), .CO(n51465));
    SB_LUT4 add_2796_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n51463), 
            .O(n8341[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_12 (.CI(n51463), .I0(n2836), .I1(n2013), .CO(n51464));
    SB_CARRY add_2799_7 (.CI(n51518), .I0(n3169), .I1(n1011), .CO(n51519));
    SB_LUT4 add_2799_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n51517), 
            .O(n8419[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_8 (.CI(n51393), .I0(n2362), .I1(n1459), .CO(n51394));
    SB_CARRY add_2799_6 (.CI(n51517), .I0(n3170), .I1(n856), .CO(n51518));
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8393[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8393[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8393[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2796_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n51462), 
            .O(n8341[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n51516), 
            .O(n8419[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_11 (.CI(n51462), .I0(n2837), .I1(n1879), .CO(n51463));
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n50455), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n61330), .I1(n25566), .I2(VCC_net), 
            .I3(n50454), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_25 (.CI(n50454), .I0(n25566), .I1(VCC_net), 
            .CO(n50455));
    SB_CARRY add_2799_5 (.CI(n51516), .I0(n3171), .I1(n698), .CO(n51517));
    SB_LUT4 add_2796_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n51461), 
            .O(n8341[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n61418), .I1(n63639), .I2(VCC_net), 
            .I3(n50453), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8393[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2792_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n51392), 
            .O(n8237[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_24 (.CI(n50453), .I0(n63639), .I1(VCC_net), 
            .CO(n50454));
    SB_CARRY add_2796_10 (.CI(n51461), .I0(n2838), .I1(n1742), .CO(n51462));
    SB_CARRY add_2792_7 (.CI(n51392), .I0(n2363), .I1(n1460), .CO(n51393));
    SB_LUT4 add_2799_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n51515), 
            .O(n8419[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n51391), 
            .O(n8237[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2796_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n51460), 
            .O(n8341[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_6 (.CI(n51391), .I0(n2364), .I1(n1011), .CO(n51392));
    SB_CARRY add_2799_4 (.CI(n51515), .I0(n3172), .I1(n858), .CO(n51516));
    SB_LUT4 add_2792_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n51390), 
            .O(n8237[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_5 (.CI(n51390), .I0(n2365), .I1(n856), .CO(n51391));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n50452), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2796_9 (.CI(n51460), .I0(n2839), .I1(n1602), .CO(n51461));
    SB_LUT4 add_2796_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n51459), 
            .O(n8341[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_23 (.CI(n50452), .I0(n294[21]), .I1(VCC_net), 
            .CO(n50453));
    SB_LUT4 add_2792_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n51389), 
            .O(n8237[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_4 (.CI(n51389), .I0(n2366), .I1(n698), .CO(n51390));
    SB_LUT4 add_2792_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n51388), 
            .O(n8237[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_22_lut (.I0(n61416), .I1(n294[20]), .I2(VCC_net), 
            .I3(n50451), .O(n61418)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_22 (.CI(n50451), .I0(n294[20]), .I1(VCC_net), 
            .CO(n50452));
    SB_LUT4 sub_38_add_2_21_lut (.I0(n61414), .I1(n294[19]), .I2(VCC_net), 
            .I3(n50450), .O(n61416)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2799_3_lut (.I0(n59058), .I1(GND_net), .I2(n538), .I3(n51514), 
            .O(n61366)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2796_8 (.CI(n51459), .I0(n2840), .I1(n1459), .CO(n51460));
    SB_CARRY add_2792_3 (.CI(n51388), .I0(n2367), .I1(n858), .CO(n51389));
    SB_CARRY add_2799_3 (.CI(n51514), .I0(GND_net), .I1(n538), .CO(n51515));
    SB_LUT4 add_2792_2_lut (.I0(n59086), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61352)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2796_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n51458), 
            .O(n8341[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51388));
    SB_CARRY sub_38_add_2_21 (.CI(n50450), .I0(n294[19]), .I1(VCC_net), 
            .CO(n50451));
    SB_LUT4 add_2791_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n51387), 
            .O(n8211[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_7 (.CI(n51458), .I0(n2841), .I1(n1460), .CO(n51459));
    SB_CARRY add_2799_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n51514));
    SB_LUT4 add_2791_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n51386), 
            .O(n8211[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_15 (.CI(n51386), .I0(n2228), .I1(n2397), .CO(n51387));
    SB_LUT4 add_2796_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n51457), 
            .O(n8341[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n51385), 
            .O(n8211[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_6 (.CI(n51457), .I0(n2842), .I1(n1011), .CO(n51458));
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8393[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2791_14 (.CI(n51385), .I0(n2229), .I1(n2272), .CO(n51386));
    SB_LUT4 add_2791_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n51384), 
            .O(n8211[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8393[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8393[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n50449), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n51513), 
            .O(n8393[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n50449), .I0(n294[18]), .I1(VCC_net), 
            .CO(n50450));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n61412), .I1(n294[17]), .I2(VCC_net), 
            .I3(n50448), .O(n61414)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i47806_2_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n63523));
    defparam i47806_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2796_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n51456), 
            .O(n8341[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_13 (.CI(n51384), .I0(n2230), .I1(n2144), .CO(n51385));
    SB_CARRY sub_38_add_2_19 (.CI(n50448), .I0(n294[17]), .I1(VCC_net), 
            .CO(n50449));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n61410), .I1(n294[16]), .I2(VCC_net), 
            .I3(n50447), .O(n61412)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i7131_4_lut (.I0(n804), .I1(n42418), .I2(n20834), .I3(baudrate[2]), 
            .O(n20836));   // verilog/uart_rx.v(119[33:55])
    defparam i7131_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2798_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n51512), 
            .O(n8393[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_18 (.CI(n50447), .I0(n294[16]), .I1(VCC_net), 
            .CO(n50448));
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8393[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8367[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8367[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8367[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2796_5 (.CI(n51456), .I0(n2843), .I1(n856), .CO(n51457));
    SB_LUT4 add_2796_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n51455), 
            .O(n8341[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n51383), 
            .O(n8211[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8367[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8367[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8367[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n61328), .I1(n294[15]), .I2(VCC_net), 
            .I3(n50446), .O(n61330)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2791_12 (.CI(n51383), .I0(n2231), .I1(n2013), .CO(n51384));
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8367[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2796_4 (.CI(n51455), .I0(n2844), .I1(n698), .CO(n51456));
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8367[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8367[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2791_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n51382), 
            .O(n8211[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4995));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8367[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4996));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_17 (.CI(n50446), .I0(n294[15]), .I1(VCC_net), 
            .CO(n50447));
    SB_LUT4 sub_38_add_2_16_lut (.I0(n61408), .I1(n294[14]), .I2(VCC_net), 
            .I3(n50445), .O(n61410)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2791_11 (.CI(n51382), .I0(n2232), .I1(n1879), .CO(n51383));
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4997));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8367[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8367[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4998));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4999));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8367[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2798_22 (.CI(n51512), .I0(n3047), .I1(n3188), .CO(n51513));
    SB_LUT4 add_2796_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n51454), 
            .O(n8341[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8367[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2798_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n51511), 
            .O(n8393[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_3 (.CI(n51454), .I0(n2845), .I1(n858), .CO(n51455));
    SB_LUT4 add_2791_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n51381), 
            .O(n8211[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_10 (.CI(n51381), .I0(n2233), .I1(n1742), .CO(n51382));
    SB_LUT4 add_2791_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n51380), 
            .O(n8211[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_16 (.CI(n50445), .I0(n294[14]), .I1(VCC_net), 
            .CO(n50446));
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8367[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8367[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5000));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8367[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2796_2_lut (.I0(n59070), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61360)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n50444), .O(n61408)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5001));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8315[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8341[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8341[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5002));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2791_9 (.CI(n51380), .I0(n2234), .I1(n1602), .CO(n51381));
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5003));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5004));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5005));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5006));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5007));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2791_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n51379), 
            .O(n8211[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n50444), .I0(n294[13]), .I1(VCC_net), 
            .CO(n50445));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n50443), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5008));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5009));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2796_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51454));
    SB_CARRY add_2791_8 (.CI(n51379), .I0(n2235), .I1(n1459), .CO(n51380));
    SB_CARRY sub_38_add_2_14 (.CI(n50443), .I0(n294[12]), .I1(VCC_net), 
            .CO(n50444));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n50442), .O(n61328)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2798_21 (.CI(n51511), .I0(n3048), .I1(n3084), .CO(n51512));
    SB_LUT4 add_2795_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n51453), 
            .O(n8315[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n51510), 
            .O(n8393[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n51378), 
            .O(n8211[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_13 (.CI(n50442), .I0(n294[11]), .I1(VCC_net), 
            .CO(n50443));
    SB_LUT4 add_2795_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n51452), 
            .O(n8315[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2791_7 (.CI(n51378), .I0(n2236), .I1(n1460), .CO(n51379));
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2791_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n51377), 
            .O(n8211[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5010));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2791_6 (.CI(n51377), .I0(n2237), .I1(n1011), .CO(n51378));
    SB_LUT4 i5760_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n59555), .I3(n44_adj_5011), 
            .O(n46_adj_5012));   // verilog/uart_rx.v(119[33:55])
    defparam i5760_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5014));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n50441), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(n69211), .I1(baudrate[11]), .I2(n1831), 
            .I3(n61348), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8419[20]), .I3(n294[1]), .O(n41_adj_5015));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8419[19]), .I3(n294[1]), .O(n39_adj_5016));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_12 (.CI(n50441), .I0(n294[10]), .I1(VCC_net), 
            .CO(n50442));
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8419[17]), .I3(n294[1]), .O(n35_adj_5017));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5018));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5019));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8419[18]), .I3(n294[1]), .O(n37_adj_5020));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8419[14]), .I3(n294[1]), .O(n29_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8289[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2795_19 (.CI(n51452), .I0(n2714), .I1(n2867), .CO(n51453));
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8419[15]), .I3(n294[1]), .O(n31_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8419[11]), .I3(n294[1]), .O(n23_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i742_4_lut (.I0(n58836), .I1(n294[18]), .I2(n46_adj_5012), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54345_2_lut_4_lut (.I0(n69211), .I1(baudrate[11]), .I2(n1831), 
            .I3(n63577), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i54345_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8419[12]), .I3(n294[1]), .O(n25_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2791_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n51376), 
            .O(n8211[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51429_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n67155));   // verilog/uart_rx.v(119[33:55])
    defparam i51429_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8419[16]), .I3(n294[1]), .O(n33_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8419[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8419[22]), .I3(n294[1]), .O(n45_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8419[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8419[8]), .I3(n294[1]), .O(n17_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8419[9]), .I3(n294[1]), .O(n19_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51176_4_lut (.I0(n37_adj_5033), .I1(n25_adj_5028), .I2(n23_adj_5025), 
            .I3(n21_adj_5024), .O(n66902));
    defparam i51176_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2791_5 (.CI(n51376), .I0(n2238), .I1(n856), .CO(n51377));
    SB_LUT4 i52080_4_lut (.I0(n19_adj_5023), .I1(n17_adj_5022), .I2(n2729), 
            .I3(baudrate[2]), .O(n67806));
    defparam i52080_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52645_4_lut (.I0(n25_adj_5028), .I1(n23_adj_5025), .I2(n21_adj_5024), 
            .I3(n67806), .O(n68371));
    defparam i52645_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52641_4_lut (.I0(n31_adj_5042), .I1(n29_adj_5039), .I2(n27_adj_5034), 
            .I3(n68371), .O(n68367));
    defparam i52641_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51178_4_lut (.I0(n37_adj_5033), .I1(n35_adj_5030), .I2(n33_adj_5029), 
            .I3(n68367), .O(n66904));
    defparam i51178_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53091_3_lut (.I0(n14), .I1(baudrate[13]), .I2(n37_adj_5033), 
            .I3(GND_net), .O(n68817));   // verilog/uart_rx.v(119[33:55])
    defparam i53091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8003[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8029[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8055[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53092_3_lut (.I0(n68817), .I1(baudrate[14]), .I2(n39_adj_5019), 
            .I3(GND_net), .O(n68818));   // verilog/uart_rx.v(119[33:55])
    defparam i53092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8081[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8107[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8133[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8159[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8185[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8211[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8237[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8263[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8289[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8315[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_978 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n62822));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_adj_979 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n62724));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_980 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n62726));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'heeee;
    SB_CARRY add_2798_20 (.CI(n51510), .I0(n3049), .I1(n2977), .CO(n51511));
    SB_LUT4 add_2795_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n51451), 
            .O(n8315[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8419[10]), .I3(n294[1]), .O(n21_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2791_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n51375), 
            .O(n8211[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n51509), 
            .O(n8393[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8419[21]), .I3(n294[1]), .O(n43_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8419[5]), .I3(n294[1]), .O(n11_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22), .I1(baudrate[17]), 
            .I2(n45), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51171_4_lut (.I0(n43), .I1(n41_adj_5018), .I2(n39_adj_5019), 
            .I3(n66902), .O(n66897));
    defparam i51171_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52665_4_lut (.I0(n40), .I1(n20), .I2(n45), .I3(n66895), 
            .O(n68391));   // verilog/uart_rx.v(119[33:55])
    defparam i52665_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8419[6]), .I3(n294[1]), .O(n13_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8419[7]), .I3(n294[1]), .O(n15_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i52988_3_lut (.I0(n68818), .I1(baudrate[15]), .I2(n41_adj_5018), 
            .I3(GND_net), .O(n68714));   // verilog/uart_rx.v(119[33:55])
    defparam i52988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8419[13]), .I3(n294[1]), .O(n27_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i50896_4_lut (.I0(n27_adj_5048), .I1(n15_adj_5047), .I2(n13_adj_5046), 
            .I3(n11_adj_5045), .O(n66622));
    defparam i50896_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50914_4_lut (.I0(n21_adj_5043), .I1(n19_adj_5041), .I2(n17_adj_5040), 
            .I3(n9), .O(n66640));
    defparam i50914_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5044), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50834_2_lut (.I0(n43_adj_5044), .I1(n19_adj_5041), .I2(GND_net), 
            .I3(GND_net), .O(n66560));
    defparam i50834_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18), .I1(baudrate[9]), 
            .I2(n29_adj_5039), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53401_4_lut (.I0(n26), .I1(n16_adj_5049), .I2(n29_adj_5039), 
            .I3(n66918), .O(n69127));   // verilog/uart_rx.v(119[33:55])
    defparam i53401_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53402_3_lut (.I0(n69127), .I1(baudrate[10]), .I2(n31_adj_5042), 
            .I3(GND_net), .O(n69128));   // verilog/uart_rx.v(119[33:55])
    defparam i53402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5040), .I3(GND_net), .O(n8_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53295_3_lut (.I0(n69128), .I1(baudrate[11]), .I2(n33_adj_5029), 
            .I3(GND_net), .O(n69021));   // verilog/uart_rx.v(119[33:55])
    defparam i53295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52939_4_lut (.I0(n43), .I1(n41_adj_5018), .I2(n39_adj_5019), 
            .I3(n66904), .O(n68665));
    defparam i52939_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53239_4_lut (.I0(n68714), .I1(n68391), .I2(n45), .I3(n66897), 
            .O(n68965));   // verilog/uart_rx.v(119[33:55])
    defparam i53239_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53238_3_lut (.I0(n69021), .I1(baudrate[12]), .I2(n35_adj_5030), 
            .I3(GND_net), .O(n68964));   // verilog/uart_rx.v(119[33:55])
    defparam i53238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53241_4_lut (.I0(n68964), .I1(n68965), .I2(n45), .I3(n68665), 
            .O(n68967));   // verilog/uart_rx.v(119[33:55])
    defparam i53241_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8289[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8315[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16), .I1(baudrate[22]), 
            .I2(n45_adj_5038), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8419[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8341[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29596));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29595));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29591));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29590));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29559));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29558));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29557));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n70507));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2795_18 (.CI(n51451), .I0(n2715), .I1(n2754), .CO(n51452));
    SB_CARRY add_2798_19 (.CI(n51509), .I0(n3050), .I1(n2867), .CO(n51510));
    SB_CARRY add_2791_4 (.CI(n51375), .I0(n2239), .I1(n698), .CO(n51376));
    SB_LUT4 add_2791_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n51374), 
            .O(n8211[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50930_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n66656));
    defparam i50930_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i51814_4_lut (.I0(n13_adj_5046), .I1(n11_adj_5045), .I2(n9), 
            .I3(n66656), .O(n67540));
    defparam i51814_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51808_4_lut (.I0(n19_adj_5041), .I1(n17_adj_5040), .I2(n15_adj_5047), 
            .I3(n67540), .O(n67534));
    defparam i51808_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53135_4_lut (.I0(n25_adj_5035), .I1(n23_adj_5032), .I2(n21_adj_5043), 
            .I3(n67534), .O(n68861));
    defparam i53135_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2798_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n51508), 
            .O(n8393[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n50440), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_3 (.CI(n51374), .I0(n2240), .I1(n858), .CO(n51375));
    SB_LUT4 i52521_4_lut (.I0(n31_adj_5027), .I1(n29_adj_5021), .I2(n27_adj_5048), 
            .I3(n68861), .O(n68247));
    defparam i52521_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53350_4_lut (.I0(n37_adj_5020), .I1(n35_adj_5017), .I2(n33_adj_5037), 
            .I3(n68247), .O(n69076));
    defparam i53350_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2791_2_lut (.I0(n59090), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61350)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5037), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61366), .I3(n48), .O(n4));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53061_3_lut (.I0(n4), .I1(baudrate[13]), .I2(n27_adj_5048), 
            .I3(GND_net), .O(n68787));   // verilog/uart_rx.v(119[33:55])
    defparam i53061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51264_4_lut (.I0(n23_adj_5062), .I1(n21_adj_5061), .I2(n19_adj_5060), 
            .I3(n17_adj_5064), .O(n66990));
    defparam i51264_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51257_4_lut (.I0(n29_adj_5059), .I1(n27_adj_5058), .I2(n25_adj_5063), 
            .I3(n66990), .O(n66983));
    defparam i51257_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52971_4_lut (.I0(n35_adj_5057), .I1(n33_adj_5056), .I2(n31_adj_5055), 
            .I3(n66983), .O(n68697));
    defparam i52971_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53097_3_lut (.I0(n16_adj_5065), .I1(baudrate[13]), .I2(n39_adj_5054), 
            .I3(GND_net), .O(n68823));   // verilog/uart_rx.v(119[33:55])
    defparam i53097_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_11 (.CI(n50440), .I0(n294[9]), .I1(VCC_net), 
            .CO(n50441));
    SB_LUT4 add_2795_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n51450), 
            .O(n8315[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53062_3_lut (.I0(n68787), .I1(baudrate[14]), .I2(n29_adj_5021), 
            .I3(GND_net), .O(n68788));   // verilog/uart_rx.v(119[33:55])
    defparam i53062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50876_2_lut (.I0(n33_adj_5037), .I1(n15_adj_5047), .I2(GND_net), 
            .I3(GND_net), .O(n66602));
    defparam i50876_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_5046), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2795_17 (.CI(n51450), .I0(n2716), .I1(n2638), .CO(n51451));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n50439), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n51449), 
            .O(n8315[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51374));
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12), .I1(baudrate[17]), 
            .I2(n35_adj_5017), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50882_4_lut (.I0(n33_adj_5037), .I1(n31_adj_5027), .I2(n29_adj_5021), 
            .I3(n66622), .O(n66608));
    defparam i50882_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53413_4_lut (.I0(n30), .I1(n10), .I2(n35_adj_5017), .I3(n66602), 
            .O(n69139));   // verilog/uart_rx.v(119[33:55])
    defparam i53413_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53098_3_lut (.I0(n68823), .I1(baudrate[14]), .I2(n41_adj_5053), 
            .I3(GND_net), .O(n68824));   // verilog/uart_rx.v(119[33:55])
    defparam i53098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52097_4_lut (.I0(n41_adj_5053), .I1(n39_adj_5054), .I2(n27_adj_5058), 
            .I3(n66986), .O(n67823));
    defparam i52097_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52663_3_lut (.I0(n22_adj_5066), .I1(baudrate[7]), .I2(n27_adj_5058), 
            .I3(GND_net), .O(n68389));   // verilog/uart_rx.v(119[33:55])
    defparam i52663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52981_3_lut (.I0(n68824), .I1(baudrate[15]), .I2(n43_adj_5052), 
            .I3(GND_net), .O(n68707));   // verilog/uart_rx.v(119[33:55])
    defparam i52981_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2798_18 (.CI(n51508), .I0(n3051), .I1(n2754), .CO(n51509));
    SB_LUT4 add_2798_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n51507), 
            .O(n8393[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5067), .I1(baudrate[9]), 
            .I2(n31_adj_5055), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53399_4_lut (.I0(n28), .I1(n18_adj_5068), .I2(n31_adj_5055), 
            .I3(n66967), .O(n69125));   // verilog/uart_rx.v(119[33:55])
    defparam i53399_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53020_3_lut (.I0(n68788), .I1(baudrate[15]), .I2(n31_adj_5027), 
            .I3(GND_net), .O(n68746));   // verilog/uart_rx.v(119[33:55])
    defparam i53020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53530_4_lut (.I0(n68746), .I1(n69139), .I2(n35_adj_5017), 
            .I3(n66608), .O(n69256));   // verilog/uart_rx.v(119[33:55])
    defparam i53530_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53400_3_lut (.I0(n69125), .I1(baudrate[10]), .I2(n33_adj_5056), 
            .I3(GND_net), .O(n69126));   // verilog/uart_rx.v(119[33:55])
    defparam i53400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53297_3_lut (.I0(n69126), .I1(baudrate[11]), .I2(n35_adj_5057), 
            .I3(GND_net), .O(n69023));   // verilog/uart_rx.v(119[33:55])
    defparam i53297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52108_4_lut (.I0(n41_adj_5053), .I1(n39_adj_5054), .I2(n37_adj_5051), 
            .I3(n68697), .O(n67834));
    defparam i52108_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53095_4_lut (.I0(n68707), .I1(n68389), .I2(n43_adj_5052), 
            .I3(n67823), .O(n68821));   // verilog/uart_rx.v(119[33:55])
    defparam i53095_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53236_3_lut (.I0(n69023), .I1(baudrate[12]), .I2(n37_adj_5051), 
            .I3(GND_net), .O(n68962));   // verilog/uart_rx.v(119[33:55])
    defparam i53236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53419_4_lut (.I0(n68962), .I1(n68821), .I2(n43_adj_5052), 
            .I3(n67834), .O(n69145));   // verilog/uart_rx.v(119[33:55])
    defparam i53419_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53531_3_lut (.I0(n69256), .I1(baudrate[18]), .I2(n37_adj_5020), 
            .I3(GND_net), .O(n69257));   // verilog/uart_rx.v(119[33:55])
    defparam i53531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_1952__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27766), .D(n1[0]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27766), .D(n1[1]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27766), .D(n1[2]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27766), .D(n1[3]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27766), .D(n1[4]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27766), .D(n1[5]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27766), .D(n1[6]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1952__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27766), .D(n1[7]), .R(n29073));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i53063_3_lut (.I0(n6), .I1(baudrate[10]), .I2(n21_adj_5043), 
            .I3(GND_net), .O(n68789));   // verilog/uart_rx.v(119[33:55])
    defparam i53063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53064_3_lut (.I0(n68789), .I1(baudrate[11]), .I2(n23_adj_5032), 
            .I3(GND_net), .O(n68790));   // verilog/uart_rx.v(119[33:55])
    defparam i53064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53420_3_lut (.I0(n69145), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n69146));   // verilog/uart_rx.v(119[33:55])
    defparam i53420_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_38_add_2_10 (.CI(n50439), .I0(n294[8]), .I1(VCC_net), 
            .CO(n50440));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n50438), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n51373), 
            .O(n8185[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n50438), .I0(n294[7]), .I1(VCC_net), 
            .CO(n50439));
    SB_LUT4 add_2790_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n51372), 
            .O(n8185[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50838_4_lut (.I0(n43_adj_5044), .I1(n25_adj_5035), .I2(n23_adj_5032), 
            .I3(n66640), .O(n66564));
    defparam i50838_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8315[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8341[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8341[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n50437), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_13 (.CI(n51372), .I0(n2099), .I1(n2272), .CO(n51373));
    SB_LUT4 i52675_4_lut (.I0(n24), .I1(n8_adj_5050), .I2(n45_adj_5038), 
            .I3(n66560), .O(n68401));   // verilog/uart_rx.v(119[33:55])
    defparam i52675_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_38_add_2_8 (.CI(n50437), .I0(n294[6]), .I1(VCC_net), 
            .CO(n50438));
    SB_LUT4 i53018_3_lut (.I0(n68790), .I1(baudrate[12]), .I2(n25_adj_5035), 
            .I3(GND_net), .O(n68744));   // verilog/uart_rx.v(119[33:55])
    defparam i53018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n50436), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8289[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8315[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8341[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53475_3_lut (.I0(n69257), .I1(baudrate[19]), .I2(n39_adj_5016), 
            .I3(GND_net), .O(n69201));   // verilog/uart_rx.v(119[33:55])
    defparam i53475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50843_4_lut (.I0(n43_adj_5044), .I1(n41_adj_5015), .I2(n39_adj_5016), 
            .I3(n69076), .O(n66569));
    defparam i50843_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53256_4_lut (.I0(n68744), .I1(n68401), .I2(n45_adj_5038), 
            .I3(n66564), .O(n68982));   // verilog/uart_rx.v(119[33:55])
    defparam i53256_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2798_17 (.CI(n51507), .I0(n3052), .I1(n2638), .CO(n51508));
    SB_LUT4 i53471_3_lut (.I0(n69201), .I1(baudrate[20]), .I2(n41_adj_5015), 
            .I3(GND_net), .O(n40_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam i53471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_981 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n61294));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8419[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47828_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n63545));
    defparam i47828_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i47884_4_lut (.I0(n63545), .I1(n62814), .I2(n63543), .I3(n62768), 
            .O(n63601));
    defparam i47884_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2795_16 (.CI(n51449), .I0(n2717), .I1(n2519), .CO(n51450));
    SB_LUT4 i51082_4_lut (.I0(n33_adj_5081), .I1(n21_adj_5080), .I2(n19_adj_5079), 
            .I3(n17_adj_5077), .O(n66808));
    defparam i51082_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47782_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n63499));
    defparam i47782_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47900_4_lut (.I0(n63499), .I1(n61988), .I2(n62726), .I3(baudrate[9]), 
            .O(n63617));
    defparam i47900_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51998_4_lut (.I0(n15_adj_5076), .I1(n13_adj_5075), .I2(n2956), 
            .I3(baudrate[2]), .O(n67724));
    defparam i51998_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53258_4_lut (.I0(n40_adj_5078), .I1(n68982), .I2(n45_adj_5038), 
            .I3(n66569), .O(n68984));   // verilog/uart_rx.v(119[33:55])
    defparam i53258_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_982 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n61664));
    defparam i1_4_lut_adj_982.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_983 (.I0(n62914), .I1(n62772), .I2(n61294), .I3(n62770), 
            .O(n61302));
    defparam i1_4_lut_adj_983.LUT_INIT = 16'hfffe;
    SB_LUT4 i54046_4_lut (.I0(n61302), .I1(n68984), .I2(baudrate[23]), 
            .I3(n3253), .O(n60390));   // verilog/uart_rx.v(119[33:55])
    defparam i54046_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52605_4_lut (.I0(n21_adj_5080), .I1(n19_adj_5079), .I2(n17_adj_5077), 
            .I3(n67724), .O(n68331));
    defparam i52605_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52603_4_lut (.I0(n27_adj_5007), .I1(n25_adj_5006), .I2(n23_adj_5005), 
            .I3(n68331), .O(n68329));
    defparam i52603_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i47846_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n63563));
    defparam i47846_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51087_4_lut (.I0(n33_adj_5081), .I1(n31), .I2(n29_adj_5008), 
            .I3(n68329), .O(n66813));
    defparam i51087_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_984 (.I0(n58877), .I1(n61664), .I2(n62914), .I3(baudrate[16]), 
            .O(n61692));
    defparam i1_4_lut_adj_984.LUT_INIT = 16'h0004;
    SB_LUT4 i47912_4_lut (.I0(n63563), .I1(n63475), .I2(n63483), .I3(n63298), 
            .O(n63629));
    defparam i47912_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53578_4_lut (.I0(n63617), .I1(n66729), .I2(n63629), .I3(n61692), 
            .O(n69304));
    defparam i53578_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i2161_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2161_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53081_3_lut (.I0(n10_adj_5084), .I1(baudrate[13]), .I2(n33_adj_5081), 
            .I3(GND_net), .O(n68807));   // verilog/uart_rx.v(119[33:55])
    defparam i53081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53082_3_lut (.I0(n68807), .I1(baudrate[14]), .I2(n35_adj_5003), 
            .I3(GND_net), .O(n68808));   // verilog/uart_rx.v(119[33:55])
    defparam i53082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i535_4_lut (.I0(n69304), .I1(n44_adj_5086), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 add_2790_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n51371), 
            .O(n8185[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5090), .I1(baudrate[17]), 
            .I2(n41), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5011), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i51076_4_lut (.I0(n39_adj_5004), .I1(n37_adj_5002), .I2(n35_adj_5003), 
            .I3(n66808), .O(n66802));
    defparam i51076_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53407_4_lut (.I0(n36), .I1(n16_adj_5092), .I2(n41), .I3(n66800), 
            .O(n69133));   // verilog/uart_rx.v(119[33:55])
    defparam i53407_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52998_3_lut (.I0(n68808), .I1(baudrate[15]), .I2(n37_adj_5002), 
            .I3(GND_net), .O(n68724));   // verilog/uart_rx.v(119[33:55])
    defparam i52998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5093), .I1(baudrate[9]), 
            .I2(n25_adj_5006), .I3(GND_net), .O(n22_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5095));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53405_4_lut (.I0(n22_adj_5094), .I1(n12_adj_5096), .I2(n25_adj_5006), 
            .I3(n66822), .O(n69131));   // verilog/uart_rx.v(119[33:55])
    defparam i53405_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2790_12 (.CI(n51371), .I0(n2100), .I1(n2144), .CO(n51372));
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n61043));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8003[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53406_3_lut (.I0(n69131), .I1(baudrate[10]), .I2(n27_adj_5007), 
            .I3(GND_net), .O(n69132));   // verilog/uart_rx.v(119[33:55])
    defparam i53406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8029[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53289_3_lut (.I0(n69132), .I1(baudrate[11]), .I2(n29_adj_5008), 
            .I3(GND_net), .O(n69015));   // verilog/uart_rx.v(119[33:55])
    defparam i53289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8055[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8081[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2795_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n51448), 
            .O(n8315[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_15 (.CI(n51448), .I0(n2718), .I1(n2397), .CO(n51449));
    SB_LUT4 i2154_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2154_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52899_4_lut (.I0(n39_adj_5004), .I1(n37_adj_5002), .I2(n35_adj_5003), 
            .I3(n66813), .O(n68625));
    defparam i52899_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53524_4_lut (.I0(n68724), .I1(n69133), .I2(n41), .I3(n66802), 
            .O(n69250));   // verilog/uart_rx.v(119[33:55])
    defparam i53524_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53247_3_lut (.I0(n69015), .I1(baudrate[12]), .I2(n31), .I3(GND_net), 
            .O(n68973));   // verilog/uart_rx.v(119[33:55])
    defparam i53247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53546_4_lut (.I0(n68973), .I1(n69250), .I2(n41), .I3(n68625), 
            .O(n69272));   // verilog/uart_rx.v(119[33:55])
    defparam i53546_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53547_3_lut (.I0(n69272), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n69273));   // verilog/uart_rx.v(119[33:55])
    defparam i53547_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53543_3_lut (.I0(n69273), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n69269));   // verilog/uart_rx.v(119[33:55])
    defparam i53543_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2790_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n51370), 
            .O(n8185[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8341[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8367[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53782_3_lut (.I0(n25593), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25566));   // verilog/uart_rx.v(119[33:55])
    defparam i53782_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50954_4_lut (.I0(n29_adj_5102), .I1(n17_adj_5101), .I2(n15_adj_5100), 
            .I3(n13_adj_5099), .O(n66680));
    defparam i50954_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8367[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_7 (.CI(n50436), .I0(n294[5]), .I1(VCC_net), 
            .CO(n50437));
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51012_4_lut (.I0(n31_adj_5108), .I1(n19_adj_5107), .I2(n17_adj_5106), 
            .I3(n15_adj_5105), .O(n66738));
    defparam i51012_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2790_11 (.CI(n51370), .I0(n2101), .I1(n2013), .CO(n51371));
    SB_LUT4 i51948_4_lut (.I0(n13), .I1(n11), .I2(n3065), .I3(baudrate[2]), 
            .O(n67674));
    defparam i51948_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51860_4_lut (.I0(n11_adj_5103), .I1(n9_adj_5098), .I2(n3171), 
            .I3(baudrate[2]), .O(n67586));
    defparam i51860_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52583_4_lut (.I0(n19_adj_5107), .I1(n17_adj_5106), .I2(n15_adj_5105), 
            .I3(n67674), .O(n68309));
    defparam i52583_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52555_4_lut (.I0(n17_adj_5101), .I1(n15_adj_5100), .I2(n13_adj_5099), 
            .I3(n67586), .O(n68281));
    defparam i52555_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52551_4_lut (.I0(n23_adj_5097), .I1(n21_adj_5091), .I2(n19_adj_5104), 
            .I3(n68281), .O(n68277));
    defparam i52551_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50956_4_lut (.I0(n29_adj_5102), .I1(n27_adj_5089), .I2(n25_adj_5088), 
            .I3(n68277), .O(n66682));
    defparam i50956_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2790_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n51369), 
            .O(n8185[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n51506), 
            .O(n8393[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n51447), 
            .O(n8315[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53069_3_lut (.I0(n6_adj_5109), .I1(baudrate[13]), .I2(n29_adj_5102), 
            .I3(GND_net), .O(n68795));   // verilog/uart_rx.v(119[33:55])
    defparam i53069_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30440));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n53943));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30436));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i52579_4_lut (.I0(n25), .I1(n23_adj_4999), .I2(n21_adj_5000), 
            .I3(n68309), .O(n68305));
    defparam i52579_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2790_10 (.CI(n51369), .I0(n2102), .I1(n1879), .CO(n51370));
    SB_LUT4 add_2790_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n51368), 
            .O(n8185[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51016_4_lut (.I0(n31_adj_5108), .I1(n29_adj_4997), .I2(n27_adj_4996), 
            .I3(n68305), .O(n66742));
    defparam i51016_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n50435), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n50435), .I0(n294[4]), .I1(VCC_net), 
            .CO(n50436));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n50434), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53075_3_lut (.I0(n8_adj_5110), .I1(baudrate[13]), .I2(n31_adj_5108), 
            .I3(GND_net), .O(n68801));   // verilog/uart_rx.v(119[33:55])
    defparam i53075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53076_3_lut (.I0(n68801), .I1(baudrate[14]), .I2(n33), .I3(GND_net), 
            .O(n68802));   // verilog/uart_rx.v(119[33:55])
    defparam i53076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5111), .I1(baudrate[17]), 
            .I2(n37_adj_5083), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53070_3_lut (.I0(n68795), .I1(baudrate[14]), .I2(n31_adj_5085), 
            .I3(GND_net), .O(n68796));   // verilog/uart_rx.v(119[33:55])
    defparam i53070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50949_4_lut (.I0(n35_adj_5087), .I1(n33_adj_5082), .I2(n31_adj_5085), 
            .I3(n66680), .O(n66675));
    defparam i50949_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5112), .I1(baudrate[17]), 
            .I2(n39), .I3(GND_net), .O(n34_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_5 (.CI(n50434), .I0(n294[3]), .I1(VCC_net), 
            .CO(n50435));
    SB_LUT4 i53411_4_lut (.I0(n32), .I1(n12_adj_5114), .I2(n37_adj_5083), 
            .I3(n66673), .O(n69137));   // verilog/uart_rx.v(119[33:55])
    defparam i53411_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51005_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n66738), 
            .O(n66731));
    defparam i51005_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53409_4_lut (.I0(n34_adj_5113), .I1(n14_adj_5115), .I2(n39), 
            .I3(n66722), .O(n69135));   // verilog/uart_rx.v(119[33:55])
    defparam i53409_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53004_3_lut (.I0(n68802), .I1(baudrate[15]), .I2(n35), .I3(GND_net), 
            .O(n68730));   // verilog/uart_rx.v(119[33:55])
    defparam i53004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53077_3_lut (.I0(n10_adj_5116), .I1(baudrate[10]), .I2(n25), 
            .I3(GND_net), .O(n68803));   // verilog/uart_rx.v(119[33:55])
    defparam i53077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53078_3_lut (.I0(n68803), .I1(baudrate[11]), .I2(n27_adj_4996), 
            .I3(GND_net), .O(n68804));   // verilog/uart_rx.v(119[33:55])
    defparam i53078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51928_4_lut (.I0(n27_adj_4996), .I1(n25), .I2(n23_adj_4999), 
            .I3(n66753), .O(n67654));
    defparam i51928_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2795_14 (.CI(n51447), .I0(n2719), .I1(n2272), .CO(n51448));
    SB_CARRY add_2790_9 (.CI(n51368), .I0(n2103), .I1(n1742), .CO(n51369));
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5117), .I1(baudrate[9]), 
            .I2(n23_adj_4999), .I3(GND_net), .O(n20_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53002_3_lut (.I0(n68804), .I1(baudrate[12]), .I2(n29_adj_4997), 
            .I3(GND_net), .O(n26_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam i53002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8107[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2790_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n51367), 
            .O(n8185[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53010_3_lut (.I0(n68796), .I1(baudrate[15]), .I2(n33_adj_5082), 
            .I3(GND_net), .O(n68736));   // verilog/uart_rx.v(119[33:55])
    defparam i53010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52885_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n66742), 
            .O(n68611));
    defparam i52885_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53526_4_lut (.I0(n68730), .I1(n69135), .I2(n39), .I3(n66731), 
            .O(n69252));   // verilog/uart_rx.v(119[33:55])
    defparam i53526_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53071_3_lut (.I0(n8_adj_5120), .I1(baudrate[10]), .I2(n23_adj_5097), 
            .I3(GND_net), .O(n68797));   // verilog/uart_rx.v(119[33:55])
    defparam i53071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53072_3_lut (.I0(n68797), .I1(baudrate[11]), .I2(n25_adj_5088), 
            .I3(GND_net), .O(n68798));   // verilog/uart_rx.v(119[33:55])
    defparam i53072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51840_4_lut (.I0(n25_adj_5088), .I1(n23_adj_5097), .I2(n21_adj_5091), 
            .I3(n66692), .O(n67566));
    defparam i51840_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52669_4_lut (.I0(n26_adj_5119), .I1(n20_adj_5118), .I2(n29_adj_4997), 
            .I3(n67654), .O(n68395));   // verilog/uart_rx.v(119[33:55])
    defparam i52669_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53550_4_lut (.I0(n68395), .I1(n69252), .I2(n39), .I3(n68611), 
            .O(n69276));   // verilog/uart_rx.v(119[33:55])
    defparam i53550_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52673_3_lut (.I0(n10_adj_5121), .I1(baudrate[9]), .I2(n21_adj_5091), 
            .I3(GND_net), .O(n68399));   // verilog/uart_rx.v(119[33:55])
    defparam i52673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53551_3_lut (.I0(n69276), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n69277));   // verilog/uart_rx.v(119[33:55])
    defparam i53551_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53539_3_lut (.I0(n69277), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n69265));   // verilog/uart_rx.v(119[33:55])
    defparam i53539_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53008_3_lut (.I0(n68798), .I1(baudrate[12]), .I2(n27_adj_5089), 
            .I3(GND_net), .O(n68734));   // verilog/uart_rx.v(119[33:55])
    defparam i53008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52858_4_lut (.I0(n35_adj_5087), .I1(n33_adj_5082), .I2(n31_adj_5085), 
            .I3(n66682), .O(n68584));
    defparam i52858_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52671_3_lut (.I0(n69265), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n68397));   // verilog/uart_rx.v(119[33:55])
    defparam i52671_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n50433), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_8 (.CI(n51367), .I0(n2104), .I1(n1602), .CO(n51368));
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8367[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2798_16 (.CI(n51506), .I0(n3053), .I1(n2519), .CO(n51507));
    SB_LUT4 add_2798_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n51505), 
            .O(n8393[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n51446), 
            .O(n8315[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_15 (.CI(n51505), .I0(n3054), .I1(n2397), .CO(n51506));
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2790_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n51366), 
            .O(n8185[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8393[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53528_4_lut (.I0(n68736), .I1(n69137), .I2(n37_adj_5083), 
            .I3(n66675), .O(n69254));   // verilog/uart_rx.v(119[33:55])
    defparam i53528_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2798_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n51504), 
            .O(n8393[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_13 (.CI(n51446), .I0(n2720), .I1(n2144), .CO(n51447));
    SB_LUT4 i53065_4_lut (.I0(n68734), .I1(n68399), .I2(n27_adj_5089), 
            .I3(n67566), .O(n68791));   // verilog/uart_rx.v(119[33:55])
    defparam i53065_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53548_4_lut (.I0(n68791), .I1(n69254), .I2(n37_adj_5083), 
            .I3(n68584), .O(n69274));   // verilog/uart_rx.v(119[33:55])
    defparam i53548_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53549_3_lut (.I0(n69274), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n69275));   // verilog/uart_rx.v(119[33:55])
    defparam i53549_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53541_3_lut (.I0(n69275), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n69267));   // verilog/uart_rx.v(119[33:55])
    defparam i53541_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2795_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n51445), 
            .O(n8315[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53344_3_lut (.I0(n69267), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n69070));   // verilog/uart_rx.v(119[33:55])
    defparam i53344_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53345_3_lut (.I0(n69070), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n69071));   // verilog/uart_rx.v(119[33:55])
    defparam i53345_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2790_7 (.CI(n51366), .I0(n2105), .I1(n1459), .CO(n51367));
    SB_CARRY add_2798_14 (.CI(n51504), .I0(n3055), .I1(n2272), .CO(n51505));
    SB_LUT4 add_2790_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n51365), 
            .O(n8185[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_12 (.CI(n51445), .I0(n2721), .I1(n2013), .CO(n51446));
    SB_LUT4 i53016_3_lut (.I0(n69071), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i53016_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2790_6 (.CI(n51365), .I0(n2106), .I1(n1460), .CO(n51366));
    SB_LUT4 add_2795_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n51444), 
            .O(n8315[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_11 (.CI(n51444), .I0(n2722), .I1(n1879), .CO(n51445));
    SB_LUT4 add_2790_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n51364), 
            .O(n8185[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n50433), .I0(n294[2]), .I1(VCC_net), 
            .CO(n50434));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n50432), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n50432), .I0(n294[1]), .I1(VCC_net), 
            .CO(n50433));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n60390), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n60390), .I1(GND_net), 
            .CO(n50432));
    SB_CARRY add_2790_5 (.CI(n51364), .I0(n2107), .I1(n1011), .CO(n51365));
    SB_LUT4 add_2790_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n51363), 
            .O(n8185[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_985 (.I0(n68397), .I1(baudrate[21]), .I2(n3046), 
            .I3(n61364), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_985.LUT_INIT = 16'h7100;
    SB_LUT4 i54389_2_lut_4_lut (.I0(n68397), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25651), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i54389_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2798_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n51503), 
            .O(n8393[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_986 (.I0(n69269), .I1(baudrate[20]), .I2(n2938), 
            .I3(n61362), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_986.LUT_INIT = 16'h7100;
    SB_LUT4 i54384_2_lut_4_lut (.I0(n69269), .I1(baudrate[20]), .I2(n2938), 
            .I3(n63601), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i54384_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2795_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n51443), 
            .O(n8315[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_4 (.CI(n51363), .I0(n2108), .I1(n856), .CO(n51364));
    SB_LUT4 i47883_1_lut (.I0(n63599), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59108));
    defparam i47883_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8289[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8315[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8341[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2790_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n51362), 
            .O(n8185[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8133[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8289[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5753_2_lut_3_lut_4_lut_4_lut (.I0(baudrate[3]), .I1(n20844), 
            .I2(n11422), .I3(n960), .O(n44_adj_5011));   // verilog/uart_rx.v(119[33:55])
    defparam i5753_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd54;
    SB_LUT4 i54209_4_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(n6_adj_5095), .I3(n61043), .O(n58988));
    defparam i54209_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_CARRY add_2798_13 (.CI(n51503), .I0(n3056), .I1(n2144), .CO(n51504));
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_4994), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8315[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8341[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2795_10 (.CI(n51443), .I0(n2723), .I1(n1742), .CO(n51444));
    SB_CARRY add_2790_3 (.CI(n51362), .I0(n2109), .I1(n698), .CO(n51363));
    SB_LUT4 i1_2_lut_4_lut_adj_987 (.I0(n69146), .I1(baudrate[17]), .I2(n2596), 
            .I3(n61356), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_987.LUT_INIT = 16'h7100;
    SB_LUT4 i54364_2_lut_4_lut (.I0(n69146), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25639), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i54364_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2790_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8185[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n51442), 
            .O(n8315[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n51362));
    SB_LUT4 add_2789_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n51361), 
            .O(n8159[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_988 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n62772));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_989 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n62770));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_990 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n62774));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_991 (.I0(n68967), .I1(baudrate[18]), .I2(n2713), 
            .I3(n61358), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_991.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_adj_992 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n62768));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28519_rep_5_2_lut (.I0(n8081[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n59102));   // verilog/uart_rx.v(119[33:55])
    defparam i28519_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n59102), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52848_3_lut (.I0(n32_adj_5126), .I1(baudrate[6]), .I2(n39_adj_5124), 
            .I3(GND_net), .O(n68574));   // verilog/uart_rx.v(119[33:55])
    defparam i52848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52849_3_lut (.I0(n68574), .I1(baudrate[7]), .I2(n41_adj_5123), 
            .I3(GND_net), .O(n68575));   // verilog/uart_rx.v(119[33:55])
    defparam i52849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52288_4_lut (.I0(n41_adj_5123), .I1(n39_adj_5124), .I2(n37_adj_5125), 
            .I3(n67155), .O(n68014));
    defparam i52288_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52959_3_lut (.I0(n34), .I1(baudrate[5]), .I2(n37_adj_5125), 
            .I3(GND_net), .O(n68685));   // verilog/uart_rx.v(119[33:55])
    defparam i52959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52102_3_lut (.I0(n68575), .I1(baudrate[8]), .I2(n43_adj_5122), 
            .I3(GND_net), .O(n67828));   // verilog/uart_rx.v(119[33:55])
    defparam i52102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54372_2_lut_4_lut (.I0(n68967), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25642), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i54372_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i53145_4_lut (.I0(n67828), .I1(n68685), .I2(n43_adj_5122), 
            .I3(n68014), .O(n68871));   // verilog/uart_rx.v(119[33:55])
    defparam i53145_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53146_3_lut (.I0(n68871), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n68872));   // verilog/uart_rx.v(119[33:55])
    defparam i53146_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n68872), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_993 (.I0(n62814), .I1(n62770), .I2(n62772), .I3(baudrate[11]), 
            .O(n62800));
    defparam i1_4_lut_adj_993.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_994 (.I0(n62800), .I1(n62802), .I2(n62790), .I3(n62724), 
            .O(n25618));
    defparam i1_4_lut_adj_994.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n25618), .I1(n48_adj_5127), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8081[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8107[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8081[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8107[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8081[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8107[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8081[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8081[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8107[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8081[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8107[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8107[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8107[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51411_4_lut (.I0(n35_adj_5134), .I1(n33_adj_5133), .I2(n31_adj_5132), 
            .I3(n29_adj_5135), .O(n67137));
    defparam i51411_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5136), .I1(baudrate[9]), 
            .I2(n43_adj_5130), .I3(GND_net), .O(n40_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52846_3_lut (.I0(n28_adj_5138), .I1(baudrate[5]), .I2(n35_adj_5134), 
            .I3(GND_net), .O(n68572));   // verilog/uart_rx.v(119[33:55])
    defparam i52846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52847_3_lut (.I0(n68572), .I1(baudrate[6]), .I2(n37_adj_5129), 
            .I3(GND_net), .O(n68573));   // verilog/uart_rx.v(119[33:55])
    defparam i52847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51405_4_lut (.I0(n41_adj_5131), .I1(n39_adj_5128), .I2(n37_adj_5129), 
            .I3(n67137), .O(n67131));
    defparam i51405_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53302_4_lut (.I0(n40_adj_5137), .I1(n30_adj_5139), .I2(n43_adj_5130), 
            .I3(n67129), .O(n69028));   // verilog/uart_rx.v(119[33:55])
    defparam i53302_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52107_3_lut (.I0(n68573), .I1(baudrate[7]), .I2(n39_adj_5128), 
            .I3(GND_net), .O(n67833));   // verilog/uart_rx.v(119[33:55])
    defparam i52107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53484_4_lut (.I0(n67833), .I1(n69028), .I2(n43_adj_5130), 
            .I3(n67131), .O(n69210));   // verilog/uart_rx.v(119[33:55])
    defparam i53484_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53485_3_lut (.I0(n69210), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n69211));   // verilog/uart_rx.v(119[33:55])
    defparam i53485_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8159[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8185[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8211[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8237[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8263[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n856), .I1(n42_adj_5140), .I2(baudrate[4]), 
            .I3(n20846), .O(n59555));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff8f;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8289[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8315[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8341[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2789_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n51360), 
            .O(n8159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n51502), 
            .O(n8393[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_995 (.I0(n698), .I1(n42_adj_5141), .I2(baudrate[3]), 
            .I3(n20836), .O(n59595));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_995.LUT_INIT = 16'hff8f;
    SB_CARRY add_2795_9 (.CI(n51442), .I0(n2724), .I1(n1602), .CO(n51443));
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8159[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8263[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8289[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8315[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2789_13 (.CI(n51360), .I0(n1967), .I1(n2144), .CO(n51361));
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8341[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2795_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n51441), 
            .O(n8315[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2789_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n51359), 
            .O(n8159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_12 (.CI(n51359), .I0(n1968), .I1(n2013), .CO(n51360));
    SB_LUT4 add_2789_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n51358), 
            .O(n8159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_11 (.CI(n51358), .I0(n1969), .I1(n1879), .CO(n51359));
    SB_CARRY add_2795_8 (.CI(n51441), .I0(n2725), .I1(n1459), .CO(n51442));
    SB_CARRY add_2798_12 (.CI(n51502), .I0(n3057), .I1(n2013), .CO(n51503));
    SB_LUT4 add_2789_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n51357), 
            .O(n8159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n51440), 
            .O(n8315[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_10 (.CI(n51357), .I0(n1970), .I1(n1742), .CO(n51358));
    SB_LUT4 add_2798_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n51501), 
            .O(n8393[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_7 (.CI(n51440), .I0(n2726), .I1(n1460), .CO(n51441));
    SB_LUT4 add_2795_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n51439), 
            .O(n8315[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2789_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n51356), 
            .O(n8159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_9 (.CI(n51356), .I0(n1971), .I1(n1602), .CO(n51357));
    SB_LUT4 add_2789_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n51355), 
            .O(n8159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_8 (.CI(n51355), .I0(n1972), .I1(n1459), .CO(n51356));
    SB_LUT4 add_2789_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n51354), 
            .O(n8159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_11 (.CI(n51501), .I0(n3058), .I1(n1879), .CO(n51502));
    SB_CARRY add_2795_6 (.CI(n51439), .I0(n2727), .I1(n1011), .CO(n51440));
    SB_CARRY add_2789_7 (.CI(n51354), .I0(n1973), .I1(n1460), .CO(n51355));
    SB_LUT4 add_2795_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n51438), 
            .O(n8315[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2789_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n51353), 
            .O(n8159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_6 (.CI(n51353), .I0(n1974), .I1(n1011), .CO(n51354));
    SB_LUT4 i1_2_lut_4_lut_adj_996 (.I0(n69259), .I1(baudrate[19]), .I2(n2827), 
            .I3(n61360), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_996.LUT_INIT = 16'h7100;
    SB_LUT4 add_2789_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n51352), 
            .O(n8159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54379_2_lut_4_lut (.I0(n69259), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25645), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i54379_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut_adj_997 (.I0(n61852), .I1(n63605), .I2(baudrate[0]), 
            .I3(n48_adj_5142), .O(n962));
    defparam i1_3_lut_4_lut_adj_997.LUT_INIT = 16'h0010;
    SB_CARRY add_2795_5 (.CI(n51438), .I0(n2728), .I1(n856), .CO(n51439));
    SB_LUT4 add_2798_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n51500), 
            .O(n8393[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_10 (.CI(n51500), .I0(n3059), .I1(n1742), .CO(n51501));
    SB_LUT4 add_2795_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n51437), 
            .O(n8315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8263[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2795_4 (.CI(n51437), .I0(n2729), .I1(n698), .CO(n51438));
    SB_CARRY add_2789_5 (.CI(n51352), .I0(n1975), .I1(n856), .CO(n51353));
    SB_LUT4 add_2789_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n51351), 
            .O(n8159[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n51499), 
            .O(n8393[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_9 (.CI(n51499), .I0(n3060), .I1(n1602), .CO(n51500));
    SB_LUT4 add_2795_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n51436), 
            .O(n8315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_4 (.CI(n51351), .I0(n1976), .I1(n698), .CO(n51352));
    SB_LUT4 add_2789_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n51350), 
            .O(n8159[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_3 (.CI(n51350), .I0(n1977), .I1(n858), .CO(n51351));
    SB_LUT4 add_2789_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8159[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n51498), 
            .O(n8393[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51350));
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8289[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2795_3 (.CI(n51436), .I0(n2730), .I1(n858), .CO(n51437));
    SB_LUT4 add_2788_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n51349), 
            .O(n8133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8315[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2795_2_lut (.I0(n59074), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61358)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2788_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n51348), 
            .O(n8133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_8 (.CI(n51498), .I0(n3061), .I1(n1459), .CO(n51499));
    SB_CARRY add_2795_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51436));
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8341[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2788_12 (.CI(n51348), .I0(n1832), .I1(n2013), .CO(n51349));
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8263[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8289[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8315[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2788_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n51347), 
            .O(n8133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_11 (.CI(n51347), .I0(n1833), .I1(n1879), .CO(n51348));
    SB_LUT4 add_2794_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n51435), 
            .O(n8289[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n51497), 
            .O(n8393[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2788_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n51346), 
            .O(n8133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n51434), 
            .O(n8289[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_10 (.CI(n51346), .I0(n1834), .I1(n1742), .CO(n51347));
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8185[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8341[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2798_7 (.CI(n51497), .I0(n3062), .I1(n1460), .CO(n51498));
    SB_LUT4 i1_3_lut_4_lut_adj_998 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61750));
    defparam i1_3_lut_4_lut_adj_998.LUT_INIT = 16'hfff7;
    SB_LUT4 add_2788_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n51345), 
            .O(n8133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n51496), 
            .O(n8393[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_18 (.CI(n51434), .I0(n2597), .I1(n2754), .CO(n51435));
    SB_CARRY add_2788_9 (.CI(n51345), .I0(n1835), .I1(n1602), .CO(n51346));
    SB_LUT4 add_2788_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n51344), 
            .O(n8133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8263[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2794_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n51433), 
            .O(n8289[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_8 (.CI(n51344), .I0(n1836), .I1(n1459), .CO(n51345));
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8289[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2788_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n51343), 
            .O(n8133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8315[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8341[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_999 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61702));
    defparam i1_3_lut_4_lut_adj_999.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_3_lut_4_lut_adj_1000 (.I0(n62726), .I1(n63577), .I2(n8081[14]), 
            .I3(n48_adj_5144), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1000.LUT_INIT = 16'h0010;
    SB_CARRY add_2788_7 (.CI(n51343), .I0(n1837), .I1(n1460), .CO(n51344));
    SB_LUT4 i1_3_lut_4_lut_adj_1001 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61734));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1001.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1002 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61814));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1002.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut_4_lut_adj_1003 (.I0(n61844), .I1(n63391), .I2(n8159[11]), 
            .I3(n48_adj_5145), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1003.LUT_INIT = 16'h0010;
    SB_LUT4 i47860_2_lut_3_lut (.I0(n61844), .I1(n63391), .I2(baudrate[12]), 
            .I3(GND_net), .O(n63577));
    defparam i47860_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i54348_2_lut_3_lut (.I0(n61844), .I1(n63391), .I2(n48_adj_5145), 
            .I3(GND_net), .O(n294[11]));
    defparam i54348_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_1004 (.I0(n62828), .I1(n61320), .I2(n61318), 
            .I3(n62818), .O(n25639));
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'hfffe;
    SB_LUT4 i43400_1_lut (.I0(n25639), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59078));
    defparam i43400_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8263[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2798_6 (.CI(n51496), .I0(n3063), .I1(n1011), .CO(n51497));
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8289[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2794_17 (.CI(n51433), .I0(n2598), .I1(n2638), .CO(n51434));
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8315[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8341[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2788_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n51342), 
            .O(n8133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2794_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n51432), 
            .O(n8289[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_6 (.CI(n51342), .I0(n1838), .I1(n1011), .CO(n51343));
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2788_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n51341), 
            .O(n8133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8237[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8237[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28498_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42420));
    defparam i28498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_2794_16 (.CI(n51432), .I0(n2599), .I1(n2519), .CO(n51433));
    SB_CARRY add_2788_5 (.CI(n51341), .I0(n1839), .I1(n856), .CO(n51342));
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8211[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1952_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n51696), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1952_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n51695), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1952_add_4_8 (.CI(n51695), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n51696));
    SB_LUT4 r_Clock_Count_1952_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n51694), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8237[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2794_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n51431), 
            .O(n8289[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2788_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n51340), 
            .O(n8133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_4 (.CI(n51340), .I0(n1840), .I1(n698), .CO(n51341));
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8237[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8237[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY r_Clock_Count_1952_add_4_7 (.CI(n51694), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n51695));
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2794_15 (.CI(n51431), .I0(n2600), .I1(n2397), .CO(n51432));
    SB_LUT4 r_Clock_Count_1952_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n51693), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2788_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n51339), 
            .O(n8133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_3 (.CI(n51339), .I0(n1841), .I1(n858), .CO(n51340));
    SB_LUT4 add_2794_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n51430), 
            .O(n8289[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2788_2_lut (.I0(n59099), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61348)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2788_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51339));
    SB_LUT4 add_2787_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n51338), 
            .O(n8107[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2787_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n51337), 
            .O(n8107[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_14 (.CI(n51430), .I0(n2601), .I1(n2272), .CO(n51431));
    SB_LUT4 add_2794_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n51429), 
            .O(n8289[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n51495), 
            .O(n8393[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_13 (.CI(n51429), .I0(n2602), .I1(n2144), .CO(n51430));
    SB_LUT4 add_2794_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n51428), 
            .O(n8289[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_5 (.CI(n51495), .I0(n3064), .I1(n856), .CO(n51496));
    SB_LUT4 add_2798_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n51494), 
            .O(n8393[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_10 (.CI(n51337), .I0(n1694), .I1(n1879), .CO(n51338));
    SB_CARRY r_Clock_Count_1952_add_4_6 (.CI(n51693), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n51694));
    SB_LUT4 add_2787_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n51336), 
            .O(n8107[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_12 (.CI(n51428), .I0(n2603), .I1(n2013), .CO(n51429));
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51303_4_lut (.I0(n25_adj_5154), .I1(n23_adj_5153), .I2(n21_adj_5152), 
            .I3(n19_adj_5159), .O(n67029));
    defparam i51303_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2787_9 (.CI(n51336), .I0(n1695), .I1(n1742), .CO(n51337));
    SB_LUT4 add_2787_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n51335), 
            .O(n8107[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n51427), 
            .O(n8289[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51297_4_lut (.I0(n31_adj_5151), .I1(n29_adj_5150), .I2(n27_adj_5155), 
            .I3(n67029), .O(n67023));
    defparam i51297_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53027_4_lut (.I0(n37_adj_5158), .I1(n35_adj_5157), .I2(n33_adj_5156), 
            .I3(n67023), .O(n68753));
    defparam i53027_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2798_4 (.CI(n51494), .I0(n3065), .I1(n698), .CO(n51495));
    SB_CARRY add_2794_11 (.CI(n51427), .I0(n2604), .I1(n1879), .CO(n51428));
    SB_CARRY add_2787_8 (.CI(n51335), .I0(n1696), .I1(n1602), .CO(n51336));
    SB_LUT4 add_2787_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n51334), 
            .O(n8107[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1952_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n51692), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_7 (.CI(n51334), .I0(n1697), .I1(n1459), .CO(n51335));
    SB_LUT4 add_2787_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n51333), 
            .O(n8107[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_6 (.CI(n51333), .I0(n1698), .I1(n1460), .CO(n51334));
    SB_LUT4 add_2798_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n51493), 
            .O(n8393[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n51426), 
            .O(n8289[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2787_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n51332), 
            .O(n8107[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_10 (.CI(n51426), .I0(n2605), .I1(n1742), .CO(n51427));
    SB_LUT4 i52817_3_lut (.I0(n18_adj_5160), .I1(baudrate[13]), .I2(n41_adj_5149), 
            .I3(GND_net), .O(n68543));   // verilog/uart_rx.v(119[33:55])
    defparam i52817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52818_3_lut (.I0(n68543), .I1(baudrate[14]), .I2(n43_adj_5148), 
            .I3(GND_net), .O(n68544));   // verilog/uart_rx.v(119[33:55])
    defparam i52818_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2787_5 (.CI(n51332), .I0(n1699), .I1(n1011), .CO(n51333));
    SB_CARRY add_2798_3 (.CI(n51493), .I0(n3066), .I1(n858), .CO(n51494));
    SB_LUT4 i52166_4_lut (.I0(n43_adj_5148), .I1(n41_adj_5149), .I2(n29_adj_5150), 
            .I3(n67025), .O(n67892));
    defparam i52166_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5161), .I1(baudrate[7]), 
            .I2(n29_adj_5150), .I3(GND_net), .O(n26_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2798_2_lut (.I0(n59062), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61364)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2794_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n51425), 
            .O(n8289[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1952_add_4_5 (.CI(n51692), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n51693));
    SB_CARRY add_2794_9 (.CI(n51425), .I0(n2606), .I1(n1602), .CO(n51426));
    SB_CARRY add_2798_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51493));
    SB_LUT4 add_2794_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n51424), 
            .O(n8289[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52147_3_lut (.I0(n68544), .I1(baudrate[15]), .I2(n45_adj_5147), 
            .I3(GND_net), .O(n67873));   // verilog/uart_rx.v(119[33:55])
    defparam i52147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1952_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n51691), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1952_add_4_4 (.CI(n51691), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n51692));
    SB_LUT4 add_2787_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n51331), 
            .O(n8107[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1952_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n51690), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1952_add_4_3 (.CI(n51690), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n51691));
    SB_LUT4 r_Clock_Count_1952_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1952_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1952_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n51690));
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5163), .I1(baudrate[9]), 
            .I2(n33_adj_5156), .I3(GND_net), .O(n30_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53334_4_lut (.I0(n30_adj_5164), .I1(n20_adj_5165), .I2(n33_adj_5156), 
            .I3(n67019), .O(n69060));   // verilog/uart_rx.v(119[33:55])
    defparam i53334_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53335_3_lut (.I0(n69060), .I1(baudrate[10]), .I2(n35_adj_5157), 
            .I3(GND_net), .O(n69061));   // verilog/uart_rx.v(119[33:55])
    defparam i53335_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2787_4 (.CI(n51331), .I0(n1700), .I1(n856), .CO(n51332));
    SB_LUT4 add_2797_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n51492), 
            .O(n8367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53128_3_lut (.I0(n69061), .I1(baudrate[11]), .I2(n37_adj_5158), 
            .I3(GND_net), .O(n68854));   // verilog/uart_rx.v(119[33:55])
    defparam i53128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52168_4_lut (.I0(n43_adj_5148), .I1(n41_adj_5149), .I2(n39_adj_5146), 
            .I3(n68753), .O(n67894));
    defparam i52168_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52975_4_lut (.I0(n67873), .I1(n26_adj_5162), .I2(n45_adj_5147), 
            .I3(n67892), .O(n68701));   // verilog/uart_rx.v(119[33:55])
    defparam i52975_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52145_3_lut (.I0(n68854), .I1(baudrate[12]), .I2(n39_adj_5146), 
            .I3(GND_net), .O(n67871));   // verilog/uart_rx.v(119[33:55])
    defparam i52145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1005 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61782));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1005.LUT_INIT = 16'hfffd;
    SB_LUT4 add_2787_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n51330), 
            .O(n8107[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n51491), 
            .O(n8367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_3 (.CI(n51330), .I0(n1701), .I1(n698), .CO(n51331));
    SB_LUT4 i52977_4_lut (.I0(n67871), .I1(n68701), .I2(n45_adj_5147), 
            .I3(n67894), .O(n68703));   // verilog/uart_rx.v(119[33:55])
    defparam i52977_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_4_lut_adj_1006 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61766));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1006.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1007 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61798));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1007.LUT_INIT = 16'hffef;
    SB_LUT4 i1_3_lut_4_lut_adj_1008 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5143), .O(n61718));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1008.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8237[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8263[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2797_21 (.CI(n51491), .I0(n2939), .I1(n3084), .CO(n51492));
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8289[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8315[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8341[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28496_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42418));
    defparam i28496_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8211[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8237[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8211[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51007_2_lut (.I0(baudrate[1]), .I1(n294[20]), .I2(GND_net), 
            .I3(GND_net), .O(n66733));   // verilog/uart_rx.v(119[33:55])
    defparam i51007_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8211[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51581_4_lut (.I0(n25593), .I1(n66733), .I2(n48_adj_5170), 
            .I3(baudrate[0]), .O(n804));
    defparam i51581_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8211[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43384_1_lut (.I0(n25651), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59062));
    defparam i43384_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8211[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8263[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8289[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8211[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8055[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8315[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51325_4_lut (.I0(n27_adj_5176), .I1(n25_adj_5175), .I2(n23_adj_5174), 
            .I3(n21_adj_5177), .O(n67051));
    defparam i51325_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51321_4_lut (.I0(n33_adj_5173), .I1(n31_adj_5172), .I2(n29_adj_5171), 
            .I3(n67051), .O(n67047));
    defparam i51321_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5179), .I1(baudrate[7]), 
            .I2(n31_adj_5172), .I3(GND_net), .O(n28_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5182), .I1(baudrate[9]), 
            .I2(n35_adj_5169), .I3(GND_net), .O(n32_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53332_4_lut (.I0(n32_adj_5183), .I1(n22_adj_5184), .I2(n35_adj_5169), 
            .I3(n67045), .O(n69058));   // verilog/uart_rx.v(119[33:55])
    defparam i53332_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n62012));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n62818));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'heeee;
    SB_LUT4 i53333_3_lut (.I0(n69058), .I1(baudrate[10]), .I2(n37_adj_5168), 
            .I3(GND_net), .O(n69059));   // verilog/uart_rx.v(119[33:55])
    defparam i53333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n62012), .I1(n62828), .I2(n62772), 
            .I3(n62768), .O(n25645));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 i53130_3_lut (.I0(n69059), .I1(baudrate[11]), .I2(n39_adj_5167), 
            .I3(GND_net), .O(n68856));   // verilog/uart_rx.v(119[33:55])
    defparam i53130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n62820));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'heeee;
    SB_LUT4 i51132_4_lut (.I0(n35_adj_4995), .I1(n23_adj_4998), .I2(n21), 
            .I3(n19), .O(n66858));
    defparam i51132_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53031_4_lut (.I0(n39_adj_5167), .I1(n37_adj_5168), .I2(n35_adj_5169), 
            .I3(n67047), .O(n68757));
    defparam i53031_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53397_4_lut (.I0(n28_adj_5180), .I1(n20_adj_5178), .I2(n31_adj_5172), 
            .I3(n67049), .O(n69123));   // verilog/uart_rx.v(119[33:55])
    defparam i53397_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52139_3_lut (.I0(n68856), .I1(baudrate[12]), .I2(n41_adj_5166), 
            .I3(GND_net), .O(n67865));   // verilog/uart_rx.v(119[33:55])
    defparam i52139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53482_4_lut (.I0(n67865), .I1(n69123), .I2(n41_adj_5166), 
            .I3(n68757), .O(n69208));   // verilog/uart_rx.v(119[33:55])
    defparam i53482_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53483_3_lut (.I0(n69208), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n69209));   // verilog/uart_rx.v(119[33:55])
    defparam i53483_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53462_3_lut (.I0(n69209), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n69188));   // verilog/uart_rx.v(119[33:55])
    defparam i53462_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52047_4_lut (.I0(n17), .I1(n15), .I2(n2844), .I3(baudrate[2]), 
            .O(n67773));
    defparam i52047_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n62730));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'heeee;
    SB_LUT4 i52625_4_lut (.I0(n23_adj_4998), .I1(n21), .I2(n19), .I3(n67773), 
            .O(n68351));
    defparam i52625_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n62728));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8263[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52623_4_lut (.I0(n29_adj_5010), .I1(n27_adj_5009), .I2(n25_adj_5001), 
            .I3(n68351), .O(n68349));
    defparam i52623_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i5744_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11422));   // verilog/uart_rx.v(119[33:55])
    defparam i5744_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8185[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8185[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8185[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8055[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47888_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), .I2(n63599), 
            .I3(GND_net), .O(n63605));
    defparam i47888_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i47861_1_lut (.I0(n63577), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59099));
    defparam i47861_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8185[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8055[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51152_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n66878));
    defparam i51152_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8185[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8185[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51352_4_lut (.I0(n29_adj_5195), .I1(n27_adj_5193), .I2(n25_adj_5190), 
            .I3(n23_adj_5200), .O(n67078));
    defparam i51352_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51348_4_lut (.I0(n35_adj_5199), .I1(n33_adj_5198), .I2(n31_adj_5197), 
            .I3(n67078), .O(n67074));
    defparam i51348_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8055[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5202), .I1(baudrate[7]), 
            .I2(n33_adj_5198), .I3(GND_net), .O(n30_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5205), .I1(baudrate[9]), 
            .I2(n37_adj_5189), .I3(GND_net), .O(n34_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53330_4_lut (.I0(n34_adj_5206), .I1(n24_adj_5207), .I2(n37_adj_5189), 
            .I3(n67072), .O(n69056));   // verilog/uart_rx.v(119[33:55])
    defparam i53330_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53331_3_lut (.I0(n69056), .I1(baudrate[10]), .I2(n39_adj_5187), 
            .I3(GND_net), .O(n69057));   // verilog/uart_rx.v(119[33:55])
    defparam i53331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53132_3_lut (.I0(n69057), .I1(baudrate[11]), .I2(n41_adj_5188), 
            .I3(GND_net), .O(n68858));   // verilog/uart_rx.v(119[33:55])
    defparam i53132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53033_4_lut (.I0(n41_adj_5188), .I1(n39_adj_5187), .I2(n37_adj_5189), 
            .I3(n67074), .O(n68759));
    defparam i53033_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8029[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53227_4_lut (.I0(n30_adj_5203), .I1(n22_adj_5201), .I2(n33_adj_5198), 
            .I3(n67076), .O(n68953));   // verilog/uart_rx.v(119[33:55])
    defparam i53227_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52133_3_lut (.I0(n68858), .I1(baudrate[12]), .I2(n43_adj_5186), 
            .I3(GND_net), .O(n67859));   // verilog/uart_rx.v(119[33:55])
    defparam i52133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53300_4_lut (.I0(n67859), .I1(n68953), .I2(n43_adj_5186), 
            .I3(n68759), .O(n69026));   // verilog/uart_rx.v(119[33:55])
    defparam i53300_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53301_3_lut (.I0(n69026), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n69027));   // verilog/uart_rx.v(119[33:55])
    defparam i53301_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47651_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25639), .I3(GND_net), .O(n59086));
    defparam i47651_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_3_lut (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n4_adj_5143));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8237[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8263[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8029[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47650_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), .I2(n25639), 
            .I3(GND_net), .O(n63361));
    defparam i47650_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i47826_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n63543));
    defparam i47826_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8029[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n62710));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8029[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47889_1_lut_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), 
            .I2(n63599), .I3(GND_net), .O(n59116));
    defparam i47889_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51122_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n66848));
    defparam i51122_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i47681_1_lut_2_lut (.I0(baudrate[15]), .I1(n63361), .I2(GND_net), 
            .I3(GND_net), .O(n59090));
    defparam i47681_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52854_3_lut (.I0(n34_adj_5213), .I1(baudrate[5]), .I2(n41_adj_5211), 
            .I3(GND_net), .O(n68580));   // verilog/uart_rx.v(119[33:55])
    defparam i52854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52855_3_lut (.I0(n68580), .I1(baudrate[6]), .I2(n43_adj_5210), 
            .I3(GND_net), .O(n68581));   // verilog/uart_rx.v(119[33:55])
    defparam i52855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52306_4_lut (.I0(n43_adj_5210), .I1(n41_adj_5211), .I2(n39_adj_5209), 
            .I3(n67173), .O(n68032));
    defparam i52306_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5215), .I1(baudrate[4]), 
            .I2(n39_adj_5209), .I3(GND_net), .O(n38_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8185[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8211[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8237[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8263[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52091_3_lut (.I0(n68581), .I1(baudrate[7]), .I2(n45_adj_5208), 
            .I3(GND_net), .O(n67817));   // verilog/uart_rx.v(119[33:55])
    defparam i52091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8289[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8315[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52951_4_lut (.I0(n67817), .I1(n38_adj_5216), .I2(n45_adj_5208), 
            .I3(n68032), .O(n68677));   // verilog/uart_rx.v(119[33:55])
    defparam i52951_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8341[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8003[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8003[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5218), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n61870));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'heeee;
    SB_LUT4 i51381_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n67107));
    defparam i51381_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8159[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8159[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51578_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i51578_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8159[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8159[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8159[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8159[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47842_2_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), .I2(baudrate[12]), 
            .I3(baudrate[13]), .O(n63559));
    defparam i47842_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8159[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51370_4_lut (.I0(n33_adj_5228), .I1(n31_adj_5227), .I2(n29_adj_5226), 
            .I3(n27_adj_5229), .O(n67096));
    defparam i51370_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5230), .I1(baudrate[10]), 
            .I2(n41_adj_5224), .I3(GND_net), .O(n38_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28530_rep_4_2_lut (.I0(n8159[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n59093));   // verilog/uart_rx.v(119[33:55])
    defparam i28530_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n59093), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52840_3_lut (.I0(n26_adj_5232), .I1(baudrate[6]), .I2(n33_adj_5228), 
            .I3(GND_net), .O(n68566));   // verilog/uart_rx.v(119[33:55])
    defparam i52840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52841_3_lut (.I0(n68566), .I1(baudrate[7]), .I2(n35_adj_5223), 
            .I3(GND_net), .O(n68567));   // verilog/uart_rx.v(119[33:55])
    defparam i52841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51364_4_lut (.I0(n39_adj_5225), .I1(n37_adj_5222), .I2(n35_adj_5223), 
            .I3(n67096), .O(n67090));
    defparam i51364_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(n62814), .I1(n62700), .I2(n61870), 
            .I3(baudrate[19]), .O(n61890));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'hfffe;
    SB_LUT4 i53328_4_lut (.I0(n38_adj_5231), .I1(n28_adj_5233), .I2(n41_adj_5224), 
            .I3(n67088), .O(n69054));   // verilog/uart_rx.v(119[33:55])
    defparam i53328_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(n61890), .I1(n62774), .I2(n62816), 
            .I3(n62772), .O(n25642));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'hfffe;
    SB_LUT4 i43396_1_lut (.I0(n25642), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59074));
    defparam i43396_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52123_3_lut (.I0(n68567), .I1(baudrate[8]), .I2(n37_adj_5222), 
            .I3(GND_net), .O(n67849));   // verilog/uart_rx.v(119[33:55])
    defparam i52123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53494_4_lut (.I0(n67849), .I1(n69054), .I2(n41_adj_5224), 
            .I3(n67090), .O(n69220));   // verilog/uart_rx.v(119[33:55])
    defparam i53494_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51362_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n67088));
    defparam i51362_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i53495_3_lut (.I0(n69220), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n69221));   // verilog/uart_rx.v(119[33:55])
    defparam i53495_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53430_3_lut (.I0(n69221), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n69156));   // verilog/uart_rx.v(119[33:55])
    defparam i53430_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52129_3_lut (.I0(n69156), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam i52129_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n62824));
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1019 (.I0(n62774), .I1(n62822), .I2(n61870), 
            .I3(GND_net), .O(n62832));
    defparam i1_3_lut_adj_1019.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1020 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n62828));
    defparam i1_2_lut_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(n62832), .I1(n62828), .I2(n62830), 
            .I3(n62824), .O(n25627));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1022 (.I0(n25627), .I1(n48_adj_5234), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1022.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8211[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5236), .I1(baudrate[4]), 
            .I2(n43_adj_5219), .I3(GND_net), .O(n42_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8237[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53304_4_lut (.I0(n42_adj_5237), .I1(n38_adj_5235), .I2(n43_adj_5219), 
            .I3(n67186), .O(n69030));   // verilog/uart_rx.v(119[33:55])
    defparam i53304_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8263[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51626_2_lut_3_lut (.I0(n25593), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n66393));   // verilog/uart_rx.v(119[33:55])
    defparam i51626_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53305_3_lut (.I0(n69030), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n69031));   // verilog/uart_rx.v(119[33:55])
    defparam i53305_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51346_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n67072));
    defparam i51346_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54327_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n63605), .I3(n48_adj_5142), .O(n294[19]));
    defparam i54327_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51350_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n67076));
    defparam i51350_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n62700));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62814));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n62916));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n62918));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n62816));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1028 (.I0(n62822), .I1(n62818), .I2(n62820), 
            .I3(n62816), .O(n62802));
    defparam i1_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1029 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n62830));
    defparam i1_2_lut_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51319_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n67045));
    defparam i51319_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51323_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n67049));
    defparam i51323_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5575_2_lut_3_lut (.I0(n20834), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam i5575_2_lut_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i7130_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n20834));   // verilog/uart_rx.v(119[33:55])
    defparam i7130_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(n62916), .I1(n62710), .I2(n62814), 
            .I3(n62700), .O(n25651));
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'hfffe;
    SB_LUT4 i28503_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59119));   // verilog/uart_rx.v(119[33:55])
    defparam i28503_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n59119), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52862_3_lut (.I0(n42_adj_5238), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n68588));   // verilog/uart_rx.v(119[33:55])
    defparam i52862_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52863_3_lut (.I0(n68588), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n68589));   // verilog/uart_rx.v(119[33:55])
    defparam i52863_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n68589), .I1(baudrate[5]), 
            .I2(n58836), .I3(GND_net), .O(n48_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(n63557), .I1(n25651), .I2(n62802), 
            .I3(n63559), .O(n25603));
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1032 (.I0(n25603), .I1(n48_adj_5239), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1032.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8003[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51293_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n67019));
    defparam i51293_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51299_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n67025));
    defparam i51299_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8159[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8185[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8211[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1033 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n61320));
    defparam i1_3_lut_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5241), .I1(baudrate[4]), 
            .I2(n41_adj_5217), .I3(GND_net), .O(n40_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54342_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n63577), .I3(n48_adj_5144), .O(n294[14]));
    defparam i54342_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i53324_4_lut (.I0(n40_adj_5242), .I1(n36_adj_5240), .I2(n41_adj_5217), 
            .I3(n67179), .O(n69050));   // verilog/uart_rx.v(119[33:55])
    defparam i53324_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53325_3_lut (.I0(n69050), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n69051));   // verilog/uart_rx.v(119[33:55])
    defparam i53325_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53154_3_lut (.I0(n69051), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n68880));   // verilog/uart_rx.v(119[33:55])
    defparam i53154_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8237[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47882_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n63577), .I3(baudrate[9]), .O(n63599));
    defparam i47882_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8263[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8289[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8315[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8341[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8055[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51136_4_lut (.I0(n35_adj_4995), .I1(n33_adj_5036), .I2(n31_adj_5013), 
            .I3(n68349), .O(n66862));
    defparam i51136_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52852_3_lut (.I0(n32_adj_5243), .I1(baudrate[5]), .I2(n39_adj_5204), 
            .I3(GND_net), .O(n68578));   // verilog/uart_rx.v(119[33:55])
    defparam i52852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52853_3_lut (.I0(n68578), .I1(baudrate[6]), .I2(n41_adj_5196), 
            .I3(GND_net), .O(n68579));   // verilog/uart_rx.v(119[33:55])
    defparam i52853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52300_4_lut (.I0(n41_adj_5196), .I1(n39_adj_5204), .I2(n37_adj_5192), 
            .I3(n67165), .O(n68026));
    defparam i52300_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52957_3_lut (.I0(n34_adj_5244), .I1(baudrate[4]), .I2(n37_adj_5192), 
            .I3(GND_net), .O(n68683));   // verilog/uart_rx.v(119[33:55])
    defparam i52957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8133[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8133[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8133[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8133[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52095_3_lut (.I0(n68579), .I1(baudrate[7]), .I2(n43_adj_5185), 
            .I3(GND_net), .O(n67821));   // verilog/uart_rx.v(119[33:55])
    defparam i52095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8133[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8133[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8133[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53149_4_lut (.I0(n67821), .I1(n68683), .I2(n43_adj_5185), 
            .I3(n68026), .O(n68875));   // verilog/uart_rx.v(119[33:55])
    defparam i53149_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53150_3_lut (.I0(n68875), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n68876));   // verilog/uart_rx.v(119[33:55])
    defparam i53150_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n68876), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8133[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51391_4_lut (.I0(n33_adj_5251), .I1(n31_adj_5250), .I2(n29_adj_5249), 
            .I3(n27_adj_5252), .O(n67117));
    defparam i51391_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5221), .I1(baudrate[9]), 
            .I2(n41_adj_5247), .I3(GND_net), .O(n38_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52844_3_lut (.I0(n26_adj_5254), .I1(baudrate[5]), .I2(n33_adj_5251), 
            .I3(GND_net), .O(n68570));   // verilog/uart_rx.v(119[33:55])
    defparam i52844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52845_3_lut (.I0(n68570), .I1(baudrate[6]), .I2(n35_adj_5246), 
            .I3(GND_net), .O(n68571));   // verilog/uart_rx.v(119[33:55])
    defparam i52845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51383_4_lut (.I0(n39_adj_5248), .I1(n37_adj_5245), .I2(n35_adj_5246), 
            .I3(n67117), .O(n67109));
    defparam i51383_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53326_4_lut (.I0(n38_adj_5253), .I1(n28_adj_5220), .I2(n41_adj_5247), 
            .I3(n67107), .O(n69052));   // verilog/uart_rx.v(119[33:55])
    defparam i53326_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52111_3_lut (.I0(n68571), .I1(baudrate[7]), .I2(n37_adj_5245), 
            .I3(GND_net), .O(n67837));   // verilog/uart_rx.v(119[33:55])
    defparam i52111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53492_4_lut (.I0(n67837), .I1(n69052), .I2(n41_adj_5247), 
            .I3(n67109), .O(n69218));   // verilog/uart_rx.v(119[33:55])
    defparam i53492_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53493_3_lut (.I0(n69218), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n69219));   // verilog/uart_rx.v(119[33:55])
    defparam i53493_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53434_3_lut (.I0(n69219), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n69160));   // verilog/uart_rx.v(119[33:55])
    defparam i53434_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52117_3_lut (.I0(n69160), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam i52117_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8185[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8211[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8237[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8263[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51661_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4939), .I3(n57927), .O(n66243));
    defparam i51661_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i51639_4_lut (.I0(n66243), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n66240));
    defparam i51639_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n66240), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27722));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i54014_2_lut_4_lut (.I0(n69156), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25627), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i54014_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i5582_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(n20834), .I2(n42418), 
            .I3(n804), .O(n44));   // verilog/uart_rx.v(119[33:55])
    defparam i5582_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf45;
    SB_LUT4 i51679_2_lut (.I0(n57703), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n66301));
    defparam i51679_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51676_4_lut (.I0(n66301), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n66298));
    defparam i51676_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50953_4_lut (.I0(n66298), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n66295));
    defparam i50953_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53666_4_lut (.I0(\r_SM_Main[2] ), .I1(n66295), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(\r_SM_Main[1] ), .O(n29073));
    defparam i53666_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n57703), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n61432));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n61432), .O(n61438));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'h0100;
    SB_LUT4 i53600_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n61438), .O(n27766));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i53600_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i51403_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n67129));
    defparam i51403_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n66393), .I1(baudrate[2]), 
            .I2(n69304), .I3(n48_adj_5170), .O(n46_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1036 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n62790));
    defparam i1_2_lut_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5255), .I1(baudrate[3]), 
            .I2(n58832), .I3(GND_net), .O(n48_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53087_3_lut (.I0(n12_adj_5256), .I1(baudrate[13]), .I2(n35_adj_4995), 
            .I3(GND_net), .O(n68813));   // verilog/uart_rx.v(119[33:55])
    defparam i53087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53597_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n27845));
    defparam i53597_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i7138_4_lut_4_lut (.I0(n960), .I1(n11422), .I2(n20844), .I3(baudrate[3]), 
            .O(n20846));   // verilog/uart_rx.v(119[33:55])
    defparam i7138_4_lut_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 i54392_2_lut_4_lut (.I0(n69071), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25654), .O(n294[1]));
    defparam i54392_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50996_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n66722));
    defparam i50996_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50947_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n66673));
    defparam i50947_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51027_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n66753));
    defparam i51027_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50966_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n66692));
    defparam i50966_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i53934_2_lut_4_lut (.I0(n68872), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25618), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i53934_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51096_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n66822));
    defparam i51096_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53900_2_lut_4_lut (.I0(n68589), .I1(baudrate[5]), .I2(n58836), 
            .I3(n25603), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i53900_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51074_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n66800));
    defparam i51074_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1037 (.I0(n25593), .I1(n48_adj_5170), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5086));
    defparam i1_3_lut_4_lut_adj_1037.LUT_INIT = 16'hefff;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51003_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5170), .I2(n25593), 
            .I3(GND_net), .O(n66729));   // verilog/uart_rx.v(119[33:55])
    defparam i51003_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i53785_2_lut_4_lut (.I0(n46_adj_5255), .I1(baudrate[3]), .I2(n58832), 
            .I3(n25597), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i53785_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51241_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n66967));
    defparam i51241_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51260_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n66986));
    defparam i51260_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1038 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n61988));
    defparam i1_2_lut_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51192_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n66918));
    defparam i51192_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51169_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n66895));
    defparam i51169_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47766_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n63483));
    defparam i47766_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i47614_1_lut_2_lut (.I0(baudrate[17]), .I1(n25639), .I2(GND_net), 
            .I3(GND_net), .O(n59082));
    defparam i47614_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(n61984), .I1(n62728), .I2(n62730), 
            .I3(n62726), .O(n61996));
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1040 (.I0(n61996), .I1(n25645), .I2(n61988), 
            .I3(n62830), .O(n25597));
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i47887_1_lut_2_lut (.I0(baudrate[8]), .I1(n63599), .I2(GND_net), 
            .I3(GND_net), .O(n59112));
    defparam i47887_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_3_lut_adj_1041 (.I0(n25597), .I1(n48_adj_5257), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1041.LUT_INIT = 16'hefef;
    SB_LUT4 i51439_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n67165));   // verilog/uart_rx.v(119[33:55])
    defparam i51439_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1042 (.I0(n68880), .I1(baudrate[7]), .I2(n1261), 
            .I3(n61344), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1042.LUT_INIT = 16'h7100;
    SB_LUT4 i54336_2_lut_4_lut (.I0(n68880), .I1(baudrate[7]), .I2(n1261), 
            .I3(n63603), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i54336_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51453_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n67179));   // verilog/uart_rx.v(119[33:55])
    defparam i51453_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5214), .I1(baudrate[17]), 
            .I2(n43_adj_5181), .I3(GND_net), .O(n38_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i53088_3_lut (.I0(n68813), .I1(baudrate[14]), .I2(n37_adj_5014), 
            .I3(GND_net), .O(n68814));   // verilog/uart_rx.v(119[33:55])
    defparam i53088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1043 (.I0(n69031), .I1(baudrate[6]), .I2(n1111), 
            .I3(n61342), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1043.LUT_INIT = 16'h7100;
    SB_LUT4 i47759_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n63475));
    defparam i47759_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54330_2_lut_4_lut (.I0(n69031), .I1(baudrate[6]), .I2(n1111), 
            .I3(n63605), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i54330_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5259));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4939), 
            .O(n15_adj_5260));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5260), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5259), 
            .I3(n57927), .O(n70507));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51460_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n67186));   // verilog/uart_rx.v(119[33:55])
    defparam i51460_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i47680_2_lut (.I0(baudrate[15]), .I1(n63361), .I2(GND_net), 
            .I3(GND_net), .O(n63391));
    defparam i47680_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n61844));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'heeee;
    SB_LUT4 i51124_4_lut (.I0(n41_adj_5031), .I1(n39_adj_5026), .I2(n37_adj_5014), 
            .I3(n66858), .O(n66850));
    defparam i51124_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53085_4_lut (.I0(n38_adj_5258), .I1(n18_adj_5212), .I2(n43_adj_5181), 
            .I3(n66848), .O(n68811));   // verilog/uart_rx.v(119[33:55])
    defparam i53085_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52992_3_lut (.I0(n68814), .I1(baudrate[15]), .I2(n39_adj_5026), 
            .I3(GND_net), .O(n68718));   // verilog/uart_rx.v(119[33:55])
    defparam i52992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43380_1_lut_4_lut (.I0(n62918), .I1(n62920), .I2(n62770), 
            .I3(n62916), .O(n59058));
    defparam i43380_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_adj_1045 (.I0(n68677), .I1(baudrate[8]), .I2(n1408), 
            .I3(n61346), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1045.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_3_lut_adj_1046 (.I0(baudrate[26]), .I1(baudrate[30]), 
            .I2(baudrate[23]), .I3(GND_net), .O(n62920));
    defparam i1_2_lut_3_lut_adj_1046.LUT_INIT = 16'hfefe;
    SB_LUT4 i54339_2_lut_4_lut (.I0(n68677), .I1(baudrate[8]), .I2(n1408), 
            .I3(n63599), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i54339_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i51447_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n67173));   // verilog/uart_rx.v(119[33:55])
    defparam i51447_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1047 (.I0(n69027), .I1(baudrate[14]), .I2(n2227), 
            .I3(n61350), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1047.LUT_INIT = 16'h7100;
    SB_LUT4 i54351_2_lut_4_lut (.I0(n69027), .I1(baudrate[14]), .I2(n2227), 
            .I3(n63391), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i54351_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47886_2_lut (.I0(baudrate[8]), .I1(n63599), .I2(GND_net), 
            .I3(GND_net), .O(n63603));
    defparam i47886_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1048 (.I0(n69188), .I1(baudrate[15]), .I2(n2353), 
            .I3(n61352), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1048.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n61852));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'heeee;
    SB_LUT4 i54358_2_lut_4_lut (.I0(n69188), .I1(baudrate[15]), .I2(n2353), 
            .I3(n63361), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i54358_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5194), .I1(baudrate[9]), 
            .I2(n27_adj_5009), .I3(GND_net), .O(n24_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52866_3_lut (.I0(n42_adj_5262), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n68592));   // verilog/uart_rx.v(119[33:55])
    defparam i52866_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52867_3_lut (.I0(n68592), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n68593));   // verilog/uart_rx.v(119[33:55])
    defparam i52867_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53403_4_lut (.I0(n24_adj_5261), .I1(n14_adj_5191), .I2(n27_adj_5009), 
            .I3(n66878), .O(n69129));   // verilog/uart_rx.v(119[33:55])
    defparam i53403_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n68593), .I1(baudrate[4]), 
            .I2(n58834), .I3(GND_net), .O(n48_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53404_3_lut (.I0(n69129), .I1(baudrate[10]), .I2(n29_adj_5010), 
            .I3(GND_net), .O(n69130));   // verilog/uart_rx.v(119[33:55])
    defparam i53404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5738_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam i5738_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i53291_3_lut (.I0(n69130), .I1(baudrate[11]), .I2(n31_adj_5013), 
            .I3(GND_net), .O(n69017));   // verilog/uart_rx.v(119[33:55])
    defparam i53291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1050 (.I0(n68703), .I1(baudrate[16]), .I2(n2476), 
            .I3(n61354), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1050.LUT_INIT = 16'h7100;
    SB_LUT4 i54361_2_lut_4_lut (.I0(n68703), .I1(baudrate[16]), .I2(n2476), 
            .I3(n63322), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i54361_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i52925_4_lut (.I0(n41_adj_5031), .I1(n39_adj_5026), .I2(n37_adj_5014), 
            .I3(n66862), .O(n68651));
    defparam i52925_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53455_4_lut (.I0(n68718), .I1(n68811), .I2(n43_adj_5181), 
            .I3(n66850), .O(n69181));   // verilog/uart_rx.v(119[33:55])
    defparam i53455_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7137_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n20844));   // verilog/uart_rx.v(119[33:55])
    defparam i7137_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i53245_3_lut (.I0(n69017), .I1(baudrate[12]), .I2(n33_adj_5036), 
            .I3(GND_net), .O(n68971));   // verilog/uart_rx.v(119[33:55])
    defparam i53245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53532_4_lut (.I0(n68971), .I1(n69181), .I2(n43_adj_5181), 
            .I3(n68651), .O(n69258));   // verilog/uart_rx.v(119[33:55])
    defparam i53532_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53533_3_lut (.I0(n69258), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n69259));   // verilog/uart_rx.v(119[33:55])
    defparam i53533_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5746_2_lut (.I0(n20844), .I1(n11422), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam i5746_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut_adj_1051 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n61318));
    defparam i1_3_lut_4_lut_adj_1051.LUT_INIT = 16'hfffe;
    SB_LUT4 i47852_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n63569));
    defparam i47852_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8315[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5141), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5140), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8003[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8341[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8029[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8055[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8081[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8107[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8133[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8159[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8185[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8211[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8237[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8263[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8289[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43392_1_lut (.I0(n25645), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59070));
    defparam i43392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1052 (.I0(baudrate[17]), .I1(n63523), .I2(baudrate[2]), 
            .I3(n42418), .O(n61282));
    defparam i1_4_lut_adj_1052.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1053 (.I0(n63575), .I1(n61282), .I2(n25639), 
            .I3(n63475), .O(n60615));
    defparam i1_4_lut_adj_1053.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1054 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n42420), .O(n61608));
    defparam i1_4_lut_adj_1054.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1055 (.I0(n61608), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n61626));
    defparam i1_4_lut_adj_1055.LUT_INIT = 16'h0002;
    SB_LUT4 i47914_4_lut (.I0(n63569), .I1(n63475), .I2(n63483), .I3(n63298), 
            .O(n63631));
    defparam i47914_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n63617), .I1(n63631), .I2(n58877), 
            .I3(n61626), .O(n59605));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1057 (.I0(n61846), .I1(n61842), .I2(n61844), 
            .I3(n63298), .O(n61864));
    defparam i1_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(n63523), .I1(n61850), .I2(n61852), 
            .I3(n61848), .O(n61866));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1059 (.I0(n61866), .I1(n25642), .I2(n61864), 
            .I3(GND_net), .O(n25593));
    defparam i1_3_lut_adj_1059.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n59605), .I1(baudrate[2]), 
            .I2(n60615), .I3(GND_net), .O(n48_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i47613_2_lut (.I0(baudrate[17]), .I1(n25639), .I2(GND_net), 
            .I3(GND_net), .O(n63322));
    defparam i47613_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i54369_2_lut (.I0(n48_adj_5170), .I1(n25593), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i54369_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i47840_2_lut_4_lut (.I0(baudrate[6]), .I1(baudrate[7]), .I2(baudrate[8]), 
            .I3(baudrate[9]), .O(n63557));
    defparam i47840_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n61984));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (GND_net, n29837, \data[15] , n29836, \data[12] , n29835, 
            \data[11] , n29834, \data[10] , n29833, \data[9] , n29832, 
            \data[8] , n29831, \data[7] , n29830, \data[6] , n29829, 
            \data[5] , n29828, \data[4] , n29827, \data[3] , n29826, 
            \data[2] , n29825, \data[1] , clk16MHz, VCC_net, CS_c, 
            CS_CLK_c, n29625, \current[0] , n30445, \data[0] , n30365, 
            \current[1] , n30364, \current[2] , n30363, \current[3] , 
            n30362, \current[4] , n30361, \current[5] , n30360, \current[6] , 
            n30359, \current[7] , n30358, \current[8] , n30357, \current[9] , 
            n30356, \current[10] , n30355, \current[11] , n6, n6_adj_4, 
            n5, n5_adj_5, n6_adj_6, state_7__N_4320, n42331, n27704, 
            \current[15] , n25555, n25573, n25579, n25563, n25544, 
            n11) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input n29837;
    output \data[15] ;
    input n29836;
    output \data[12] ;
    input n29835;
    output \data[11] ;
    input n29834;
    output \data[10] ;
    input n29833;
    output \data[9] ;
    input n29832;
    output \data[8] ;
    input n29831;
    output \data[7] ;
    input n29830;
    output \data[6] ;
    input n29829;
    output \data[5] ;
    input n29828;
    output \data[4] ;
    input n29827;
    output \data[3] ;
    input n29826;
    output \data[2] ;
    input n29825;
    output \data[1] ;
    input clk16MHz;
    input VCC_net;
    output CS_c;
    output CS_CLK_c;
    input n29625;
    output \current[0] ;
    input n30445;
    output \data[0] ;
    input n30365;
    output \current[1] ;
    input n30364;
    output \current[2] ;
    input n30363;
    output \current[3] ;
    input n30362;
    output \current[4] ;
    input n30361;
    output \current[5] ;
    input n30360;
    output \current[6] ;
    input n30359;
    output \current[7] ;
    input n30358;
    output \current[8] ;
    input n30357;
    output \current[9] ;
    input n30356;
    output \current[10] ;
    input n30355;
    output \current[11] ;
    output n6;
    output n6_adj_4;
    output n5;
    output n5_adj_5;
    output n6_adj_6;
    output state_7__N_4320;
    output n42331;
    output n27704;
    output \current[15] ;
    output n25555;
    output n25573;
    output n25579;
    output n25563;
    output n25544;
    output n11;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n51686;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n51687;
    wire [11:0]n53;
    
    wire n51685, n51684, n51683, clk_slow_N_4233, n51682, n51681, 
        n51680, n51679, n51678, n51677;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n2;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4234;
    wire [1:0]n1859;
    wire [7:0]n37;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n51583, clk_out, n51582, n51581, n51580, n66358, n51579, 
        n66357, n51578, n66353, n51577, n66362, n9, n29627, n12142, 
        n27868, n28812, n22540, n27761, delay_counter_15__N_4315;
    wire [2:0]n17;
    
    wire n29083, n22542, n22544, n22546, n42874, n51689, n51688, 
        n15, n8, n12, n10, n6_adj_4992;
    
    SB_CARRY delay_counter_1947_1948_add_4_12 (.CI(n51686), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n51687));
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29837));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29836));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29835));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29834));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29833));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29832));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29831));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29830));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29829));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29828));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29827));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29826));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29825));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 delay_counter_1947_1948_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n51685), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_11 (.CI(n51685), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n51686));
    SB_LUT4 delay_counter_1947_1948_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n51684), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_10 (.CI(n51684), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n51685));
    SB_LUT4 delay_counter_1947_1948_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n51683), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4233));   // verilog/tli4970.v(13[10] 19[6])
    SB_CARRY delay_counter_1947_1948_add_4_9 (.CI(n51683), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n51684));
    SB_LUT4 delay_counter_1947_1948_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n51682), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_8 (.CI(n51682), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n51683));
    SB_LUT4 delay_counter_1947_1948_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n51681), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_7 (.CI(n51681), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n51682));
    SB_LUT4 delay_counter_1947_1948_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n51680), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_6 (.CI(n51680), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n51681));
    SB_LUT4 delay_counter_1947_1948_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n51679), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_5 (.CI(n51679), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n51680));
    SB_LUT4 delay_counter_1947_1948_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n51678), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_4 (.CI(n51678), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n51679));
    SB_LUT4 delay_counter_1947_1948_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n51677), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_3 (.CI(n51677), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n51678));
    SB_LUT4 delay_counter_1947_1948_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1947_1948_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n51677));
    SB_LUT4 i2394_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));
    defparam i2394_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2064_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4234));
    defparam i2064_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4234), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4233));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2120_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1859[0]));
    defparam i2120_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_counter_1941_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n51583), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 bit_counter_1941_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n51582), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1941_add_4_8 (.CI(n51582), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n51583));
    SB_LUT4 bit_counter_1941_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n51581), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1941_add_4_7 (.CI(n51581), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n51582));
    SB_LUT4 bit_counter_1941_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n51580), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1941_add_4_6 (.CI(n51580), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n51581));
    SB_LUT4 bit_counter_1941_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n51579), .O(n66358)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1941_add_4_5 (.CI(n51579), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n51580));
    SB_LUT4 bit_counter_1941_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n51578), .O(n66357)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1941_add_4_4 (.CI(n51578), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n51579));
    SB_LUT4 bit_counter_1941_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n51577), .O(n66353)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1941_add_4_3 (.CI(n51577), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n51578));
    SB_LUT4 bit_counter_1941_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n66362)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1941_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1941_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n51577));
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29627));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29625));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n27868), .D(n12142), 
            .R(n28812));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1941__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27761), 
            .D(n22540));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1947_1948__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1949_1950__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4234));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1949_1950__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4234));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1949_1950__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4234));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_1947_1948__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1947_1948__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4315));   // verilog/tli4970.v(40[24:39])
    SB_DFFNESR bit_counter_1941__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27761), 
            .D(n37[4]), .R(n29083));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1941__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27761), 
            .D(n37[5]), .R(n29083));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1941__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27761), 
            .D(n37[6]), .R(n29083));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1941__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27761), 
            .D(n37[7]), .R(n29083));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1941__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27761), 
            .D(n22542));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1941__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27761), 
            .D(n22544));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1941__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27761), 
            .D(n22546));   // verilog/tli4970.v(55[24:39])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30445));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30365));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30364));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30363));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30362));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30361));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30360));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30359));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30358));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30357));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30356));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30355));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_336_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_336_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_334_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4));   // verilog/tli4970.v(54[9:26])
    defparam equal_334_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_334_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_334_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_325_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5));   // verilog/tli4970.v(54[9:26])
    defparam equal_325_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_329_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_6));   // verilog/tli4970.v(54[9:26])
    defparam equal_329_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4320));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28409_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n42331));
    defparam i28409_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27704), 
            .D(n1859[0]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n27868), .D(n42874), 
            .S(n28812));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 counter_1949_1950_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n51689), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1949_1950_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1949_1950_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n51688), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1949_1950_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1949_1950_add_4_3 (.CI(n51688), .I0(GND_net), .I1(counter[1]), 
            .CO(n51689));
    SB_LUT4 counter_1949_1950_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1949_1950_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1949_1950_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n51688));
    SB_LUT4 delay_counter_1947_1948_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n51687), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1947_1948_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n51686), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1947_1948_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(delay_counter_15__N_4315), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n27868));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i14781_2_lut_4_lut (.I0(delay_counter_15__N_4315), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n28812));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14781_2_lut_4_lut.LUT_INIT = 16'h2202;
    SB_LUT4 i15052_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29083));   // verilog/tli4970.v(55[24:39])
    defparam i15052_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8785_3_lut (.I0(state[0]), .I1(n66353), .I2(state[1]), .I3(GND_net), 
            .O(n22546));   // verilog/tli4970.v(55[24:39])
    defparam i8785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8783_3_lut (.I0(state[0]), .I1(n66357), .I2(state[1]), .I3(GND_net), 
            .O(n22544));   // verilog/tli4970.v(55[24:39])
    defparam i8783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8781_3_lut (.I0(state[0]), .I1(n66358), .I2(state[1]), .I3(GND_net), 
            .O(n22542));   // verilog/tli4970.v(55[24:39])
    defparam i8781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(state[0]), 
            .I3(state[1]), .O(n25555));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_4_lut_adj_964 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25573));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_964.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_965 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25579));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_965.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_966 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25563));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_966.LUT_INIT = 16'hfffb;
    SB_LUT4 i54375_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9));
    defparam i54375_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i15596_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n29627));
    defparam i15596_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(state[0]), .I3(state[1]), .O(n25544));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_265_i11_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_265_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13927_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27761));
    defparam i13927_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8779_3_lut (.I0(state[0]), .I1(n66362), .I2(state[1]), .I3(GND_net), 
            .O(n22540));   // verilog/tli4970.v(55[24:39])
    defparam i8779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53624_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n42874));
    defparam i53624_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2065_4_lut (.I0(delay_counter[0]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[3]), .O(n12));
    defparam i2065_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(delay_counter[11]), .I1(delay_counter[7]), .I2(delay_counter[8]), 
            .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4315));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_2032_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n12142));
    defparam mux_2032_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i53613_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n27704));
    defparam i53613_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4992));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_967 (.I0(n11), .I1(bit_counter[7]), .I2(bit_counter[6]), 
            .I3(n6_adj_4992), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut_adj_967.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (\a_new[1] , \b_new[1] , debounce_cnt_N_3834, 
            a_prev, b_prev, position_31__N_3837, GND_net, ENCODER0_B_N_keep, 
            n1779, ENCODER0_A_N_keep, n29707, n1742, n29706, n29672, 
            n1744, \encoder0_position[30] , \encoder0_position[29] , \encoder0_position[28] , 
            \encoder0_position[27] , \encoder0_position[26] , \encoder0_position[25] , 
            \encoder0_position[24] , \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    output \b_new[1] ;
    output debounce_cnt_N_3834;
    output a_prev;
    output b_prev;
    output position_31__N_3837;
    input GND_net;
    input ENCODER0_B_N_keep;
    input n1779;
    input ENCODER0_A_N_keep;
    input n29707;
    output n1742;
    input n29706;
    input n29672;
    output n1744;
    output \encoder0_position[30] ;
    output \encoder0_position[29] ;
    output \encoder0_position[28] ;
    output \encoder0_position[27] ;
    output \encoder0_position[26] ;
    output \encoder0_position[25] ;
    output \encoder0_position[24] ;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire direction_N_3841;
    wire [31:0]n133;
    
    wire n51740, n51739, n51738, n51737, n51736, n51735, n51734, 
        n51733, n51732, n51731, n51730, n51729, n51728, n51727, 
        n51726, n51725, n51724, n51723, n51722, n51721, n51720, 
        n51719, n51718, n51717, n51716, n51715, n51714, n51713, 
        n51712, n51711, n51710;
    
    SB_LUT4 debounce_cnt_I_937_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3834));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_938_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3837));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_938_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3841));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1742), .C(n1779), .D(n29707));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n29706));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29672));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1957_add_4_33_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(n1744), .I3(n51740), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1957_add_4_32_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[30] ), .I3(n51739), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_32 (.CI(n51739), .I0(direction_N_3841), 
            .I1(\encoder0_position[30] ), .CO(n51740));
    SB_LUT4 position_1957_add_4_31_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[29] ), .I3(n51738), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_31 (.CI(n51738), .I0(direction_N_3841), 
            .I1(\encoder0_position[29] ), .CO(n51739));
    SB_LUT4 position_1957_add_4_30_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[28] ), .I3(n51737), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_30 (.CI(n51737), .I0(direction_N_3841), 
            .I1(\encoder0_position[28] ), .CO(n51738));
    SB_LUT4 position_1957_add_4_29_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[27] ), .I3(n51736), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_29 (.CI(n51736), .I0(direction_N_3841), 
            .I1(\encoder0_position[27] ), .CO(n51737));
    SB_LUT4 position_1957_add_4_28_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[26] ), .I3(n51735), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1957__i31 (.Q(n1744), .C(n1779), .E(position_31__N_3837), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1957_add_4_28 (.CI(n51735), .I0(direction_N_3841), 
            .I1(\encoder0_position[26] ), .CO(n51736));
    SB_LUT4 position_1957_add_4_27_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[25] ), .I3(n51734), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1957__i30 (.Q(\encoder0_position[30] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i29 (.Q(\encoder0_position[29] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i28 (.Q(\encoder0_position[28] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i27 (.Q(\encoder0_position[27] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i26 (.Q(\encoder0_position[26] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i25 (.Q(\encoder0_position[25] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i24 (.Q(\encoder0_position[24] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i23 (.Q(\encoder0_position[23] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i22 (.Q(\encoder0_position[22] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i21 (.Q(\encoder0_position[21] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i20 (.Q(\encoder0_position[20] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i19 (.Q(\encoder0_position[19] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i18 (.Q(\encoder0_position[18] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i17 (.Q(\encoder0_position[17] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i16 (.Q(\encoder0_position[16] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i15 (.Q(\encoder0_position[15] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i14 (.Q(\encoder0_position[14] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i13 (.Q(\encoder0_position[13] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i12 (.Q(\encoder0_position[12] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i11 (.Q(\encoder0_position[11] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i10 (.Q(\encoder0_position[10] ), .C(n1779), 
            .E(position_31__N_3837), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i9 (.Q(\encoder0_position[9] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i8 (.Q(\encoder0_position[8] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i7 (.Q(\encoder0_position[7] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i6 (.Q(\encoder0_position[6] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i5 (.Q(\encoder0_position[5] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i4 (.Q(\encoder0_position[4] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i3 (.Q(\encoder0_position[3] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i2 (.Q(\encoder0_position[2] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1957__i1 (.Q(\encoder0_position[1] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1957_add_4_27 (.CI(n51734), .I0(direction_N_3841), 
            .I1(\encoder0_position[25] ), .CO(n51735));
    SB_LUT4 position_1957_add_4_26_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[24] ), .I3(n51733), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_26 (.CI(n51733), .I0(direction_N_3841), 
            .I1(\encoder0_position[24] ), .CO(n51734));
    SB_LUT4 position_1957_add_4_25_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[23] ), .I3(n51732), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1957__i0 (.Q(\encoder0_position[0] ), .C(n1779), .E(position_31__N_3837), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1957_add_4_25 (.CI(n51732), .I0(direction_N_3841), 
            .I1(\encoder0_position[23] ), .CO(n51733));
    SB_LUT4 position_1957_add_4_24_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[22] ), .I3(n51731), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_24 (.CI(n51731), .I0(direction_N_3841), 
            .I1(\encoder0_position[22] ), .CO(n51732));
    SB_LUT4 position_1957_add_4_23_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[21] ), .I3(n51730), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_23 (.CI(n51730), .I0(direction_N_3841), 
            .I1(\encoder0_position[21] ), .CO(n51731));
    SB_LUT4 position_1957_add_4_22_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[20] ), .I3(n51729), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_22 (.CI(n51729), .I0(direction_N_3841), 
            .I1(\encoder0_position[20] ), .CO(n51730));
    SB_LUT4 position_1957_add_4_21_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[19] ), .I3(n51728), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_21 (.CI(n51728), .I0(direction_N_3841), 
            .I1(\encoder0_position[19] ), .CO(n51729));
    SB_LUT4 position_1957_add_4_20_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[18] ), .I3(n51727), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_20 (.CI(n51727), .I0(direction_N_3841), 
            .I1(\encoder0_position[18] ), .CO(n51728));
    SB_LUT4 position_1957_add_4_19_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[17] ), .I3(n51726), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_19 (.CI(n51726), .I0(direction_N_3841), 
            .I1(\encoder0_position[17] ), .CO(n51727));
    SB_LUT4 position_1957_add_4_18_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[16] ), .I3(n51725), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_18 (.CI(n51725), .I0(direction_N_3841), 
            .I1(\encoder0_position[16] ), .CO(n51726));
    SB_LUT4 position_1957_add_4_17_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[15] ), .I3(n51724), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_17 (.CI(n51724), .I0(direction_N_3841), 
            .I1(\encoder0_position[15] ), .CO(n51725));
    SB_LUT4 position_1957_add_4_16_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[14] ), .I3(n51723), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_16 (.CI(n51723), .I0(direction_N_3841), 
            .I1(\encoder0_position[14] ), .CO(n51724));
    SB_LUT4 position_1957_add_4_15_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[13] ), .I3(n51722), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_15 (.CI(n51722), .I0(direction_N_3841), 
            .I1(\encoder0_position[13] ), .CO(n51723));
    SB_LUT4 position_1957_add_4_14_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[12] ), .I3(n51721), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_14 (.CI(n51721), .I0(direction_N_3841), 
            .I1(\encoder0_position[12] ), .CO(n51722));
    SB_LUT4 position_1957_add_4_13_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[11] ), .I3(n51720), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_13 (.CI(n51720), .I0(direction_N_3841), 
            .I1(\encoder0_position[11] ), .CO(n51721));
    SB_LUT4 position_1957_add_4_12_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[10] ), .I3(n51719), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_12 (.CI(n51719), .I0(direction_N_3841), 
            .I1(\encoder0_position[10] ), .CO(n51720));
    SB_LUT4 position_1957_add_4_11_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[9] ), .I3(n51718), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_11 (.CI(n51718), .I0(direction_N_3841), 
            .I1(\encoder0_position[9] ), .CO(n51719));
    SB_LUT4 position_1957_add_4_10_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[8] ), .I3(n51717), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_10 (.CI(n51717), .I0(direction_N_3841), 
            .I1(\encoder0_position[8] ), .CO(n51718));
    SB_LUT4 position_1957_add_4_9_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[7] ), .I3(n51716), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_9 (.CI(n51716), .I0(direction_N_3841), 
            .I1(\encoder0_position[7] ), .CO(n51717));
    SB_LUT4 position_1957_add_4_8_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[6] ), .I3(n51715), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_8 (.CI(n51715), .I0(direction_N_3841), 
            .I1(\encoder0_position[6] ), .CO(n51716));
    SB_LUT4 position_1957_add_4_7_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[5] ), .I3(n51714), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_7 (.CI(n51714), .I0(direction_N_3841), 
            .I1(\encoder0_position[5] ), .CO(n51715));
    SB_LUT4 position_1957_add_4_6_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[4] ), .I3(n51713), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_6 (.CI(n51713), .I0(direction_N_3841), 
            .I1(\encoder0_position[4] ), .CO(n51714));
    SB_LUT4 position_1957_add_4_5_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[3] ), .I3(n51712), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_5 (.CI(n51712), .I0(direction_N_3841), 
            .I1(\encoder0_position[3] ), .CO(n51713));
    SB_LUT4 position_1957_add_4_4_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[2] ), .I3(n51711), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_1957_add_4_4 (.CI(n51711), .I0(direction_N_3841), 
            .I1(\encoder0_position[2] ), .CO(n51712));
    SB_LUT4 position_1957_add_4_3_lut (.I0(GND_net), .I1(direction_N_3841), 
            .I2(\encoder0_position[1] ), .I3(n51710), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_3 (.CI(n51710), .I0(direction_N_3841), 
            .I1(\encoder0_position[1] ), .CO(n51711));
    SB_LUT4 position_1957_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1957_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1957_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n51710));
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (GND_net, n2874, pwm_out, clk32MHz, reset, VCC_net, pwm_setpoint) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n2874;
    output pwm_out;
    input clk32MHz;
    input reset;
    input VCC_net;
    input [23:0]pwm_setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n59859, n14, n13, n8, n10, n48, pwm_out_N_577, n56571, 
        n51576, n56599, n51575, n56619, n51574, n56647, n51573, 
        n57493, n56675, n51572, n56703, n51571, n56737, n51570, 
        n56779, n56821, n56859, n56893, n56917, n56943, n56975, 
        n57001, n57031, n57061, n57097, n57151, n57359, n57497, 
        n57499, n57501, n51569, n51568, n51567, n51566, n51565, 
        n51564, n51563, n51562, n51561, n51560, n51559, n51558, 
        n51557, n51556, n51555, n51554, n8_adj_4986, n66779, n16, 
        n10_adj_4987, n66815, n12, n41, n39, n45, n43, n37, 
        n29, n31, n23, n25, n35, n11, n13_adj_4988, n27, n15, 
        n33, n9, n17, n19, n21, n66873, n66842, n30, n66936, 
        n67804, n67796, n68933, n68335, n69098, n6, n68359, n68360, 
        n24, n66783, n68279, n67571, n4, n68357, n68358, n66826, 
        n68939, n67573, n69179, n69180, n69107, n66798, n68883, 
        n67579, n69084;
    
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n59859));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[16]), .I1(pwm_counter[14]), .I2(pwm_counter[19]), 
            .I3(pwm_counter[17]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(pwm_counter[11]), .I1(pwm_counter[18]), .I2(pwm_counter[22]), 
            .I3(pwm_counter[15]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n59859), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n8));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut (.I0(pwm_counter[21]), .I1(n8), .I2(n13), .I3(n14), 
            .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[13]), .I2(n10), 
            .I3(pwm_counter[20]), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2874), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_1940_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n51576), .O(n56571)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1940_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n51575), .O(n56599)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_24 (.CI(n51575), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n51576));
    SB_LUT4 pwm_counter_1940_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n51574), .O(n56619)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_23 (.CI(n51574), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n51575));
    SB_LUT4 pwm_counter_1940_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n51573), .O(n56647)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_DFFR pwm_counter_1940__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n57493), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_1940_add_4_22 (.CI(n51573), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n51574));
    SB_LUT4 pwm_counter_1940_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n51572), .O(n56675)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_21 (.CI(n51572), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n51573));
    SB_LUT4 pwm_counter_1940_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n51571), .O(n56703)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_20 (.CI(n51571), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n51572));
    SB_LUT4 pwm_counter_1940_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n51570), .O(n56737)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_DFFR pwm_counter_1940__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n56571), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n56599), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n56619), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n56647), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n56675), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n56703), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n56737), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n56779), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n56821), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n56859), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n56893), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n56917), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n56943), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n56975), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n57001), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n57031), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n57061), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n57097), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n57151), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n57359), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n57497), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n57499), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1940__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n57501), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_1940_add_4_19 (.CI(n51570), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n51571));
    SB_LUT4 pwm_counter_1940_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n51569), .O(n56779)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_18 (.CI(n51569), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n51570));
    SB_LUT4 pwm_counter_1940_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n51568), .O(n56821)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_17 (.CI(n51568), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n51569));
    SB_LUT4 pwm_counter_1940_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n51567), .O(n56859)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_16 (.CI(n51567), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n51568));
    SB_LUT4 pwm_counter_1940_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n51566), .O(n56893)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_15 (.CI(n51566), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n51567));
    SB_LUT4 pwm_counter_1940_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n51565), .O(n56917)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_14 (.CI(n51565), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n51566));
    SB_LUT4 pwm_counter_1940_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n51564), .O(n56943)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_13 (.CI(n51564), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n51565));
    SB_LUT4 pwm_counter_1940_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n51563), .O(n56975)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_12 (.CI(n51563), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n51564));
    SB_LUT4 pwm_counter_1940_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n51562), .O(n57001)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_11 (.CI(n51562), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n51563));
    SB_LUT4 pwm_counter_1940_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n51561), .O(n57031)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_10 (.CI(n51561), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n51562));
    SB_LUT4 pwm_counter_1940_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n51560), .O(n57061)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_9 (.CI(n51560), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n51561));
    SB_LUT4 pwm_counter_1940_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n51559), .O(n57097)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_8 (.CI(n51559), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n51560));
    SB_LUT4 pwm_counter_1940_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n51558), .O(n57151)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_7 (.CI(n51558), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n51559));
    SB_LUT4 pwm_counter_1940_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n51557), .O(n57359)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_6 (.CI(n51557), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n51558));
    SB_LUT4 pwm_counter_1940_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n51556), .O(n57497)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_5 (.CI(n51556), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n51557));
    SB_LUT4 pwm_counter_1940_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n51555), .O(n57499)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_4 (.CI(n51555), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n51556));
    SB_LUT4 pwm_counter_1940_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n51554), .O(n57501)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_3 (.CI(n51554), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n51555));
    SB_LUT4 pwm_counter_1940_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n57493)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1940_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1940_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n51554));
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4986));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51053_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n66779));
    defparam i51053_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4987));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51089_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n66815));
    defparam i51089_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4988));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51147_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n66873));
    defparam i51147_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51116_4_lut (.I0(n27), .I1(n15), .I2(n13_adj_4988), .I3(n11), 
            .O(n66842));
    defparam i51116_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52078_4_lut (.I0(n13_adj_4988), .I1(n11), .I2(n9), .I3(n66936), 
            .O(n67804));
    defparam i52078_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52070_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n67804), 
            .O(n67796));
    defparam i52070_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53207_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n67796), 
            .O(n68933));
    defparam i53207_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52609_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n68933), 
            .O(n68335));
    defparam i52609_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53372_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n68335), 
            .O(n69098));
    defparam i53372_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52633_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n68359));   // verilog/pwm.v(21[8:24])
    defparam i52633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52634_3_lut (.I0(n68359), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n68360));   // verilog/pwm.v(21[8:24])
    defparam i52634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51057_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n66873), 
            .O(n66783));
    defparam i51057_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52553_4_lut (.I0(n24), .I1(n8_adj_4986), .I2(n45), .I3(n66779), 
            .O(n68279));   // verilog/pwm.v(21[8:24])
    defparam i52553_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51845_3_lut (.I0(n68360), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n67571));   // verilog/pwm.v(21[8:24])
    defparam i51845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52631_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n68357));   // verilog/pwm.v(21[8:24])
    defparam i52631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52632_3_lut (.I0(n68357), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n68358));   // verilog/pwm.v(21[8:24])
    defparam i52632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51100_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n66842), 
            .O(n66826));
    defparam i51100_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53213_4_lut (.I0(n30), .I1(n10_adj_4987), .I2(n35), .I3(n66815), 
            .O(n68939));   // verilog/pwm.v(21[8:24])
    defparam i53213_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51847_3_lut (.I0(n68358), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n67573));   // verilog/pwm.v(21[8:24])
    defparam i51847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53453_4_lut (.I0(n67573), .I1(n68939), .I2(n35), .I3(n66826), 
            .O(n69179));   // verilog/pwm.v(21[8:24])
    defparam i53453_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53454_3_lut (.I0(n69179), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n69180));   // verilog/pwm.v(21[8:24])
    defparam i53454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53381_3_lut (.I0(n69180), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n69107));   // verilog/pwm.v(21[8:24])
    defparam i53381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51072_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n69098), 
            .O(n66798));
    defparam i51072_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53157_4_lut (.I0(n67571), .I1(n68279), .I2(n45), .I3(n66783), 
            .O(n68883));   // verilog/pwm.v(21[8:24])
    defparam i53157_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51853_3_lut (.I0(n69107), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n67579));   // verilog/pwm.v(21[8:24])
    defparam i51853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53358_4_lut (.I0(n67579), .I1(n68883), .I2(n45), .I3(n66798), 
            .O(n69084));   // verilog/pwm.v(21[8:24])
    defparam i53358_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53359_3_lut (.I0(n69084), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i53359_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51210_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n66936));   // verilog/pwm.v(21[8:24])
    defparam i51210_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, n182, IntegralLimit, n156, \Kp[1] , 
            \Kp[0] , \Kp[2] , \Ki[7] , \Kp[3] , \Kp[4] , \Kp[5] , 
            \Ki[8] , \Kp[6] , \Kp[7] , \Ki[9] , \Ki[1] , \Kp[8] , 
            \Kp[9] , \Kp[10] , \Ki[2] , \Ki[3] , n150, \Ki[0] , 
            \Ki[4] , \Ki[5] , n6, n37154, n20194, \Kp[13] , n20185, 
            n214, \Ki[6] , \Kp[14] , clk16MHz, duty, reset, n37050, 
            n4, \Kp[11] , \Kp[12] , PWMLimit, n406, setpoint, n15, 
            n405, \Kp[15] , n478, n135, n500, \Ki[10] , VCC_net, 
            n187, \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , 
            n41, deadband, \motor_state[23] , \motor_state[22] , n219, 
            \motor_state[21] , \motor_state[20] , \motor_state[19] , \motor_state[18] , 
            \motor_state[17] , n20112, n20113, n7, n56, \motor_state[15] , 
            \motor_state[14] , \motor_state[13] , \motor_state[12] , \motor_state[11] , 
            \motor_state[10] , \motor_state[9] , n10, \motor_state[7] , 
            \motor_state[6] , \motor_state[5] , \motor_state[4] , \motor_state[3] , 
            \motor_state[2] , \motor_state[1] , n18, \duty_23__N_3602[7] , 
            \duty_23__N_3602[4] , n624, n551, n478_adj_1, n405_adj_2, 
            n332, n259, n186, n113, n244, n36515, n41_adj_3, \data_in_frame[9][7] , 
            \data_in_frame[6][3] , \data_in_frame[8][4] , \data_in_frame[8][2] , 
            n58520, \data_in_frame[4][2] , \data_in_frame[8][6] , \data_in_frame[1][6] , 
            \data_in_frame[12][0] , n58075, n58405, n58556, \data_in_frame[3][7] , 
            \data_in_frame[4][1] , \data_in_frame[8][3] , n58766, n50204, 
            n50001, n62, n20158, n20159, n42880) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n182;
    input [23:0]IntegralLimit;
    output n156;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Ki[7] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Ki[8] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Ki[9] ;
    input \Ki[1] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Ki[2] ;
    input \Ki[3] ;
    output n150;
    input \Ki[0] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input n6;
    input n37154;
    output n20194;
    input \Kp[13] ;
    input n20185;
    output n214;
    input \Ki[6] ;
    input \Kp[14] ;
    input clk16MHz;
    output [23:0]duty;
    input reset;
    input n37050;
    input n4;
    input \Kp[11] ;
    input \Kp[12] ;
    input [23:0]PWMLimit;
    output n406;
    input [23:0]setpoint;
    input n15;
    output n405;
    input \Kp[15] ;
    output n478;
    output n135;
    output n500;
    input \Ki[10] ;
    input VCC_net;
    output n187;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input n41;
    input [23:0]deadband;
    input \motor_state[23] ;
    input \motor_state[22] ;
    output n219;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input n20112;
    input n20113;
    input n7;
    input n56;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input n10;
    input \motor_state[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input n18;
    input \duty_23__N_3602[7] ;
    input \duty_23__N_3602[4] ;
    input n624;
    input n551;
    input n478_adj_1;
    input n405_adj_2;
    input n332;
    input n259;
    input n186;
    input n113;
    input n244;
    input n36515;
    input n41_adj_3;
    input \data_in_frame[9][7] ;
    input \data_in_frame[6][3] ;
    input \data_in_frame[8][4] ;
    input \data_in_frame[8][2] ;
    input n58520;
    input \data_in_frame[4][2] ;
    input \data_in_frame[8][6] ;
    input \data_in_frame[1][6] ;
    input \data_in_frame[12][0] ;
    input n58075;
    input n58405;
    input n58556;
    input \data_in_frame[3][7] ;
    input \data_in_frame[4][1] ;
    input \data_in_frame[8][3] ;
    output n58766;
    output n50204;
    output n50001;
    input n62;
    output n20158;
    output n20159;
    output n42880;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n50826;
    wire [15:0]n16950;
    
    wire n603, n50827, n50500;
    wire [23:0]n46;
    
    wire n50501, n51808;
    wire [11:0]n18947;
    
    wire n834, n51809;
    wire [21:0]n12695;
    wire [20:0]n13661;
    
    wire n51986;
    wire [23:0]n379;
    
    wire n50499;
    wire [16:0]n16339;
    
    wire n530, n50825, n50388;
    wire [43:0]n258;
    wire [47:0]n303;
    
    wire n50389;
    wire [23:0]n353;
    
    wire n50387, n50498, n51987, n51985, n51984;
    wire [23:0]n48;
    wire [23:0]n49;
    wire [23:0]n208;
    wire [23:0]n233;
    wire [23:0]n105;
    
    wire n113_c, n44, n186_c, n554, n259_c, n332_c, n405_c, n627, 
        n478_c, n551_c, n700, n83, n14, n51983, n156_adj_4431, 
        n229, n302, n375_adj_4432, n125, n624_c, n697, n770, n51982, 
        n198, n448;
    wire [12:0]n18613;
    
    wire n761, n51807, n271, n521, n86, n17, n344, n688, n51806, 
        n594, n159, n417;
    wire [3:0]n20155;
    wire [4:0]n20109;
    
    wire n51981, n204, n1099, n51980, n615, n51805, n542, n51804, 
        n314, n131, n1026, n51979, n451, n953, n51978, n950, 
        n387, n4_adj_4434, n524, n457, n50824, n597, n460, n1023, 
        n469, n51803, n880, n51977, n807, n51976, n734, n51975, 
        n396, n51802, n661, n51974, n588, n51973, n384, n50823, 
        counter_31__N_3714, control_update;
    wire [23:0]duty_23__N_3602;
    
    wire n27916, n490, n323, n51801, n250_adj_4436, n51800, n62866, 
        n311, n50822, n62868, n177, n51799, n515, n51972, n442, 
        n51971, n35, n104, n50153, n62856, n533, n369, n51970, 
        n8, n6_adj_4437, n62874, n60827, n238_adj_4439, n50821, 
        n50386;
    wire [6:0]n19869;
    wire [5:0]n19980;
    
    wire n560, n51798, n296, n51969, n165, n50820, n232, n487, 
        n51797, n23, n92, n606, n50497, n670, n679, n667, n101, 
        n50496, n414, n51796, n32, n223, n51968, n305, n174, 
        n50495, n740, n247, n150_adj_4444, n51967, n341, n51795, 
        n378;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n50385, n813, n320, n50494, n50384, n886, n50493, n393, 
        n8_adj_4446, n77, n451_adj_4447, n466, n539, n959;
    wire [19:0]n14539;
    
    wire n51966, n612, n1032, n685;
    wire [23:0]n433;
    
    wire n432;
    wire [23:0]n458;
    wire [23:0]n483;
    
    wire n1, n3_adj_4449, n1105, n268, n51794, n50492, n50491, 
        n50383, n51965, n50490, n758, n50382, n50489, n50488, 
        n195, n51793, n524_adj_4454, n50381, n50487, n50380, n50486, 
        n50379, n50485, n597_adj_4458, n50378, n831, n53, n122_adj_4459;
    wire [14:0]n17493;
    
    wire n50801, n50484, n1117, n50800;
    wire [10:0]n19231;
    
    wire n910, n51792, n50483, n1044, n50799, n971, n50798;
    wire [23:0]n51;
    
    wire n837, n51791, n51964, n51963, n898, n50797, n825, n50796, 
        n904, n752, n50795, n977, n1050, n679_adj_4462, n50794;
    wire [20:0]n13134;
    wire [19:0]n14058;
    
    wire n51006, n50377, n51005, n50482, n764, n51790, n606_adj_4463, 
        n50793, n691, n51789, n618, n51788, n51962, n51961, n51004, 
        n533_adj_4464, n50792, n1102, n51960, n51003, n50376, n460_adj_4465, 
        n50791, n1029, n51959, n51002, n50481, n387_adj_4466, n50790, 
        n50375, n314_adj_4467, n50789, n50480, n545, n51787, n50374, 
        n241, n50788, n50479, n472_adj_4470, n51786, n956, n51958, 
        n883, n51957, n168, n50787, n670_adj_4471, n810, n51956, 
        n743, n399_adj_4473, n51785, n66320, n42898, n326, n51784, 
        n51001, n26, n95, n1102_adj_4477, n51000, n737, n51955;
    wire [6:0]n19947;
    wire [5:0]n20041;
    
    wire n560_adj_4478, n50786, n1029_adj_4479, n50999, n487_adj_4480, 
        n50785, n956_adj_4481, n50998, n50373, n414_adj_4482, n50784, 
        n50478, n253_adj_4483, n51783, n341_adj_4485, n50783, n664, 
        n51954, n50477, n180, n51782, n268_adj_4487, n50782, n50372, 
        n883_adj_4488, n50997, n50476, n810_adj_4490, n50996, n195_adj_4491, 
        n50781, n591, n51953, n737_adj_4492, n50995, n53_adj_4493, 
        n122_adj_4494, n50475, n50371, n518, n51952, n50474, n38, 
        n107_adj_4497, n50370, n664_adj_4498, n50994, n50473;
    wire [9:0]n19469;
    
    wire n840, n51781, n445_adj_4500, n51951, n767, n51780, n591_adj_4501, 
        n50993, n50472, n1_adj_4503, n518_adj_4504, n50992, n372_adj_4505, 
        n51950, n445_adj_4506, n50991, n50369, n299_adj_4507, n51949, 
        n372_adj_4508, n50990, n3_adj_4509, n299_adj_4510, n50989, 
        n226_adj_4511, n50988, n816, n1_adj_4512, n3_adj_4513, n50471, 
        n50470, n153, n50987, n50469;
    wire [11:0]n18754;
    wire [10:0]n19065;
    
    wire n910_adj_4517, n50593, n837_adj_4518, n50592, n764_adj_4519, 
        n50591, n694, n51779, n60191, n490_adj_4521, n51312, n11_adj_4522, 
        n80, n226_adj_4523, n51948;
    wire [4:0]n20063;
    
    wire n417_adj_4524, n51311, n153_adj_4525, n51947, n621, n51778, 
        n11_adj_4526, n80_adj_4527, n691_adj_4528, n50590, n618_adj_4529, 
        n50589, n50368, n50468;
    wire [18:0]n15335;
    
    wire n51946, n548, n51777, n344_adj_4532, n51310, n743_adj_4533;
    wire [13:0]n17972;
    
    wire n1120, n50763, n1047, n50762, n51945, n475_adj_4534, n51776, 
        n402_adj_4535, n51775, n271_adj_4537, n51309, n50367, n889, 
        n329, n51774, n50467, n198_adj_4540, n51308, n51944, n256_adj_4541, 
        n51773, n51943, n974, n50761, n545_adj_4542, n50588, n472_adj_4543, 
        n50587, n56_c, n125_adj_4544, n901, n50760, n828, n50759, 
        n399_adj_4545, n50586, n50366, n755, n50758, n51942, n326_adj_4546, 
        n50585, n1105_adj_4547, n51941, n752_adj_4548, n825_adj_4549, 
        n1096, n816_adj_4550, n962, n1035, n1032_adj_4552, n51940, 
        n682, n50757, n889_adj_4553, n609, n50756, n962_adj_4554, 
        n1035_adj_4555, n183, n51772, n536, n50755, n959_adj_4556, 
        n51939, n463, n50754, n1108, n886_adj_4557, n51938, n813_adj_4558, 
        n51937, n253_adj_4559, n50584, n110_adj_4560, n41_adj_4561, 
        n1108_adj_4562, n39, n45, n37, n43, n390_adj_4567, n50753, 
        n21_adj_4568, n317, n50752, n23_adj_4569, n180_adj_4570, n50583, 
        n50466, n244_c, n50751, n171, n50750, n740_adj_4572, n51936, 
        n50465, n38_adj_4574, n107_adj_4575, n50365, n25_adj_4576, 
        n29, n98, n50464, n50463, n29_adj_4580, n31, n17_adj_4581, 
        n667_adj_4582, n51935, n594_adj_4583, n51934, n50364, n19_adj_4586, 
        n9_adj_4587, n35_adj_4588, n11_adj_4589, n898_adj_4590, n521_adj_4591, 
        n51933, n448_adj_4592, n51932, n375_adj_4593, n51931, n13_adj_4594, 
        n15_adj_4595, n27, n33, n67318, n302_adj_4596, n51930, n229_adj_4597, 
        n51929, n68158, n70652, n156_adj_4598, n51928, n14_adj_4599, 
        n83_adj_4600;
    wire [17:0]n16053;
    
    wire n51927, n51926, n68140, n70647, n67308, n971_adj_4601, 
        n68152, n51925, n70667, n68146, n70662, n16_adj_4602, n67281, 
        n8_adj_4603, n24_adj_4604, n67329, n70660, n67326, n70688, 
        n68513, n51924, n50462, n70685, n50461, n50460, n50363, 
        n50459, n50458, n51923, n68156, n68779, n67300, n51922, 
        n70651, n51921, n68507, n70677, n69018, n51920, n50457, 
        n50362, n51919, n70641, n69227, n50361, n50456, n70638;
    wire [18:0]n14897;
    
    wire n50964, n67355, n12_adj_4606, n50963, n51918, n10_adj_4607, 
        n30, n67418, n68195, n68191, n69072, n68523, n69143, n16_adj_4608, 
        n8_adj_4609, n24_adj_4610, n6_adj_4611, n68655, n68656, n67399, 
        n67334, n67332, n68289, n67599, n4_adj_4612, n68645, n68646, 
        n12_adj_4613, n67292, n70673, n10_adj_4614, n30_adj_4615, 
        n67294, n69034, n67611, n69214, n69215, n69172, n6_adj_4616, 
        n68647, n68648, n67283, n70636, n68291, n67609, n67285, 
        n68899, n67617, n50962, n69090, n51917, n4_adj_4617, n68653, 
        n68654, n67345, n67342, n69100, n67601, n69212, n69213, 
        n69176, n67336;
    wire [12:0]n18391;
    
    wire n50733, n50732, n50731, n68897, n67607, n50961, n50730, 
        n51916, n50960, n51915, n50729, n50360, n50959, n47, n69091, 
        n50728, n69088, n50958, n50359, n50727, n50957, n50726, 
        n50725, n51914, n50358, n50724, n50956, n50723, n50955, 
        n51913, n50722, n50954, n50721, n51912, n9_adj_4618, n13_adj_4619, 
        n15_adj_4620, n50953, n50357, n51911, n21_adj_4621, n50720, 
        n50719, n19_adj_4622, n17_adj_4623, n51910, n50952, n50356, 
        n9_adj_4624, n11_adj_4625, n50049, n62910, n13_adj_4626, n50718, 
        n15_adj_4627, n50951, n50717, n50950, n50716, n50355, n21_adj_4629;
    wire [9:0]n19328;
    wire [8:0]n19547;
    
    wire n51909, n19_adj_4630, n51908, n51907, n50949, n50948, n17_adj_4632, 
        n1044_adj_4633, n50354, n50947, n1117_adj_4634;
    wire [3:0]n20122;
    
    wire n4_adj_4635, n50946, n50353, n50352, n29696;
    wire [8:0]n19665;
    wire [7:0]n19823;
    
    wire n50945, n51906, n51905, n50944, n51904, n51903, n51902, 
        n50943, n50351, n29668, n29667, n29665, n51901, n29663;
    wire [16:0]n16697;
    
    wire n51900, n51899, n51898, n29662, n29661, n29660, n481_adj_4637, 
        n50942, n408, n50941, n1111, n51897, n50350, n45_adj_4638, 
        n335, n50940, n50349, n25_adj_4639, n31_adj_4640, n27_adj_4641, 
        n29_adj_4642, n19_adj_4643, n21_adj_4644, n29632, n1038, n51896, 
        n965, n51895, n23_adj_4645, n50348, n15_adj_4646, n17_adj_4647, 
        n262, n50939, n980, n50700, n907, n50699, n189_adj_4648, 
        n50938, n50347, n7_adj_4650, n47_adj_4651, n116_adj_4652, 
        n834_adj_4653, n50698, n9_adj_4654, n892, n51894, n761_adj_4655, 
        n50697, n11_adj_4656, n819, n51893, n13_adj_4657, n746, 
        n51892, n673, n51891, n600, n51890, n5_adj_4658, n67277, 
        n67273, n68773, n4_adj_4659, n68635, n68636, n10_adj_4660, 
        n67275, n68096, n12_adj_4661, n67623, n116_adj_4662, n47_adj_4663, 
        n50346, n8_adj_4664, n527, n51889, n6_adj_4665, n16_adj_4666, 
        n67271, n69038, n69039, n68926, n68098, n68602, n67621, 
        n68604, n34, n454_adj_4667, n51888, n36, n381_adj_4668, 
        n51887, n308, n51886, n38_adj_4669, n235_adj_4670, n51885;
    wire [31:0]n52;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n51645, n688_adj_4672, n50696, n40, n42, n44_adj_4673, 
        n67242, n68605, n41_adj_4674, n27_adj_4675, n25_adj_4676, 
        n23_adj_4677, n162, n51884, n51644, n20_adj_4679, n89, n615_adj_4680, 
        n50695, n21_adj_4681, n4_adj_4683, n15_adj_4684, n17_adj_4685, 
        n19_adj_4686, n9_adj_4687;
    wire [15:0]n17271;
    
    wire n51883, n11_adj_4688, n13_adj_4689, n7_adj_4690, n67236, 
        n67231, n12_adj_4691, n6_adj_4692, n14_adj_4693, n10_adj_4694, 
        n8_adj_4695, n18_adj_4696, n67229, n69040, n69041, n68924, 
        n68769, n67234, n69121, n67627, n69198, n69199, n29619, 
        n51882, n69118, n34_adj_4697, n36_adj_4698, n38_adj_4699, 
        n40_adj_4700, n67216, n69042, n69043, n68920, n8_adj_4701, 
        n12_adj_4702, n1114, n51881, n16_adj_4703, n10_adj_4704, n61067, 
        n8_adj_4705, n60808, n10_adj_4706, n12_adj_4707, n16_adj_4708, 
        n11_adj_4709, n542_adj_4710, n50694, n50345, n469_adj_4711, 
        n50693, n396_adj_4712, n50692, n1041, n51880, n51643, n51642, 
        n968, n51879, n51641, n895, n51878, n822, n51877, n51640, 
        n749, n51876, n676, n51875, n603_adj_4718, n51874, n51639, 
        n323_adj_4738, n50691, n250_adj_4739, n50690, n50344, n530_adj_4740, 
        n51873, n50343, n457_adj_4741, n51872, n177_adj_4742, n50689, 
        n35_adj_4743, n104_adj_4744, n30459, n30458, n30457, n30456, 
        n30450, n30449, n30447, n30446, n30444, n30411, n30410, 
        n30407, n30406, n51638, n50342, n384_adj_4745, n51871, n311_adj_4746, 
        n51870, n51637, n238_adj_4747, n51869, n50341, n30227, n165_adj_4748, 
        n51868, n23_adj_4749, n92_adj_4750;
    wire [7:0]n19726;
    
    wire n700_adj_4751, n51867, n347, n6_adj_4752, n58043, n627_adj_4753, 
        n51866, n62906, n62_c, n51636, n51635, n554_adj_4754, n51865, 
        n481_adj_4755, n51864, n408_adj_4756, n51863, n51634, n335_adj_4757, 
        n51862, n189_adj_4758, n262_adj_4759, n51861, n50063, n50278, 
        n51860, n62896, n70741, n62900, n8_adj_4760;
    wire [0:0]n11613;
    wire [21:0]n12072;
    
    wire n51105, n50340;
    wire [14:0]n17779;
    
    wire n51859, n51633, n6_adj_4761, n51104, n51632, n51631, n51103, 
        n51102, n51101, n51630, n51629, n51628, n51627, n51858, 
        n51857;
    wire [17:0]n15656;
    
    wire n50916, n51856, n50915, n51626, n51855, n51100, n50914, 
        n50913, n51099, n50912, n50911, n51098, n50910, n50909, 
        n51625, n50908, n51097, n51854, n51853, n50907, n51852, 
        n50906, n51851, n51850, n51096, n51849, n50905, n50904, 
        n51848, n51095, n50903, n51624, n51847, n378_adj_4764, n50902, 
        n877, n51094, n305_adj_4765, n50901, n232_adj_4766, n50900, 
        n804, n51093, n159_adj_4767, n50899, n731, n51092, n658, 
        n51091, n17_adj_4768, n86_adj_4769, n585, n51090, n512, 
        n51089, n439_adj_4771, n51088, n241_adj_4772, n51846, n51623, 
        n366_adj_4773, n51087, n168_adj_4774, n51845, n293_adj_4775, 
        n51086, n220_adj_4776, n51085, n26_adj_4777, n95_adj_4778, 
        n147_adj_4779, n51084;
    wire [13:0]n18225;
    
    wire n1120_adj_4780, n51844, n5_adj_4781, n74, n1047_adj_4782, 
        n51843, n50878, n50877, n50876, n77_adj_4783, n1111_adj_4784, 
        n50875, n974_adj_4785, n51842, n1038_adj_4786, n50874, n8_adj_4787, 
        n965_adj_4788, n50873, n51622, n892_adj_4789, n50872, n819_adj_4790, 
        n50871, n746_adj_4791, n50870, n673_adj_4792, n50869, n600_adj_4793, 
        n50868;
    wire [23:0]n54;
    
    wire n50524, n50523, n527_adj_4796, n50867, n901_adj_4797, n51841, 
        n454_adj_4798, n50866, n51621, n381_adj_4799, n50865, n828_adj_4800, 
        n51840, n50522;
    wire [0:0]n12188;
    
    wire n50408, n50407, n50521, n51620, n308_adj_4804, n50864, 
        n755_adj_4805, n51839, n235_adj_4806, n50863, n162_adj_4807, 
        n50862, n20_adj_4808, n89_adj_4809, n50406, n630, n50861, 
        n557, n50860, n484_adj_4810, n50859, n51619, n50405, n50520, 
        n50404, n682_adj_4813, n51838, n411, n50858, n338, n50857, 
        n50519, n265, n50856, n609_adj_4815, n51837, n51618, n50403, 
        n192_adj_4816, n50855, n50, n119_adj_4817, n50402, n50518, 
        n50401, n50517, n50400, n50399, n51617, n50516, n770_adj_4822, 
        n51059, n50515, n697_adj_4824, n51058, n536_adj_4825, n51836, 
        n463_adj_4826, n51835, n390_adj_4827, n51834, n317_adj_4828, 
        n51833, n907_adj_4829, n51616, n244_adj_4830, n51832, n51615, 
        n171_adj_4831, n51831, n29_adj_4832, n98_adj_4833, n980_adj_4834, 
        n51057, n50398, n51056, n676_adj_4838, n749_adj_4839, n51055, 
        n50397, n51054, n50514, n630_adj_4843, n51830, n557_adj_4844, 
        n51829, n484_adj_4845, n51828, n411_adj_4846, n51827, n50396, 
        n51053, n338_adj_4848, n51826, n101_adj_4849, n32_adj_4850, 
        n66612, n265_adj_4851, n51825, n192_adj_4852, n51824, n174_adj_4853, 
        n50_adj_4854, n119_adj_4855, n51052, n150_adj_4857, n247_adj_4858, 
        n74_adj_4859, n1050_adj_4860, n51823, n5_adj_4861, n977_adj_4862, 
        n51822, n6_adj_4863, n51051, n50513, n840_adj_4867, n52019, 
        n767_adj_4868, n52018, n694_adj_4869, n52017, n621_adj_4870, 
        n52016, n548_adj_4871, n52015, n475_adj_4872, n52014, n44_adj_4873, 
        n402_adj_4875, n52013, n147_adj_4876, n329_adj_4877, n52012, 
        n256_adj_4879, n52011, n904_adj_4880, n51821, n183_adj_4881, 
        n52010, n41_adj_4882, n110_adj_4883, n52009, n51050, n51049, 
        n51048, n831_adj_4884, n51820, n52008, n223_adj_4885, n220_adj_4887, 
        n52007, n51047, n52006, n52005, n52004, n52003, n52002, 
        n1096_adj_4888, n52001, n50512, n51046, n51045, n293_adj_4890, 
        n50395, n51044, n1099_adj_4892, n51043, n758_adj_4893, n51819, 
        n1026_adj_4894, n51042, n50511, n953_adj_4896, n51041, n50394, 
        n50510, n50393, n366_adj_4898, n1023_adj_4899, n52000, n66769, 
        n50392, n50509, n880_adj_4902, n51040, n807_adj_4903, n51039, 
        n50508, n50835, n50391, n50834, n734_adj_4905, n51038, n50390, 
        n661_adj_4906, n51037, n1114_adj_4907, n50833, n1041_adj_4908, 
        n50832, n588_adj_4909, n51036, n968_adj_4911, n50831, n895_adj_4912, 
        n50830, n515_adj_4913, n51035, n50507, n685_adj_4915, n51818, 
        n612_adj_4916, n51817, n539_adj_4917, n51816, n442_adj_4918, 
        n51034, n50506, n369_adj_4920, n51033, n50505, n466_adj_4922, 
        n51815, n950_adj_4923, n51999, n877_adj_4924, n51998, n804_adj_4925, 
        n51997, n393_adj_4926, n51814, n731_adj_4927, n51996, n6_adj_4928, 
        n50504, n822_adj_4930, n50829, n296_adj_4931, n51032, n658_adj_4932, 
        n51995, n439_adj_4933, n50503, n585_adj_4935, n51994, n320_adj_4936, 
        n51813, n512_adj_4937, n51993, n51992, n51991, n51990, n51989, 
        n50502, n51031, n51988, n51812, n51030, n51811, n50828, 
        n51810, n67420, n67443, n66619, n66653, n37_adj_4939, n39_adj_4940, 
        n41_adj_4941, n35_adj_4942, n33_adj_4943, n29_adj_4944, n27_adj_4945, 
        n31_adj_4946, n23_adj_4947, n25_adj_4948, n43_adj_4949, n45_adj_4950, 
        n66748, n66716, n12_adj_4952, n10_adj_4953, n30_adj_4954, 
        n67670, n67660, n68905, n68293, n69080, n16_adj_4955, n68347, 
        n68348, n8_adj_4956, n24_adj_4957, n66625, n68285, n67591, 
        n4_adj_4958, n68885, n68886, n66664, n69119, n68595, n69248, 
        n69249, n69217, n66628, n68891, n40_adj_4959, n68893, n37_adj_4960, 
        n39_adj_4961, n35_adj_4962, n33_adj_4963, n29_adj_4964, n31_adj_4965, 
        n27_adj_4966, n45_adj_4967, n23_adj_4968, n25_adj_4969, n43_adj_4970, 
        n66598, n66539, n12_adj_4971, n10_adj_4972, n30_adj_4973, 
        n67500, n67494, n68849, n68215, n69074, n16_adj_4974, n68835, 
        n68836, n8_adj_4975, n24_adj_4976, n67422, n68287, n68599, 
        n4_adj_4977, n68833, n68834, n66505, n69032, n28, n69177, 
        n69178, n69105, n67425, n68895, n67597, n69086, n16_adj_4979, 
        n18_adj_4980, n24_adj_4981, n22_adj_4982, n26_adj_4983;
    wire [2:0]n20183;
    
    SB_CARRY add_6214_9 (.CI(n50826), .I0(n16950[6]), .I1(n603), .CO(n50827));
    SB_CARRY unary_minus_21_add_3_24 (.CI(n50500), .I0(GND_net), .I1(n46[22]), 
            .CO(n50501));
    SB_CARRY add_6349_12 (.CI(n51808), .I0(n18947[9]), .I1(n834), .CO(n51809));
    SB_LUT4 add_6041_22_lut (.I0(GND_net), .I1(n13661[19]), .I2(GND_net), 
            .I3(n51986), .O(n12695[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n46[21]), 
            .I3(n50499), .O(n379[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6214_8_lut (.I0(GND_net), .I1(n16950[5]), .I2(n530), .I3(n50825), 
            .O(n16339[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_5 (.CI(n50388), .I0(n258[3]), .I1(n303[3]), .CO(n50389));
    SB_LUT4 add_19_4_lut (.I0(GND_net), .I1(n258[2]), .I2(n303[2]), .I3(n50387), 
            .O(n353[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_23 (.CI(n50499), .I0(GND_net), .I1(n46[21]), 
            .CO(n50500));
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n46[20]), 
            .I3(n50498), .O(n379[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_22 (.CI(n51986), .I0(n13661[19]), .I1(GND_net), 
            .CO(n51987));
    SB_LUT4 add_6041_21_lut (.I0(GND_net), .I1(n13661[18]), .I2(GND_net), 
            .I3(n51985), .O(n12695[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_21 (.CI(n51985), .I0(n13661[18]), .I1(GND_net), 
            .CO(n51986));
    SB_LUT4 add_6041_20_lut (.I0(GND_net), .I1(n13661[17]), .I2(GND_net), 
            .I3(n51984), .O(n12695[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i7_3_lut (.I0(n48[6]), .I1(n49[6]), .I2(n182), .I3(GND_net), 
            .O(n208[6]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i7_3_lut (.I0(n208[6]), .I1(IntegralLimit[6]), .I2(n156), 
            .I3(GND_net), .O(n233[6]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Kp[1] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Kp[0] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Kp[2] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i373_2_lut (.I0(\Ki[7] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Kp[3] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Kp[4] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Kp[5] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i422_2_lut (.I0(\Ki[8] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Kp[6] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Kp[7] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i15_3_lut (.I0(n48[14]), .I1(n49[14]), .I2(n182), .I3(GND_net), 
            .O(n208[14]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i15_3_lut (.I0(n208[14]), .I1(IntegralLimit[14]), .I2(n156), 
            .I3(GND_net), .O(n233[14]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i471_2_lut (.I0(\Ki[9] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Kp[1] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Kp[0] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6041_20 (.CI(n51984), .I0(n13661[17]), .I1(GND_net), 
            .CO(n51985));
    SB_LUT4 add_6041_19_lut (.I0(GND_net), .I1(n13661[16]), .I2(GND_net), 
            .I3(n51983), .O(n12695[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Kp[2] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4431));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Kp[3] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Kp[4] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Kp[5] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4432));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i85_2_lut (.I0(\Ki[1] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Kp[8] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n50498), .I0(GND_net), .I1(n46[20]), 
            .CO(n50499));
    SB_CARRY add_6041_19 (.CI(n51983), .I0(n13661[16]), .I1(GND_net), 
            .CO(n51984));
    SB_LUT4 mult_17_i469_2_lut (.I0(\Kp[9] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Kp[10] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_18_lut (.I0(GND_net), .I1(n13661[15]), .I2(GND_net), 
            .I3(n51982), .O(n12695[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i134_2_lut (.I0(\Ki[2] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Kp[6] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6349_11_lut (.I0(GND_net), .I1(n18947[8]), .I2(n761), 
            .I3(n51807), .O(n18613[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_11 (.CI(n51807), .I0(n18947[8]), .I1(n761), .CO(n51808));
    SB_LUT4 mult_18_i183_2_lut (.I0(\Ki[3] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Kp[7] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i6_3_lut (.I0(n150), .I1(n49[5]), .I2(n182), .I3(GND_net), 
            .O(n208[5]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i6_3_lut (.I0(n208[5]), .I1(IntegralLimit[5]), .I2(n156), 
            .I3(GND_net), .O(n233[5]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i59_2_lut (.I0(\Ki[1] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i12_2_lut (.I0(\Ki[0] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i232_2_lut (.I0(\Ki[4] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6041_18 (.CI(n51982), .I0(n13661[15]), .I1(GND_net), 
            .CO(n51983));
    SB_LUT4 add_6349_10_lut (.I0(GND_net), .I1(n18947[7]), .I2(n688), 
            .I3(n51806), .O(n18613[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_10 (.CI(n51806), .I0(n18947[7]), .I1(n688), .CO(n51807));
    SB_LUT4 mult_17_i400_2_lut (.I0(\Kp[8] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i108_2_lut (.I0(\Ki[2] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i281_2_lut (.I0(\Ki[5] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n20155[2]), .I1(n6), .I2(n37154), .I3(\Ki[4] ), 
            .O(n20109[3]));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 add_6041_17_lut (.I0(GND_net), .I1(n13661[14]), .I2(GND_net), 
            .I3(n51981), .O(n12695[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_17 (.CI(n51981), .I0(n13661[14]), .I1(GND_net), 
            .CO(n51982));
    SB_LUT4 mult_18_i138_2_lut (.I0(\Ki[2] ), .I1(n233[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_16_lut (.I0(GND_net), .I1(n13661[13]), .I2(n1099), 
            .I3(n51980), .O(n12695[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_16 (.CI(n51980), .I0(n13661[13]), .I1(n1099), .CO(n51981));
    SB_LUT4 add_6349_9_lut (.I0(GND_net), .I1(n18947[6]), .I2(n615), .I3(n51805), 
            .O(n18613[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_9 (.CI(n51805), .I0(n18947[6]), .I1(n615), .CO(n51806));
    SB_LUT4 add_6349_8_lut (.I0(GND_net), .I1(n18947[5]), .I2(n542), .I3(n51804), 
            .O(n18613[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i212_2_lut (.I0(\Ki[4] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36230_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(n233[22]), .I3(n233[21]), 
            .O(n20194));   // verilog/motorControl.v(55[31:42])
    defparam i36230_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_18_i89_2_lut (.I0(\Ki[1] ), .I1(n233[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_15_lut (.I0(GND_net), .I1(n13661[12]), .I2(n1026), 
            .I3(n51979), .O(n12695[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_15 (.CI(n51979), .I0(n13661[12]), .I1(n1026), .CO(n51980));
    SB_LUT4 mult_17_i304_2_lut (.I0(\Kp[6] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_14_lut (.I0(GND_net), .I1(n13661[11]), .I2(n953), 
            .I3(n51978), .O(n12695[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Kp[13] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i261_2_lut (.I0(\Ki[5] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_945 (.I0(n20185), .I1(n4_adj_4434), .I2(\Ki[3] ), 
            .I3(n233[19]), .O(n20155[2]));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h9666;
    SB_LUT4 mux_15_i24_3_lut (.I0(n48[23]), .I1(n49[23]), .I2(n182), .I3(GND_net), 
            .O(n208[23]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Kp[7] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_16_i24_3_lut (.I0(n208[23]), .I1(IntegralLimit[23]), .I2(n156), 
            .I3(GND_net), .O(n233[23]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6041_14 (.CI(n51978), .I0(n13661[11]), .I1(n953), .CO(n51979));
    SB_LUT4 mux_15_i19_3_lut (.I0(n48[18]), .I1(n49[18]), .I2(n182), .I3(GND_net), 
            .O(n214));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i20_3_lut (.I0(n48[19]), .I1(n49[19]), .I2(n182), .I3(GND_net), 
            .O(n208[19]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6214_8 (.CI(n50825), .I0(n16950[5]), .I1(n530), .CO(n50826));
    SB_LUT4 add_6214_7_lut (.I0(GND_net), .I1(n16950[4]), .I2(n457), .I3(n50824), 
            .O(n16339[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Kp[8] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6214_7 (.CI(n50824), .I0(n16950[4]), .I1(n457), .CO(n50825));
    SB_CARRY add_19_4 (.CI(n50387), .I0(n258[2]), .I1(n303[2]), .CO(n50388));
    SB_CARRY add_6349_8 (.CI(n51804), .I0(n18947[5]), .I1(n542), .CO(n51805));
    SB_LUT4 mult_18_i310_2_lut (.I0(\Ki[6] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Kp[14] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_16_i20_3_lut (.I0(n208[19]), .I1(IntegralLimit[19]), .I2(n156), 
            .I3(GND_net), .O(n233[19]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6349_7_lut (.I0(GND_net), .I1(n18947[4]), .I2(n469), .I3(n51803), 
            .O(n18613[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_13_lut (.I0(GND_net), .I1(n13661[10]), .I2(n880), 
            .I3(n51977), .O(n12695[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_13 (.CI(n51977), .I0(n13661[10]), .I1(n880), .CO(n51978));
    SB_LUT4 add_6041_12_lut (.I0(GND_net), .I1(n13661[9]), .I2(n807), 
            .I3(n51976), .O(n12695[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_12 (.CI(n51976), .I0(n13661[9]), .I1(n807), .CO(n51977));
    SB_LUT4 add_6041_11_lut (.I0(GND_net), .I1(n13661[8]), .I2(n734), 
            .I3(n51975), .O(n12695[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_7 (.CI(n51803), .I0(n18947[4]), .I1(n469), .CO(n51804));
    SB_LUT4 add_6349_6_lut (.I0(GND_net), .I1(n18947[3]), .I2(n396), .I3(n51802), 
            .O(n18613[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_11 (.CI(n51975), .I0(n13661[8]), .I1(n734), .CO(n51976));
    SB_LUT4 add_6041_10_lut (.I0(GND_net), .I1(n13661[7]), .I2(n661), 
            .I3(n51974), .O(n12695[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_6 (.CI(n51802), .I0(n18947[3]), .I1(n396), .CO(n51803));
    SB_CARRY add_6041_10 (.CI(n51974), .I0(n13661[7]), .I1(n661), .CO(n51975));
    SB_LUT4 add_6041_9_lut (.I0(GND_net), .I1(n13661[6]), .I2(n588), .I3(n51973), 
            .O(n12695[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6214_6_lut (.I0(GND_net), .I1(n16950[3]), .I2(n384), .I3(n50823), 
            .O(n16339[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF control_update_40 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_LUT4 mux_15_i22_3_lut (.I0(n48[21]), .I1(n49[21]), .I2(n182), .I3(GND_net), 
            .O(n208[21]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i22_3_lut (.I0(n208[21]), .I1(IntegralLimit[21]), .I2(n156), 
            .I3(GND_net), .O(n233[21]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i23_3_lut (.I0(n48[22]), .I1(n49[22]), .I2(n182), .I3(GND_net), 
            .O(n208[22]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i23_3_lut (.I0(n208[22]), .I1(IntegralLimit[22]), .I2(n156), 
            .I3(GND_net), .O(n233[22]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER result_i0 (.Q(duty[0]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[0]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_LUT4 mult_18_i330_2_lut (.I0(\Ki[6] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6214_6 (.CI(n50823), .I0(n16950[3]), .I1(n384), .CO(n50824));
    SB_LUT4 add_6349_5_lut (.I0(GND_net), .I1(n18947[2]), .I2(n323), .I3(n51801), 
            .O(n18613[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_5 (.CI(n51801), .I0(n18947[2]), .I1(n323), .CO(n51802));
    SB_CARRY add_6041_9 (.CI(n51973), .I0(n13661[6]), .I1(n588), .CO(n51974));
    SB_LUT4 add_6349_4_lut (.I0(GND_net), .I1(n18947[1]), .I2(n250_adj_4436), 
            .I3(n51800), .O(n18613[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\Ki[2] ), .I1(\Ki[1] ), .I2(n233[21]), 
            .I3(n233[22]), .O(n62866));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h6ca0;
    SB_CARRY add_6349_4 (.CI(n51800), .I0(n18947[1]), .I1(n250_adj_4436), 
            .CO(n51801));
    SB_LUT4 add_6214_5_lut (.I0(GND_net), .I1(n16950[2]), .I2(n311), .I3(n50822), 
            .O(n16339[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_947 (.I0(\Ki[4] ), .I1(n37050), .I2(n233[19]), 
            .I3(\Ki[3] ), .O(n62868));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_6349_3_lut (.I0(GND_net), .I1(n18947[0]), .I2(n177), .I3(n51799), 
            .O(n18613[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_8_lut (.I0(GND_net), .I1(n13661[5]), .I2(n515), .I3(n51972), 
            .O(n12695[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_3 (.CI(n51799), .I0(n18947[0]), .I1(n177), .CO(n51800));
    SB_CARRY add_6041_8 (.CI(n51972), .I0(n13661[5]), .I1(n515), .CO(n51973));
    SB_LUT4 add_6041_7_lut (.I0(GND_net), .I1(n13661[4]), .I2(n442), .I3(n51971), 
            .O(n12695[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6349_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n18613[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_5 (.CI(n50822), .I0(n16950[2]), .I1(n311), .CO(n50823));
    SB_LUT4 i36232_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(n233[22]), .I3(n233[21]), 
            .O(n50153));   // verilog/motorControl.v(55[31:42])
    defparam i36232_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n37154), .I1(\Ki[0] ), .I2(\Ki[5] ), 
            .I3(n233[23]), .O(n62856));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h93a0;
    SB_LUT4 mult_18_i359_2_lut (.I0(\Ki[7] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6041_7 (.CI(n51971), .I0(n13661[4]), .I1(n442), .CO(n51972));
    SB_LUT4 add_6041_6_lut (.I0(GND_net), .I1(n13661[3]), .I2(n369), .I3(n51970), 
            .O(n12695[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_6 (.CI(n51970), .I0(n13661[3]), .I1(n369), .CO(n51971));
    SB_CARRY add_6349_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n51799));
    SB_LUT4 i36125_4_lut (.I0(n20155[2]), .I1(n37154), .I2(n6), .I3(\Ki[4] ), 
            .O(n8));   // verilog/motorControl.v(55[31:42])
    defparam i36125_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i36324_4_lut (.I0(n20185), .I1(\Ki[3] ), .I2(n4_adj_4434), 
            .I3(n233[19]), .O(n6_adj_4437));   // verilog/motorControl.v(55[31:42])
    defparam i36324_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n4), .I1(n50153), .I2(n62868), .I3(n62866), 
            .O(n62874));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n62874), .I1(n6_adj_4437), .I2(n8), 
            .I3(n62856), .O(n60827));   // verilog/motorControl.v(55[31:42])
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 add_6214_4_lut (.I0(GND_net), .I1(n16950[1]), .I2(n238_adj_4439), 
            .I3(n50821), .O(n16339[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_19_3_lut (.I0(GND_net), .I1(n258[1]), .I2(n303[1]), .I3(n50386), 
            .O(n353[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_4 (.CI(n50821), .I0(n16950[1]), .I1(n238_adj_4439), 
            .CO(n50822));
    SB_LUT4 add_6454_8_lut (.I0(GND_net), .I1(n19980[5]), .I2(n560), .I3(n51798), 
            .O(n19869[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_5_lut (.I0(GND_net), .I1(n13661[2]), .I2(n296), .I3(n51969), 
            .O(n12695[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_3 (.CI(n50386), .I0(n258[1]), .I1(n303[1]), .CO(n50387));
    SB_LUT4 add_6214_3_lut (.I0(GND_net), .I1(n16950[0]), .I2(n165), .I3(n50820), 
            .O(n16339[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_3 (.CI(n50820), .I0(n16950[0]), .I1(n165), .CO(n50821));
    SB_LUT4 mult_18_i157_2_lut (.I0(\Ki[3] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6454_7_lut (.I0(GND_net), .I1(n19980[4]), .I2(n487), .I3(n51797), 
            .O(n19869[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6214_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n16339[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i408_2_lut (.I0(\Ki[8] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n46[19]), 
            .I3(n50497), .O(n379[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Kp[9] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i457_2_lut (.I0(\Ki[9] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_19_2_lut (.I0(GND_net), .I1(n258[0]), .I2(n303[0]), .I3(GND_net), 
            .O(n353[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Kp[9] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6454_7 (.CI(n51797), .I0(n19980[4]), .I1(n487), .CO(n51798));
    SB_CARRY unary_minus_21_add_3_21 (.CI(n50497), .I0(GND_net), .I1(n46[19]), 
            .CO(n50498));
    SB_CARRY add_6214_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n50820));
    SB_LUT4 mult_17_i69_2_lut (.I0(\Kp[1] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n46[18]), 
            .I3(n50496), .O(n379[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_5 (.CI(n51969), .I0(n13661[2]), .I1(n296), .CO(n51970));
    SB_LUT4 add_6454_6_lut (.I0(GND_net), .I1(n19980[3]), .I2(n414), .I3(n51796), 
            .O(n19869[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_20 (.CI(n50496), .I0(GND_net), .I1(n46[18]), 
            .CO(n50497));
    SB_LUT4 mult_17_i22_2_lut (.I0(\Kp[0] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_4_lut (.I0(GND_net), .I1(n13661[1]), .I2(n223), .I3(n51968), 
            .O(n12695[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i206_2_lut (.I0(\Ki[4] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6041_4 (.CI(n51968), .I0(n13661[1]), .I1(n223), .CO(n51969));
    SB_LUT4 mult_17_i118_2_lut (.I0(\Kp[2] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n46[17]), 
            .I3(n50495), .O(n379[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Kp[10] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6454_6 (.CI(n51796), .I0(n19980[3]), .I1(n414), .CO(n51797));
    SB_CARRY add_19_2 (.CI(GND_net), .I0(n258[0]), .I1(n303[0]), .CO(n50386));
    SB_LUT4 mult_17_i167_2_lut (.I0(\Kp[3] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_3_lut (.I0(GND_net), .I1(n13661[0]), .I2(n150_adj_4444), 
            .I3(n51967), .O(n12695[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_5_lut (.I0(GND_net), .I1(n19980[2]), .I2(n341), .I3(n51795), 
            .O(n19869[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i255_2_lut (.I0(\Ki[5] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_21_add_3_19 (.CI(n50495), .I0(GND_net), .I1(n46[17]), 
            .CO(n50496));
    SB_LUT4 add_10_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n105[23]), .I3(n50385), .O(n48[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Kp[11] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Kp[4] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n46[16]), 
            .I3(n50494), .O(n379[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_18 (.CI(n50494), .I0(GND_net), .I1(n46[16]), 
            .CO(n50495));
    SB_LUT4 add_10_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n105[23]), .I3(n50384), .O(n48[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Kp[12] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n46[15]), 
            .I3(n50493), .O(n379[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Kp[5] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6041_3 (.CI(n51967), .I0(n13661[0]), .I1(n150_adj_4444), 
            .CO(n51968));
    SB_LUT4 add_6041_2_lut (.I0(GND_net), .I1(n8_adj_4446), .I2(n77), 
            .I3(GND_net), .O(n12695[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i304_2_lut (.I0(\Ki[6] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4447));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Kp[6] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Kp[7] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Kp[13] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6454_5 (.CI(n51795), .I0(n19980[2]), .I1(n341), .CO(n51796));
    SB_CARRY add_6041_2 (.CI(GND_net), .I0(n8_adj_4446), .I1(n77), .CO(n51967));
    SB_LUT4 add_6085_22_lut (.I0(GND_net), .I1(n14539[19]), .I2(GND_net), 
            .I3(n51966), .O(n13661[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Kp[8] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Kp[14] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Kp[9] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_28_i2_3_lut (.I0(n353[1]), .I1(n433[1]), .I2(n432), .I3(GND_net), 
            .O(n458[1]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i2_3_lut (.I0(n458[1]), .I1(PWMLimit[1]), .I2(n406), 
            .I3(GND_net), .O(n483[1]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_4_lut (.I0(setpoint[1]), .I1(n483[1]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[1]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i2_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i27582_3_lut (.I0(n353[2]), .I1(n433[2]), .I2(n432), .I3(GND_net), 
            .O(n1));
    defparam i27582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27584_3_lut (.I0(n1), .I1(PWMLimit[2]), .I2(n406), .I3(GND_net), 
            .O(n3_adj_4449));
    defparam i27584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27585_4_lut (.I0(setpoint[2]), .I1(n3_adj_4449), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[2]));
    defparam i27585_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_28_i4_3_lut (.I0(n353[3]), .I1(n433[3]), .I2(n432), .I3(GND_net), 
            .O(n458[3]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i4_3_lut (.I0(n458[3]), .I1(PWMLimit[3]), .I2(n406), 
            .I3(GND_net), .O(n483[3]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Kp[15] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(setpoint[3]), .I1(n483[3]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[3]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_6454_4_lut (.I0(GND_net), .I1(n19980[1]), .I2(n268), .I3(n51794), 
            .O(n19869[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_17 (.CI(n50493), .I0(GND_net), .I1(n46[15]), 
            .CO(n50494));
    SB_CARRY add_10_24 (.CI(n50384), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n105[23]), .CO(n50385));
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n46[14]), 
            .I3(n50492), .O(n379[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_16 (.CI(n50492), .I0(GND_net), .I1(n46[14]), 
            .CO(n50493));
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n46[13]), 
            .I3(n50491), .O(n379[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n105[23]), .I3(n50383), .O(n48[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_15 (.CI(n50491), .I0(GND_net), .I1(n46[13]), 
            .CO(n50492));
    SB_LUT4 mux_28_i5_3_lut (.I0(n353[4]), .I1(n433[4]), .I2(n432), .I3(GND_net), 
            .O(n478));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6085_21_lut (.I0(GND_net), .I1(n14539[18]), .I2(GND_net), 
            .I3(n51965), .O(n13661[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n46[12]), 
            .I3(n50490), .O(n379[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i6_3_lut (.I0(n353[5]), .I1(n433[5]), .I2(n432), .I3(GND_net), 
            .O(n458[5]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Kp[10] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_10_23 (.CI(n50383), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n105[23]), .CO(n50384));
    SB_CARRY unary_minus_21_add_3_14 (.CI(n50490), .I0(GND_net), .I1(n46[12]), 
            .CO(n50491));
    SB_LUT4 add_10_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n105[23]), .I3(n50382), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_4 (.CI(n51794), .I0(n19980[1]), .I1(n268), .CO(n51795));
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n46[11]), 
            .I3(n50489), .O(n379[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_22 (.CI(n50382), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n105[23]), .CO(n50383));
    SB_CARRY unary_minus_21_add_3_13 (.CI(n50489), .I0(GND_net), .I1(n46[11]), 
            .CO(n50490));
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n46[10]), 
            .I3(n50488), .O(n379[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_3_lut (.I0(GND_net), .I1(n19980[0]), .I2(n195), .I3(n51793), 
            .O(n19869[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i353_2_lut (.I0(\Ki[7] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4454));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_10_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n105[23]), .I3(n50381), .O(n48[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_21 (.CI(n50381), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n105[23]), .CO(n50382));
    SB_CARRY unary_minus_21_add_3_12 (.CI(n50488), .I0(GND_net), .I1(n46[10]), 
            .CO(n50489));
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n46[9]), 
            .I3(n50487), .O(n379[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_29_i6_3_lut (.I0(n458[5]), .I1(PWMLimit[5]), .I2(n406), 
            .I3(GND_net), .O(n483[5]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6085_21 (.CI(n51965), .I0(n14539[18]), .I1(GND_net), 
            .CO(n51966));
    SB_LUT4 duty_23__I_0_i6_4_lut (.I0(setpoint[5]), .I1(n483[5]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[5]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i6_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_10_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n105[22]), .I3(n50380), .O(n48[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n50487), .I0(GND_net), .I1(n46[9]), 
            .CO(n50488));
    SB_CARRY add_10_20 (.CI(n50380), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n105[22]), .CO(n50381));
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n46[8]), 
            .I3(n50486), .O(n379[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i7_3_lut (.I0(n353[6]), .I1(n433[6]), .I2(n432), .I3(GND_net), 
            .O(n458[6]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n50486), .I0(GND_net), .I1(n46[8]), 
            .CO(n50487));
    SB_LUT4 add_10_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n105[21]), .I3(n50379), .O(n48[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n46[7]), 
            .I3(n50485), .O(n379[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_29_i7_3_lut (.I0(n458[6]), .I1(PWMLimit[6]), .I2(n406), 
            .I3(GND_net), .O(n483[6]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n50485), .I0(GND_net), .I1(n46[7]), 
            .CO(n50486));
    SB_CARRY add_10_19 (.CI(n50379), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n105[21]), .CO(n50380));
    SB_LUT4 mult_18_i402_2_lut (.I0(\Ki[8] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4458));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_10_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n105[20]), .I3(n50378), .O(n48[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Kp[11] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_10_18 (.CI(n50378), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n105[20]), .CO(n50379));
    SB_CARRY add_6454_3 (.CI(n51793), .I0(n19980[0]), .I1(n195), .CO(n51794));
    SB_LUT4 add_6454_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_4459), 
            .I3(GND_net), .O(n19869[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i7_4_lut (.I0(setpoint[6]), .I1(n483[6]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[6]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_6454_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_4459), .CO(n51793));
    SB_LUT4 add_6247_17_lut (.I0(GND_net), .I1(n17493[14]), .I2(GND_net), 
            .I3(n50801), .O(n16950[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n46[6]), 
            .I3(n50484), .O(n379[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6247_16_lut (.I0(GND_net), .I1(n17493[13]), .I2(n1117), 
            .I3(n50800), .O(n16950[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6373_13_lut (.I0(GND_net), .I1(n19231[10]), .I2(n910), 
            .I3(n51792), .O(n18947[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i8_3_lut (.I0(n353[7]), .I1(n433[7]), .I2(n432), .I3(GND_net), 
            .O(n458[7]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n50484), .I0(GND_net), .I1(n46[6]), 
            .CO(n50485));
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n46[5]), 
            .I3(n50483), .O(n379[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_16 (.CI(n50800), .I0(n17493[13]), .I1(n1117), .CO(n50801));
    SB_LUT4 add_6247_15_lut (.I0(GND_net), .I1(n17493[12]), .I2(n1044), 
            .I3(n50799), .O(n16950[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_15 (.CI(n50799), .I0(n17493[12]), .I1(n1044), .CO(n50800));
    SB_LUT4 add_6247_14_lut (.I0(GND_net), .I1(n17493[11]), .I2(n971), 
            .I3(n50798), .O(n16950[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_14 (.CI(n50798), .I0(n17493[11]), .I1(n971), .CO(n50799));
    SB_LUT4 mux_29_i8_3_lut (.I0(n458[7]), .I1(PWMLimit[7]), .I2(n406), 
            .I3(GND_net), .O(n500));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_28_i9_3_lut (.I0(n353[8]), .I1(n433[8]), .I2(n432), .I3(GND_net), 
            .O(n458[8]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i9_3_lut (.I0(n458[8]), .I1(PWMLimit[8]), .I2(n406), 
            .I3(GND_net), .O(n483[8]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_14_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[0]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_i9_4_lut (.I0(setpoint[8]), .I1(n483[8]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[8]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i9_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Kp[1] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Kp[0] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_28_i10_3_lut (.I0(n353[9]), .I1(n433[9]), .I2(n432), .I3(GND_net), 
            .O(n458[9]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6373_12_lut (.I0(GND_net), .I1(n19231[9]), .I2(n837), 
            .I3(n51791), .O(n18947[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_20_lut (.I0(GND_net), .I1(n14539[17]), .I2(GND_net), 
            .I3(n51964), .O(n13661[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_20 (.CI(n51964), .I0(n14539[17]), .I1(GND_net), 
            .CO(n51965));
    SB_LUT4 add_6085_19_lut (.I0(GND_net), .I1(n14539[16]), .I2(GND_net), 
            .I3(n51963), .O(n13661[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_29_i10_3_lut (.I0(n458[9]), .I1(PWMLimit[9]), .I2(n406), 
            .I3(GND_net), .O(n483[9]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Kp[6] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6247_13_lut (.I0(GND_net), .I1(n17493[10]), .I2(n898), 
            .I3(n50797), .O(n16950[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_13 (.CI(n50797), .I0(n17493[10]), .I1(n898), .CO(n50798));
    SB_LUT4 add_6247_12_lut (.I0(GND_net), .I1(n17493[9]), .I2(n825), 
            .I3(n50796), .O(n16950[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i10_4_lut (.I0(setpoint[9]), .I1(n483[9]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[9]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i10_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Kp[12] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6247_12 (.CI(n50796), .I0(n17493[9]), .I1(n825), .CO(n50797));
    SB_LUT4 add_6247_11_lut (.I0(GND_net), .I1(n17493[8]), .I2(n752), 
            .I3(n50795), .O(n16950[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_7 (.CI(n50483), .I0(GND_net), .I1(n46[5]), 
            .CO(n50484));
    SB_LUT4 mult_17_i657_2_lut (.I0(\Kp[13] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Kp[14] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Kp[2] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6247_11 (.CI(n50795), .I0(n17493[8]), .I1(n752), .CO(n50796));
    SB_LUT4 add_6247_10_lut (.I0(GND_net), .I1(n17493[7]), .I2(n679_adj_4462), 
            .I3(n50794), .O(n16950[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6061_22_lut (.I0(GND_net), .I1(n14058[19]), .I2(GND_net), 
            .I3(n51006), .O(n13134[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6373_12 (.CI(n51791), .I0(n19231[9]), .I1(n837), .CO(n51792));
    SB_LUT4 add_10_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n105[19]), .I3(n50377), .O(n48[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_10 (.CI(n50794), .I0(n17493[7]), .I1(n679_adj_4462), 
            .CO(n50795));
    SB_LUT4 add_6061_21_lut (.I0(GND_net), .I1(n14058[18]), .I2(GND_net), 
            .I3(n51005), .O(n13134[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i11_3_lut (.I0(n353[10]), .I1(n433[10]), .I2(n432), 
            .I3(GND_net), .O(n458[10]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6085_19 (.CI(n51963), .I0(n14539[16]), .I1(GND_net), 
            .CO(n51964));
    SB_CARRY add_6061_21 (.CI(n51005), .I0(n14058[18]), .I1(GND_net), 
            .CO(n51006));
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n46[4]), 
            .I3(n50482), .O(n379[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_29_i11_3_lut (.I0(n458[10]), .I1(PWMLimit[10]), .I2(n406), 
            .I3(GND_net), .O(n483[10]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6373_11_lut (.I0(GND_net), .I1(n19231[8]), .I2(n764), 
            .I3(n51790), .O(n18947[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6247_9_lut (.I0(GND_net), .I1(n17493[6]), .I2(n606_adj_4463), 
            .I3(n50793), .O(n16950[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6373_11 (.CI(n51790), .I0(n19231[8]), .I1(n764), .CO(n51791));
    SB_CARRY add_6247_9 (.CI(n50793), .I0(n17493[6]), .I1(n606_adj_4463), 
            .CO(n50794));
    SB_LUT4 add_6373_10_lut (.I0(GND_net), .I1(n19231[7]), .I2(n691), 
            .I3(n51789), .O(n18947[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6373_10 (.CI(n51789), .I0(n19231[7]), .I1(n691), .CO(n51790));
    SB_LUT4 add_6373_9_lut (.I0(GND_net), .I1(n19231[6]), .I2(n618), .I3(n51788), 
            .O(n18947[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_18_lut (.I0(GND_net), .I1(n14539[15]), .I2(GND_net), 
            .I3(n51962), .O(n13661[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i11_4_lut (.I0(setpoint[10]), .I1(n483[10]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[10]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i11_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_28_i12_3_lut (.I0(n353[11]), .I1(n433[11]), .I2(n432), 
            .I3(GND_net), .O(n458[11]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i12_3_lut (.I0(n458[11]), .I1(PWMLimit[11]), .I2(n406), 
            .I3(GND_net), .O(n483[11]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6085_18 (.CI(n51962), .I0(n14539[15]), .I1(GND_net), 
            .CO(n51963));
    SB_CARRY add_6373_9 (.CI(n51788), .I0(n19231[6]), .I1(n618), .CO(n51789));
    SB_LUT4 add_6085_17_lut (.I0(GND_net), .I1(n14539[14]), .I2(GND_net), 
            .I3(n51961), .O(n13661[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_17 (.CI(n51961), .I0(n14539[14]), .I1(GND_net), 
            .CO(n51962));
    SB_LUT4 add_6061_20_lut (.I0(GND_net), .I1(n14058[17]), .I2(GND_net), 
            .I3(n51004), .O(n13134[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6247_8_lut (.I0(GND_net), .I1(n17493[5]), .I2(n533_adj_4464), 
            .I3(n50792), .O(n16950[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_6 (.CI(n50482), .I0(GND_net), .I1(n46[4]), 
            .CO(n50483));
    SB_LUT4 duty_23__I_0_i12_4_lut (.I0(setpoint[11]), .I1(n483[11]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[11]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i12_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_6061_20 (.CI(n51004), .I0(n14058[17]), .I1(GND_net), 
            .CO(n51005));
    SB_CARRY add_10_17 (.CI(n50377), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n105[19]), .CO(n50378));
    SB_LUT4 add_6085_16_lut (.I0(GND_net), .I1(n14539[13]), .I2(n1102), 
            .I3(n51960), .O(n13661[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6061_19_lut (.I0(GND_net), .I1(n14058[16]), .I2(GND_net), 
            .I3(n51003), .O(n13134[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_19 (.CI(n51003), .I0(n14058[16]), .I1(GND_net), 
            .CO(n51004));
    SB_LUT4 add_10_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n105[18]), .I3(n50376), .O(n48[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_16 (.CI(n51960), .I0(n14539[13]), .I1(n1102), .CO(n51961));
    SB_CARRY add_6247_8 (.CI(n50792), .I0(n17493[5]), .I1(n533_adj_4464), 
            .CO(n50793));
    SB_LUT4 add_6247_7_lut (.I0(GND_net), .I1(n17493[4]), .I2(n460_adj_4465), 
            .I3(n50791), .O(n16950[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_15_lut (.I0(GND_net), .I1(n14539[12]), .I2(n1029), 
            .I3(n51959), .O(n13661[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_7 (.CI(n50791), .I0(n17493[4]), .I1(n460_adj_4465), 
            .CO(n50792));
    SB_LUT4 add_6061_18_lut (.I0(GND_net), .I1(n14058[15]), .I2(GND_net), 
            .I3(n51002), .O(n13134[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n46[3]), 
            .I3(n50481), .O(n379[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6247_6_lut (.I0(GND_net), .I1(n17493[3]), .I2(n387_adj_4466), 
            .I3(n50790), .O(n16950[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n50481), .I0(GND_net), .I1(n46[3]), 
            .CO(n50482));
    SB_CARRY add_6247_6 (.CI(n50790), .I0(n17493[3]), .I1(n387_adj_4466), 
            .CO(n50791));
    SB_CARRY add_10_16 (.CI(n50376), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n105[18]), .CO(n50377));
    SB_LUT4 add_10_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n105[17]), .I3(n50375), .O(n48[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6247_5_lut (.I0(GND_net), .I1(n17493[2]), .I2(n314_adj_4467), 
            .I3(n50789), .O(n16950[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n46[2]), 
            .I3(n50480), .O(n379[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6373_8_lut (.I0(GND_net), .I1(n19231[5]), .I2(n545), .I3(n51787), 
            .O(n18947[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_15 (.CI(n50375), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n105[17]), .CO(n50376));
    SB_CARRY add_6247_5 (.CI(n50789), .I0(n17493[2]), .I1(n314_adj_4467), 
            .CO(n50790));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n50480), .I0(GND_net), .I1(n46[2]), 
            .CO(n50481));
    SB_LUT4 add_10_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n105[16]), .I3(n50374), .O(n48[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_18 (.CI(n51002), .I0(n14058[15]), .I1(GND_net), 
            .CO(n51003));
    SB_LUT4 add_6247_4_lut (.I0(GND_net), .I1(n17493[1]), .I2(n241), .I3(n50788), 
            .O(n16950[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n46[1]), 
            .I3(n50479), .O(n379[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_15 (.CI(n51959), .I0(n14539[12]), .I1(n1029), .CO(n51960));
    SB_CARRY add_6373_8 (.CI(n51787), .I0(n19231[5]), .I1(n545), .CO(n51788));
    SB_LUT4 add_6373_7_lut (.I0(GND_net), .I1(n19231[4]), .I2(n472_adj_4470), 
            .I3(n51786), .O(n18947[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_14_lut (.I0(GND_net), .I1(n14539[11]), .I2(n956), 
            .I3(n51958), .O(n13661[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_14 (.CI(n51958), .I0(n14539[11]), .I1(n956), .CO(n51959));
    SB_CARRY unary_minus_21_add_3_3 (.CI(n50479), .I0(GND_net), .I1(n46[1]), 
            .CO(n50480));
    SB_CARRY add_6373_7 (.CI(n51786), .I0(n19231[4]), .I1(n472_adj_4470), 
            .CO(n51787));
    SB_LUT4 add_6085_13_lut (.I0(GND_net), .I1(n14539[10]), .I2(n883), 
            .I3(n51957), .O(n13661[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i13_3_lut (.I0(n353[12]), .I1(n433[12]), .I2(n432), 
            .I3(GND_net), .O(n458[12]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6247_4 (.CI(n50788), .I0(n17493[1]), .I1(n241), .CO(n50789));
    SB_LUT4 add_6247_3_lut (.I0(GND_net), .I1(n17493[0]), .I2(n168), .I3(n50787), 
            .O(n16950[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_29_i13_3_lut (.I0(n458[12]), .I1(PWMLimit[12]), .I2(n406), 
            .I3(GND_net), .O(n483[12]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i451_2_lut (.I0(\Ki[9] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4471));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i451_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6085_13 (.CI(n51957), .I0(n14539[10]), .I1(n883), .CO(n51958));
    SB_LUT4 add_6085_12_lut (.I0(GND_net), .I1(n14539[9]), .I2(n810), 
            .I3(n51956), .O(n13661[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i13_4_lut (.I0(setpoint[12]), .I1(n483[12]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[12]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i13_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mult_18_i500_2_lut (.I0(\Ki[10] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_28_i14_3_lut (.I0(n353[13]), .I1(n433[13]), .I2(n432), 
            .I3(GND_net), .O(n458[13]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i14_3_lut (.I0(n458[13]), .I1(PWMLimit[13]), .I2(n406), 
            .I3(GND_net), .O(n483[13]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6373_6_lut (.I0(GND_net), .I1(n19231[3]), .I2(n399_adj_4473), 
            .I3(n51785), .O(n18947[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6373_6 (.CI(n51785), .I0(n19231[3]), .I1(n399_adj_4473), 
            .CO(n51786));
    SB_LUT4 duty_23__I_0_i14_4_lut (.I0(setpoint[13]), .I1(n483[13]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[13]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i14_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_28_i15_3_lut (.I0(n353[14]), .I1(n433[14]), .I2(n432), 
            .I3(GND_net), .O(n458[14]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6085_12 (.CI(n51956), .I0(n14539[9]), .I1(n810), .CO(n51957));
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n42898), .I1(GND_net), .I2(n46[0]), 
            .I3(VCC_net), .O(n66320)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_29_i15_3_lut (.I0(n458[14]), .I1(PWMLimit[14]), .I2(n406), 
            .I3(GND_net), .O(n483[14]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_4_lut (.I0(setpoint[14]), .I1(n483[14]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[14]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i15_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 unary_minus_14_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[1]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6373_5_lut (.I0(GND_net), .I1(n19231[2]), .I2(n326), .I3(n51784), 
            .O(n18947[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i16_3_lut (.I0(n353[15]), .I1(n433[15]), .I2(n432), 
            .I3(GND_net), .O(n458[15]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n46[0]), 
            .CO(n50479));
    SB_CARRY add_6247_3 (.CI(n50787), .I0(n17493[0]), .I1(n168), .CO(n50788));
    SB_LUT4 add_6061_17_lut (.I0(GND_net), .I1(n14058[14]), .I2(GND_net), 
            .I3(n51001), .O(n13134[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6247_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n16950[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6247_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_17 (.CI(n51001), .I0(n14058[14]), .I1(GND_net), 
            .CO(n51002));
    SB_CARRY add_6373_5 (.CI(n51784), .I0(n19231[2]), .I1(n326), .CO(n51785));
    SB_LUT4 add_6061_16_lut (.I0(GND_net), .I1(n14058[13]), .I2(n1102_adj_4477), 
            .I3(n51000), .O(n13134[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6247_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n50787));
    SB_CARRY add_6061_16 (.CI(n51000), .I0(n14058[13]), .I1(n1102_adj_4477), 
            .CO(n51001));
    SB_CARRY add_10_14 (.CI(n50374), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n105[16]), .CO(n50375));
    SB_LUT4 add_6085_11_lut (.I0(GND_net), .I1(n14539[8]), .I2(n737), 
            .I3(n51955), .O(n13661[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6463_8_lut (.I0(GND_net), .I1(n20041[5]), .I2(n560_adj_4478), 
            .I3(n50786), .O(n19947[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6061_15_lut (.I0(GND_net), .I1(n14058[12]), .I2(n1029_adj_4479), 
            .I3(n50999), .O(n13134[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_29_i16_3_lut (.I0(n458[15]), .I1(PWMLimit[15]), .I2(n406), 
            .I3(GND_net), .O(n483[15]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_4_lut (.I0(setpoint[15]), .I1(n483[15]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[15]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i16_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_6085_11 (.CI(n51955), .I0(n14539[8]), .I1(n737), .CO(n51956));
    SB_LUT4 add_6463_7_lut (.I0(GND_net), .I1(n20041[4]), .I2(n487_adj_4480), 
            .I3(n50785), .O(n19947[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_15 (.CI(n50999), .I0(n14058[12]), .I1(n1029_adj_4479), 
            .CO(n51000));
    SB_LUT4 add_6061_14_lut (.I0(GND_net), .I1(n14058[11]), .I2(n956_adj_4481), 
            .I3(n50998), .O(n13134[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n105[15]), .I3(n50373), .O(n48[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_7 (.CI(n50785), .I0(n20041[4]), .I1(n487_adj_4480), 
            .CO(n50786));
    SB_LUT4 add_6463_6_lut (.I0(GND_net), .I1(n20041[3]), .I2(n414_adj_4482), 
            .I3(n50784), .O(n19947[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_13 (.CI(n50373), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n105[15]), .CO(n50374));
    SB_LUT4 unary_minus_14_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n51[23]), 
            .I3(n50478), .O(n49[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6373_4_lut (.I0(GND_net), .I1(n19231[1]), .I2(n253_adj_4483), 
            .I3(n51783), .O(n18947[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6373_4 (.CI(n51783), .I0(n19231[1]), .I1(n253_adj_4483), 
            .CO(n51784));
    SB_LUT4 mux_28_i17_3_lut (.I0(n353[16]), .I1(n433[16]), .I2(n432), 
            .I3(GND_net), .O(n458[16]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6061_14 (.CI(n50998), .I0(n14058[11]), .I1(n956_adj_4481), 
            .CO(n50999));
    SB_CARRY add_6463_6 (.CI(n50784), .I0(n20041[3]), .I1(n414_adj_4482), 
            .CO(n50785));
    SB_LUT4 mux_29_i17_3_lut (.I0(n458[16]), .I1(PWMLimit[16]), .I2(n406), 
            .I3(GND_net), .O(n483[16]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6463_5_lut (.I0(GND_net), .I1(n20041[2]), .I2(n341_adj_4485), 
            .I3(n50783), .O(n19947[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_10_lut (.I0(GND_net), .I1(n14539[7]), .I2(n664), 
            .I3(n51954), .O(n13661[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_5 (.CI(n50783), .I0(n20041[2]), .I1(n341_adj_4485), 
            .CO(n50784));
    SB_LUT4 unary_minus_14_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n51[22]), 
            .I3(n50477), .O(n49[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6373_3_lut (.I0(GND_net), .I1(n19231[0]), .I2(n180), .I3(n51782), 
            .O(n18947[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6463_4_lut (.I0(GND_net), .I1(n20041[1]), .I2(n268_adj_4487), 
            .I3(n50782), .O(n19947[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n105[14]), .I3(n50372), .O(n48[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_10 (.CI(n51954), .I0(n14539[7]), .I1(n664), .CO(n51955));
    SB_CARRY unary_minus_14_add_3_24 (.CI(n50477), .I0(GND_net), .I1(n51[22]), 
            .CO(n50478));
    SB_CARRY add_6463_4 (.CI(n50782), .I0(n20041[1]), .I1(n268_adj_4487), 
            .CO(n50783));
    SB_LUT4 add_6061_13_lut (.I0(GND_net), .I1(n14058[10]), .I2(n883_adj_4488), 
            .I3(n50997), .O(n13134[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_12 (.CI(n50372), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n105[14]), .CO(n50373));
    SB_LUT4 unary_minus_14_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n51[21]), 
            .I3(n50476), .O(n49[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_23 (.CI(n50476), .I0(GND_net), .I1(n51[21]), 
            .CO(n50477));
    SB_CARRY add_6061_13 (.CI(n50997), .I0(n14058[10]), .I1(n883_adj_4488), 
            .CO(n50998));
    SB_CARRY add_6373_3 (.CI(n51782), .I0(n19231[0]), .I1(n180), .CO(n51783));
    SB_LUT4 add_6061_12_lut (.I0(GND_net), .I1(n14058[9]), .I2(n810_adj_4490), 
            .I3(n50996), .O(n13134[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6463_3_lut (.I0(GND_net), .I1(n20041[0]), .I2(n195_adj_4491), 
            .I3(n50781), .O(n19947[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_9_lut (.I0(GND_net), .I1(n14539[6]), .I2(n591), .I3(n51953), 
            .O(n13661[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_12 (.CI(n50996), .I0(n14058[9]), .I1(n810_adj_4490), 
            .CO(n50997));
    SB_LUT4 add_6061_11_lut (.I0(GND_net), .I1(n14058[8]), .I2(n737_adj_4492), 
            .I3(n50995), .O(n13134[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_9 (.CI(n51953), .I0(n14539[6]), .I1(n591), .CO(n51954));
    SB_CARRY add_6463_3 (.CI(n50781), .I0(n20041[0]), .I1(n195_adj_4491), 
            .CO(n50782));
    SB_LUT4 add_6463_2_lut (.I0(GND_net), .I1(n53_adj_4493), .I2(n122_adj_4494), 
            .I3(GND_net), .O(n19947[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n51[20]), 
            .I3(n50475), .O(n187)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n105[13]), .I3(n50371), .O(n48[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_8_lut (.I0(GND_net), .I1(n14539[5]), .I2(n518), .I3(n51952), 
            .O(n13661[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_22 (.CI(n50475), .I0(GND_net), .I1(n51[20]), 
            .CO(n50476));
    SB_CARRY add_6463_2 (.CI(GND_net), .I0(n53_adj_4493), .I1(n122_adj_4494), 
            .CO(n50781));
    SB_CARRY add_10_11 (.CI(n50371), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n105[13]), .CO(n50372));
    SB_CARRY add_6061_11 (.CI(n50995), .I0(n14058[8]), .I1(n737_adj_4492), 
            .CO(n50996));
    SB_LUT4 unary_minus_14_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n51[19]), 
            .I3(n50474), .O(n49[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6373_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_4497), 
            .I3(GND_net), .O(n18947[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6373_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n105[12]), .I3(n50370), .O(n48[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_10 (.CI(n50370), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n105[12]), .CO(n50371));
    SB_CARRY add_6085_8 (.CI(n51952), .I0(n14539[5]), .I1(n518), .CO(n51953));
    SB_LUT4 add_6061_10_lut (.I0(GND_net), .I1(n14058[7]), .I2(n664_adj_4498), 
            .I3(n50994), .O(n13134[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_21 (.CI(n50474), .I0(GND_net), .I1(n51[19]), 
            .CO(n50475));
    SB_LUT4 unary_minus_14_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n51[18]), 
            .I3(n50473), .O(n49[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6373_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_4497), .CO(n51782));
    SB_LUT4 add_6395_12_lut (.I0(GND_net), .I1(n19469[9]), .I2(n840), 
            .I3(n51781), .O(n19231[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_7_lut (.I0(GND_net), .I1(n14539[4]), .I2(n445_adj_4500), 
            .I3(n51951), .O(n13661[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6395_11_lut (.I0(GND_net), .I1(n19469[8]), .I2(n767), 
            .I3(n51780), .O(n19231[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_10 (.CI(n50994), .I0(n14058[7]), .I1(n664_adj_4498), 
            .CO(n50995));
    SB_LUT4 add_6061_9_lut (.I0(GND_net), .I1(n14058[6]), .I2(n591_adj_4501), 
            .I3(n50993), .O(n13134[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_9 (.CI(n50993), .I0(n14058[6]), .I1(n591_adj_4501), 
            .CO(n50994));
    SB_CARRY unary_minus_14_add_3_20 (.CI(n50473), .I0(GND_net), .I1(n51[18]), 
            .CO(n50474));
    SB_LUT4 unary_minus_14_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n51[17]), 
            .I3(n50472), .O(n49[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i17_4_lut (.I0(setpoint[16]), .I1(n483[16]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[16]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i17_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i22390_3_lut (.I0(n353[17]), .I1(n433[17]), .I2(n432), .I3(GND_net), 
            .O(n1_adj_4503));
    defparam i22390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i200_2_lut (.I0(\Ki[4] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6061_8_lut (.I0(GND_net), .I1(n14058[5]), .I2(n518_adj_4504), 
            .I3(n50992), .O(n13134[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_8 (.CI(n50992), .I0(n14058[5]), .I1(n518_adj_4504), 
            .CO(n50993));
    SB_CARRY add_6085_7 (.CI(n51951), .I0(n14539[4]), .I1(n445_adj_4500), 
            .CO(n51952));
    SB_LUT4 add_6085_6_lut (.I0(GND_net), .I1(n14539[3]), .I2(n372_adj_4505), 
            .I3(n51950), .O(n13661[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6061_7_lut (.I0(GND_net), .I1(n14058[4]), .I2(n445_adj_4506), 
            .I3(n50991), .O(n13134[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_19 (.CI(n50472), .I0(GND_net), .I1(n51[17]), 
            .CO(n50473));
    SB_LUT4 mult_17_i377_2_lut (.I0(\Kp[7] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_10_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n105[11]), .I3(n50369), .O(n48[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_7 (.CI(n50991), .I0(n14058[4]), .I1(n445_adj_4506), 
            .CO(n50992));
    SB_CARRY add_6085_6 (.CI(n51950), .I0(n14539[3]), .I1(n372_adj_4505), 
            .CO(n51951));
    SB_LUT4 add_6085_5_lut (.I0(GND_net), .I1(n14539[2]), .I2(n299_adj_4507), 
            .I3(n51949), .O(n13661[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6395_11 (.CI(n51780), .I0(n19469[8]), .I1(n767), .CO(n51781));
    SB_LUT4 add_6061_6_lut (.I0(GND_net), .I1(n14058[3]), .I2(n372_adj_4508), 
            .I3(n50990), .O(n13134[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_6 (.CI(n50990), .I0(n14058[3]), .I1(n372_adj_4508), 
            .CO(n50991));
    SB_LUT4 i22392_3_lut (.I0(n1_adj_4503), .I1(PWMLimit[17]), .I2(n406), 
            .I3(GND_net), .O(n3_adj_4509));
    defparam i22392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_4_lut (.I0(setpoint[17]), .I1(n3_adj_4509), 
            .I2(n15), .I3(n405), .O(duty_23__N_3602[17]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i18_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_6061_5_lut (.I0(GND_net), .I1(n14058[2]), .I2(n299_adj_4510), 
            .I3(n50989), .O(n13134[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6061_5 (.CI(n50989), .I0(n14058[2]), .I1(n299_adj_4510), 
            .CO(n50990));
    SB_LUT4 mux_28_i19_3_lut (.I0(n353[18]), .I1(n433[18]), .I2(n432), 
            .I3(GND_net), .O(n458[18]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i19_3_lut (.I0(n458[18]), .I1(PWMLimit[18]), .I2(n406), 
            .I3(GND_net), .O(n483[18]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6061_4_lut (.I0(GND_net), .I1(n14058[1]), .I2(n226_adj_4511), 
            .I3(n50988), .O(n13134[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i19_4_lut (.I0(setpoint[18]), .I1(n483[18]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[18]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i19_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mult_18_i549_2_lut (.I0(\Ki[11] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23371_3_lut (.I0(n353[19]), .I1(n433[19]), .I2(n432), .I3(GND_net), 
            .O(n1_adj_4512));
    defparam i23371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23373_3_lut (.I0(n1_adj_4512), .I1(PWMLimit[19]), .I2(n406), 
            .I3(GND_net), .O(n3_adj_4513));
    defparam i23373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_14_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n51[16]), 
            .I3(n50471), .O(n49[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_18 (.CI(n50471), .I0(GND_net), .I1(n51[16]), 
            .CO(n50472));
    SB_LUT4 unary_minus_14_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n51[15]), 
            .I3(n50470), .O(n49[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_17 (.CI(n50470), .I0(GND_net), .I1(n51[15]), 
            .CO(n50471));
    SB_CARRY add_6061_4 (.CI(n50988), .I0(n14058[1]), .I1(n226_adj_4511), 
            .CO(n50989));
    SB_LUT4 add_6061_3_lut (.I0(GND_net), .I1(n14058[0]), .I2(n153), .I3(n50987), 
            .O(n13134[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n51[14]), 
            .I3(n50469), .O(n49[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_9 (.CI(n50369), .I0(\PID_CONTROLLER.integral [7]), .I1(n105[11]), 
            .CO(n50370));
    SB_LUT4 add_6359_13_lut (.I0(GND_net), .I1(n19065[10]), .I2(n910_adj_4517), 
            .I3(n50593), .O(n18754[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_12_lut (.I0(GND_net), .I1(n19065[9]), .I2(n837_adj_4518), 
            .I3(n50592), .O(n18754[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_12 (.CI(n50592), .I0(n19065[9]), .I1(n837_adj_4518), 
            .CO(n50593));
    SB_LUT4 add_6359_11_lut (.I0(GND_net), .I1(n19065[8]), .I2(n764_adj_4519), 
            .I3(n50591), .O(n18754[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6395_10_lut (.I0(GND_net), .I1(n19469[7]), .I2(n694), 
            .I3(n51779), .O(n19231[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23374_4_lut (.I0(setpoint[19]), .I1(n3_adj_4513), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[19]));
    defparam i23374_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_28_i21_3_lut (.I0(n353[20]), .I1(n433[20]), .I2(n432), 
            .I3(GND_net), .O(n458[20]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Kp[3] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4439));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_29_i21_3_lut (.I0(n458[20]), .I1(PWMLimit[20]), .I2(n406), 
            .I3(GND_net), .O(n483[20]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_4_lut (.I0(setpoint[20]), .I1(n483[20]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[20]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i21_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY add_6061_3 (.CI(n50987), .I0(n14058[0]), .I1(n153), .CO(n50988));
    SB_CARRY add_6085_5 (.CI(n51949), .I0(n14539[2]), .I1(n299_adj_4507), 
            .CO(n51950));
    SB_LUT4 add_6467_7_lut (.I0(GND_net), .I1(n60191), .I2(n490_adj_4521), 
            .I3(n51312), .O(n19980[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6061_2_lut (.I0(GND_net), .I1(n11_adj_4522), .I2(n80), 
            .I3(GND_net), .O(n13134[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6061_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_4_lut (.I0(GND_net), .I1(n14539[1]), .I2(n226_adj_4523), 
            .I3(n51948), .O(n13661[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6467_6_lut (.I0(GND_net), .I1(n20063[3]), .I2(n417_adj_4524), 
            .I3(n51311), .O(n19980[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_6 (.CI(n51311), .I0(n20063[3]), .I1(n417_adj_4524), 
            .CO(n51312));
    SB_CARRY add_6085_4 (.CI(n51948), .I0(n14539[1]), .I1(n226_adj_4523), 
            .CO(n51949));
    SB_CARRY add_6061_2 (.CI(GND_net), .I0(n11_adj_4522), .I1(n80), .CO(n50987));
    SB_LUT4 add_6085_3_lut (.I0(GND_net), .I1(n14539[0]), .I2(n153_adj_4525), 
            .I3(n51947), .O(n13661[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6085_3 (.CI(n51947), .I0(n14539[0]), .I1(n153_adj_4525), 
            .CO(n51948));
    SB_CARRY add_6395_10 (.CI(n51779), .I0(n19469[7]), .I1(n694), .CO(n51780));
    SB_CARRY add_6359_11 (.CI(n50591), .I0(n19065[8]), .I1(n764_adj_4519), 
            .CO(n50592));
    SB_LUT4 add_6395_9_lut (.I0(GND_net), .I1(n19469[6]), .I2(n621), .I3(n51778), 
            .O(n19231[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6085_2_lut (.I0(GND_net), .I1(n11_adj_4526), .I2(n80_adj_4527), 
            .I3(GND_net), .O(n13661[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6085_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i22_3_lut (.I0(n353[21]), .I1(n433[21]), .I2(n432), 
            .I3(GND_net), .O(n458[21]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6085_2 (.CI(GND_net), .I0(n11_adj_4526), .I1(n80_adj_4527), 
            .CO(n51947));
    SB_LUT4 mux_29_i22_3_lut (.I0(n458[21]), .I1(PWMLimit[21]), .I2(n406), 
            .I3(GND_net), .O(n483[21]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6359_10_lut (.I0(GND_net), .I1(n19065[7]), .I2(n691_adj_4528), 
            .I3(n50590), .O(n18754[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_10 (.CI(n50590), .I0(n19065[7]), .I1(n691_adj_4528), 
            .CO(n50591));
    SB_LUT4 add_6359_9_lut (.I0(GND_net), .I1(n19065[6]), .I2(n618_adj_4529), 
            .I3(n50589), .O(n18754[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_16 (.CI(n50469), .I0(GND_net), .I1(n51[14]), 
            .CO(n50470));
    SB_LUT4 add_10_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n105[10]), .I3(n50368), .O(n48[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n51[13]), 
            .I3(n50468), .O(n49[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i22_4_lut (.I0(setpoint[21]), .I1(n483[21]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[21]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i22_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_6125_21_lut (.I0(GND_net), .I1(n15335[18]), .I2(GND_net), 
            .I3(n51946), .O(n14539[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6395_9 (.CI(n51778), .I0(n19469[6]), .I1(n621), .CO(n51779));
    SB_LUT4 add_6395_8_lut (.I0(GND_net), .I1(n19469[5]), .I2(n548), .I3(n51777), 
            .O(n19231[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_28_i23_3_lut (.I0(n353[22]), .I1(n433[22]), .I2(n432), 
            .I3(GND_net), .O(n458[22]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i23_3_lut (.I0(n458[22]), .I1(PWMLimit[22]), .I2(n406), 
            .I3(GND_net), .O(n483[22]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_4_lut (.I0(setpoint[22]), .I1(n483[22]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[22]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i23_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mux_28_i24_3_lut (.I0(n353[23]), .I1(n433[23]), .I2(n432), 
            .I3(GND_net), .O(n458[23]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i24_3_lut (.I0(n458[23]), .I1(PWMLimit[23]), .I2(n406), 
            .I3(GND_net), .O(n483[23]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_4_lut (.I0(setpoint[23]), .I1(n483[23]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[23]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i24_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_6467_5_lut (.I0(GND_net), .I1(n20063[2]), .I2(n344_adj_4532), 
            .I3(n51310), .O(n19980[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Kp[10] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4533));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6278_16_lut (.I0(GND_net), .I1(n17972[13]), .I2(n1120), 
            .I3(n50763), .O(n17493[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6395_8 (.CI(n51777), .I0(n19469[5]), .I1(n548), .CO(n51778));
    SB_LUT4 add_6278_15_lut (.I0(GND_net), .I1(n17972[12]), .I2(n1047), 
            .I3(n50762), .O(n17493[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6125_20_lut (.I0(GND_net), .I1(n15335[17]), .I2(GND_net), 
            .I3(n51945), .O(n14539[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6395_7_lut (.I0(GND_net), .I1(n19469[4]), .I2(n475_adj_4534), 
            .I3(n51776), .O(n19231[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6395_7 (.CI(n51776), .I0(n19469[4]), .I1(n475_adj_4534), 
            .CO(n51777));
    SB_CARRY add_6467_5 (.CI(n51310), .I0(n20063[2]), .I1(n344_adj_4532), 
            .CO(n51311));
    SB_LUT4 add_6395_6_lut (.I0(GND_net), .I1(n19469[3]), .I2(n402_adj_4535), 
            .I3(n51775), .O(n19231[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[2]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6395_6 (.CI(n51775), .I0(n19469[3]), .I1(n402_adj_4535), 
            .CO(n51776));
    SB_CARRY unary_minus_14_add_3_15 (.CI(n50468), .I0(GND_net), .I1(n51[13]), 
            .CO(n50469));
    SB_LUT4 add_6467_4_lut (.I0(GND_net), .I1(n20063[1]), .I2(n271_adj_4537), 
            .I3(n51309), .O(n19980[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_8 (.CI(n50368), .I0(\PID_CONTROLLER.integral [6]), .I1(n105[10]), 
            .CO(n50369));
    SB_CARRY add_6359_9 (.CI(n50589), .I0(n19065[6]), .I1(n618_adj_4529), 
            .CO(n50590));
    SB_LUT4 add_10_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n105[9]), .I3(n50367), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_15 (.CI(n50762), .I0(n17972[12]), .I1(n1047), .CO(n50763));
    SB_LUT4 mult_18_i598_2_lut (.I0(\Ki[12] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6125_20 (.CI(n51945), .I0(n15335[17]), .I1(GND_net), 
            .CO(n51946));
    SB_LUT4 add_6395_5_lut (.I0(GND_net), .I1(n19469[2]), .I2(n329), .I3(n51774), 
            .O(n19231[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6395_5 (.CI(n51774), .I0(n19469[2]), .I1(n329), .CO(n51775));
    SB_LUT4 unary_minus_14_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n51[12]), 
            .I3(n50467), .O(n49[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_4 (.CI(n51309), .I0(n20063[1]), .I1(n271_adj_4537), 
            .CO(n51310));
    SB_LUT4 add_6467_3_lut (.I0(GND_net), .I1(n20063[0]), .I2(n198_adj_4540), 
            .I3(n51308), .O(n19980[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6467_3 (.CI(n51308), .I0(n20063[0]), .I1(n198_adj_4540), 
            .CO(n51309));
    SB_LUT4 add_6125_19_lut (.I0(GND_net), .I1(n15335[16]), .I2(GND_net), 
            .I3(n51944), .O(n14539[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6395_4_lut (.I0(GND_net), .I1(n19469[1]), .I2(n256_adj_4541), 
            .I3(n51773), .O(n19231[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_19 (.CI(n51944), .I0(n15335[16]), .I1(GND_net), 
            .CO(n51945));
    SB_LUT4 add_6125_18_lut (.I0(GND_net), .I1(n15335[15]), .I2(GND_net), 
            .I3(n51943), .O(n14539[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i249_2_lut (.I0(\Ki[5] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6278_14_lut (.I0(GND_net), .I1(n17972[11]), .I2(n974), 
            .I3(n50761), .O(n17493[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_14 (.CI(n50761), .I0(n17972[11]), .I1(n974), .CO(n50762));
    SB_LUT4 add_6359_8_lut (.I0(GND_net), .I1(n19065[5]), .I2(n545_adj_4542), 
            .I3(n50588), .O(n18754[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_8 (.CI(n50588), .I0(n19065[5]), .I1(n545_adj_4542), 
            .CO(n50589));
    SB_LUT4 add_6359_7_lut (.I0(GND_net), .I1(n19065[4]), .I2(n472_adj_4543), 
            .I3(n50587), .O(n18754[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6467_2_lut (.I0(GND_net), .I1(n56_c), .I2(n125_adj_4544), 
            .I3(GND_net), .O(n19980[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6467_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6278_13_lut (.I0(GND_net), .I1(n17972[10]), .I2(n901), 
            .I3(n50760), .O(n17493[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_7 (.CI(n50367), .I0(\PID_CONTROLLER.integral [5]), .I1(n105[9]), 
            .CO(n50368));
    SB_CARRY add_6467_2 (.CI(GND_net), .I0(n56_c), .I1(n125_adj_4544), 
            .CO(n51308));
    SB_CARRY add_6278_13 (.CI(n50760), .I0(n17972[10]), .I1(n901), .CO(n50761));
    SB_LUT4 add_6278_12_lut (.I0(GND_net), .I1(n17972[9]), .I2(n828), 
            .I3(n50759), .O(n17493[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_7 (.CI(n50587), .I0(n19065[4]), .I1(n472_adj_4543), 
            .CO(n50588));
    SB_LUT4 add_6359_6_lut (.I0(GND_net), .I1(n19065[3]), .I2(n399_adj_4545), 
            .I3(n50586), .O(n18754[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_6 (.CI(n50586), .I0(n19065[3]), .I1(n399_adj_4545), 
            .CO(n50587));
    SB_LUT4 add_10_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n105[8]), .I3(n50366), .O(n48[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_18 (.CI(n51943), .I0(n15335[15]), .I1(GND_net), 
            .CO(n51944));
    SB_CARRY add_6278_12 (.CI(n50759), .I0(n17972[9]), .I1(n828), .CO(n50760));
    SB_LUT4 add_6278_11_lut (.I0(GND_net), .I1(n17972[8]), .I2(n755), 
            .I3(n50758), .O(n17493[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6125_17_lut (.I0(GND_net), .I1(n15335[14]), .I2(GND_net), 
            .I3(n51942), .O(n14539[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_5_lut (.I0(GND_net), .I1(n19065[2]), .I2(n326_adj_4546), 
            .I3(n50585), .O(n18754[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_17 (.CI(n51942), .I0(n15335[14]), .I1(GND_net), 
            .CO(n51943));
    SB_LUT4 add_6125_16_lut (.I0(GND_net), .I1(n15335[13]), .I2(n1105_adj_4547), 
            .I3(n51941), .O(n14539[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_16 (.CI(n51941), .I0(n15335[13]), .I1(n1105_adj_4547), 
            .CO(n51942));
    SB_CARRY add_6359_5 (.CI(n50585), .I0(n19065[2]), .I1(n326_adj_4546), 
            .CO(n50586));
    SB_LUT4 mult_18_i506_2_lut (.I0(\Ki[10] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4548));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i555_2_lut (.I0(\Ki[11] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4549));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Kp[15] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Kp[11] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4550));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i12_3_lut (.I0(n48[11]), .I1(n49[11]), .I2(n182), .I3(GND_net), 
            .O(n208[11]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i12_3_lut (.I0(n208[11]), .I1(IntegralLimit[11]), .I2(n156), 
            .I3(GND_net), .O(n233[11]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6278_11 (.CI(n50758), .I0(n17972[8]), .I1(n755), .CO(n50759));
    SB_LUT4 mult_18_i71_2_lut (.I0(\Ki[1] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i24_2_lut (.I0(\Ki[0] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i298_2_lut (.I0(\Ki[6] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i347_2_lut (.I0(\Ki[7] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i120_2_lut (.I0(\Ki[2] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Kp[4] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i647_2_lut (.I0(\Ki[13] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i169_2_lut (.I0(\Ki[3] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4436));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i696_2_lut (.I0(\Ki[14] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6125_15_lut (.I0(GND_net), .I1(n15335[12]), .I2(n1032_adj_4552), 
            .I3(n51940), .O(n14539[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6278_10_lut (.I0(GND_net), .I1(n17972[7]), .I2(n682), 
            .I3(n50757), .O(n17493[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_15 (.CI(n51940), .I0(n15335[12]), .I1(n1032_adj_4552), 
            .CO(n51941));
    SB_CARRY add_6395_4 (.CI(n51773), .I0(n19469[1]), .I1(n256_adj_4541), 
            .CO(n51774));
    SB_CARRY add_6278_10 (.CI(n50757), .I0(n17972[7]), .I1(n682), .CO(n50758));
    SB_LUT4 mult_17_i598_2_lut (.I0(\Kp[12] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4553));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6278_9_lut (.I0(GND_net), .I1(n17972[6]), .I2(n609), .I3(n50756), 
            .O(n17493[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Kp[13] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4554));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Kp[14] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4555));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6395_3_lut (.I0(GND_net), .I1(n19469[0]), .I2(n183), .I3(n51772), 
            .O(n19231[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_9 (.CI(n50756), .I0(n17972[6]), .I1(n609), .CO(n50757));
    SB_LUT4 add_6278_8_lut (.I0(GND_net), .I1(n17972[5]), .I2(n536), .I3(n50755), 
            .O(n17493[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_8 (.CI(n50755), .I0(n17972[5]), .I1(n536), .CO(n50756));
    SB_LUT4 add_6125_14_lut (.I0(GND_net), .I1(n15335[11]), .I2(n959_adj_4556), 
            .I3(n51939), .O(n14539[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6278_7_lut (.I0(GND_net), .I1(n17972[4]), .I2(n463), .I3(n50754), 
            .O(n17493[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i745_2_lut (.I0(\Ki[15] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6395_3 (.CI(n51772), .I0(n19469[0]), .I1(n183), .CO(n51773));
    SB_LUT4 mult_18_i218_2_lut (.I0(\Ki[4] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6125_14 (.CI(n51939), .I0(n15335[11]), .I1(n959_adj_4556), 
            .CO(n51940));
    SB_LUT4 add_6125_13_lut (.I0(GND_net), .I1(n15335[10]), .I2(n886_adj_4557), 
            .I3(n51938), .O(n14539[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_13 (.CI(n51938), .I0(n15335[10]), .I1(n886_adj_4557), 
            .CO(n51939));
    SB_LUT4 add_6125_12_lut (.I0(GND_net), .I1(n15335[9]), .I2(n813_adj_4558), 
            .I3(n51937), .O(n14539[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_4_lut (.I0(GND_net), .I1(n19065[1]), .I2(n253_adj_4559), 
            .I3(n50584), .O(n18754[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6395_2_lut (.I0(GND_net), .I1(n41), .I2(n110_adj_4560), 
            .I3(GND_net), .O(n19231[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6395_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_12 (.CI(n51937), .I0(n15335[9]), .I1(n813_adj_4558), 
            .CO(n51938));
    SB_LUT4 LessThan_20_i41_2_lut (.I0(deadband[20]), .I1(n353[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4561));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Kp[15] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4562));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[3]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_20_i39_2_lut (.I0(deadband[19]), .I1(n353[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i45_2_lut (.I0(deadband[22]), .I1(n353[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i37_2_lut (.I0(deadband[18]), .I1(n353[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_14_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[4]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6278_7 (.CI(n50754), .I0(n17972[4]), .I1(n463), .CO(n50755));
    SB_LUT4 unary_minus_14_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[5]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6395_2 (.CI(GND_net), .I0(n41), .I1(n110_adj_4560), .CO(n51772));
    SB_LUT4 unary_minus_14_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[6]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_20_i43_2_lut (.I0(deadband[21]), .I1(n353[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6278_6_lut (.I0(GND_net), .I1(n17972[3]), .I2(n390_adj_4567), 
            .I3(n50753), .O(n17493[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_4 (.CI(n50584), .I0(n19065[1]), .I1(n253_adj_4559), 
            .CO(n50585));
    SB_LUT4 LessThan_20_i21_2_lut (.I0(deadband[10]), .I1(n353[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4568));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6278_6 (.CI(n50753), .I0(n17972[3]), .I1(n390_adj_4567), 
            .CO(n50754));
    SB_LUT4 add_6278_5_lut (.I0(GND_net), .I1(n17972[2]), .I2(n317), .I3(n50752), 
            .O(n17493[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i23_2_lut (.I0(deadband[11]), .I1(n353[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4569));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6359_3_lut (.I0(GND_net), .I1(n19065[0]), .I2(n180_adj_4570), 
            .I3(n50583), .O(n18754[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_14 (.CI(n50467), .I0(GND_net), .I1(n51[12]), 
            .CO(n50468));
    SB_LUT4 unary_minus_14_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n51[11]), 
            .I3(n50466), .O(n49[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_5 (.CI(n50752), .I0(n17972[2]), .I1(n317), .CO(n50753));
    SB_CARRY add_6359_3 (.CI(n50583), .I0(n19065[0]), .I1(n180_adj_4570), 
            .CO(n50584));
    SB_CARRY add_10_6 (.CI(n50366), .I0(\PID_CONTROLLER.integral [4]), .I1(n105[8]), 
            .CO(n50367));
    SB_LUT4 add_6278_4_lut (.I0(GND_net), .I1(n17972[1]), .I2(n244_c), 
            .I3(n50751), .O(n17493[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_4 (.CI(n50751), .I0(n17972[1]), .I1(n244_c), .CO(n50752));
    SB_LUT4 add_6278_3_lut (.I0(GND_net), .I1(n17972[0]), .I2(n171), .I3(n50750), 
            .O(n17493[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_13 (.CI(n50466), .I0(GND_net), .I1(n51[11]), 
            .CO(n50467));
    SB_LUT4 add_6125_11_lut (.I0(GND_net), .I1(n15335[8]), .I2(n740_adj_4572), 
            .I3(n51936), .O(n14539[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n51[10]), 
            .I3(n50465), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_12 (.CI(n50465), .I0(GND_net), .I1(n51[10]), 
            .CO(n50466));
    SB_LUT4 add_6359_2_lut (.I0(GND_net), .I1(n38_adj_4574), .I2(n107_adj_4575), 
            .I3(GND_net), .O(n18754[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n105[7]), .I3(n50365), .O(n48[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_3 (.CI(n50750), .I0(n17972[0]), .I1(n171), .CO(n50751));
    SB_LUT4 LessThan_20_i25_2_lut (.I0(deadband[12]), .I1(n353[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4576));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6125_11 (.CI(n51936), .I0(n15335[8]), .I1(n740_adj_4572), 
            .CO(n51937));
    SB_CARRY add_6359_2 (.CI(GND_net), .I0(n38_adj_4574), .I1(n107_adj_4575), 
            .CO(n50583));
    SB_LUT4 add_6278_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n17493[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6278_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6278_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n50750));
    SB_LUT4 unary_minus_14_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n51[9]), 
            .I3(n50464), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_11 (.CI(n50464), .I0(GND_net), .I1(n51[9]), 
            .CO(n50465));
    SB_CARRY add_10_5 (.CI(n50365), .I0(\PID_CONTROLLER.integral [3]), .I1(n105[7]), 
            .CO(n50366));
    SB_LUT4 unary_minus_14_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n51[8]), 
            .I3(n50463), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i29_2_lut (.I0(deadband[14]), .I1(n353[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4580));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i31_2_lut (.I0(deadband[15]), .I1(n353[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(deadband[8]), .I1(n353[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4581));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6125_10_lut (.I0(GND_net), .I1(n15335[7]), .I2(n667_adj_4582), 
            .I3(n51935), .O(n14539[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_10 (.CI(n51935), .I0(n15335[7]), .I1(n667_adj_4582), 
            .CO(n51936));
    SB_LUT4 add_6125_9_lut (.I0(GND_net), .I1(n15335[6]), .I2(n594_adj_4583), 
            .I3(n51934), .O(n14539[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[7]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_14_add_3_10 (.CI(n50463), .I0(GND_net), .I1(n51[8]), 
            .CO(n50464));
    SB_LUT4 add_10_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n105[6]), .I3(n50364), .O(n48[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(deadband[9]), .I1(n353[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4586));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(deadband[4]), .I1(n353[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4587));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_2_lut (.I0(deadband[17]), .I1(n353[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4588));
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i11_2_lut (.I0(deadband[5]), .I1(n353[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4589));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_18_i604_2_lut (.I0(\Ki[12] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4590));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6125_9 (.CI(n51934), .I0(n15335[6]), .I1(n594_adj_4583), 
            .CO(n51935));
    SB_LUT4 add_6125_8_lut (.I0(GND_net), .I1(n15335[5]), .I2(n521_adj_4591), 
            .I3(n51933), .O(n14539[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_8 (.CI(n51933), .I0(n15335[5]), .I1(n521_adj_4591), 
            .CO(n51934));
    SB_LUT4 add_6125_7_lut (.I0(GND_net), .I1(n15335[4]), .I2(n448_adj_4592), 
            .I3(n51932), .O(n14539[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_7 (.CI(n51932), .I0(n15335[4]), .I1(n448_adj_4592), 
            .CO(n51933));
    SB_LUT4 add_6125_6_lut (.I0(GND_net), .I1(n15335[3]), .I2(n375_adj_4593), 
            .I3(n51931), .O(n14539[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_6 (.CI(n51931), .I0(n15335[3]), .I1(n375_adj_4593), 
            .CO(n51932));
    SB_LUT4 LessThan_20_i13_2_lut (.I0(deadband[6]), .I1(n353[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4594));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_15_i5_3_lut (.I0(n48[4]), .I1(n49[4]), .I2(n182), .I3(GND_net), 
            .O(n208[4]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(deadband[7]), .I1(n353[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4595));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i27_2_lut (.I0(deadband[13]), .I1(n353[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i33_2_lut (.I0(deadband[16]), .I1(n353[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51592_4_lut (.I0(n353[6]), .I1(n353[5]), .I2(n379[6]), .I3(n379[5]), 
            .O(n67318));
    defparam i51592_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 add_6125_5_lut (.I0(GND_net), .I1(n15335[2]), .I2(n302_adj_4596), 
            .I3(n51930), .O(n14539[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_5 (.CI(n51930), .I0(n15335[2]), .I1(n302_adj_4596), 
            .CO(n51931));
    SB_LUT4 add_6125_4_lut (.I0(GND_net), .I1(n15335[1]), .I2(n229_adj_4597), 
            .I3(n51929), .O(n14539[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_4 (.CI(n51929), .I0(n15335[1]), .I1(n229_adj_4597), 
            .CO(n51930));
    SB_LUT4 i52432_3_lut (.I0(n353[7]), .I1(n67318), .I2(n379[7]), .I3(GND_net), 
            .O(n68158));
    defparam i52432_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_22_i27_rep_167_2_lut (.I0(n353[13]), .I1(n379[13]), 
            .I2(GND_net), .I3(GND_net), .O(n70652));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i27_rep_167_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6125_3_lut (.I0(GND_net), .I1(n15335[0]), .I2(n156_adj_4598), 
            .I3(n51928), .O(n14539[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_3 (.CI(n51928), .I0(n15335[0]), .I1(n156_adj_4598), 
            .CO(n51929));
    SB_LUT4 add_6125_2_lut (.I0(GND_net), .I1(n14_adj_4599), .I2(n83_adj_4600), 
            .I3(GND_net), .O(n14539[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6125_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6125_2 (.CI(GND_net), .I0(n14_adj_4599), .I1(n83_adj_4600), 
            .CO(n51928));
    SB_LUT4 add_6163_20_lut (.I0(GND_net), .I1(n16053[17]), .I2(GND_net), 
            .I3(n51927), .O(n15335[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_19_lut (.I0(GND_net), .I1(n16053[16]), .I2(GND_net), 
            .I3(n51926), .O(n15335[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_19 (.CI(n51926), .I0(n16053[16]), .I1(GND_net), 
            .CO(n51927));
    SB_LUT4 i52414_4_lut (.I0(n353[14]), .I1(n70652), .I2(n379[14]), .I3(n68158), 
            .O(n68140));
    defparam i52414_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_22_i31_rep_162_2_lut (.I0(n353[15]), .I1(n379[15]), 
            .I2(GND_net), .I3(GND_net), .O(n70647));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i31_rep_162_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51582_4_lut (.I0(n353[8]), .I1(n353[4]), .I2(n379[8]), .I3(n379[4]), 
            .O(n67308));
    defparam i51582_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mux_16_i5_3_lut (.I0(n208[4]), .I1(IntegralLimit[4]), .I2(n156), 
            .I3(GND_net), .O(n233[4]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i653_2_lut (.I0(\Ki[13] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4601));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i57_2_lut (.I0(\Ki[1] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4600));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i10_2_lut (.I0(\Ki[0] ), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4599));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i106_2_lut (.I0(\Ki[2] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4598));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i155_2_lut (.I0(\Ki[3] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4597));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i204_2_lut (.I0(\Ki[4] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4596));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52426_3_lut (.I0(n353[9]), .I1(n67308), .I2(n379[9]), .I3(GND_net), 
            .O(n68152));
    defparam i52426_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 mult_18_i253_2_lut (.I0(\Ki[5] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4593));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6163_18_lut (.I0(GND_net), .I1(n16053[15]), .I2(GND_net), 
            .I3(n51925), .O(n15335[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_18 (.CI(n51925), .I0(n16053[15]), .I1(GND_net), 
            .CO(n51926));
    SB_LUT4 mult_18_i302_2_lut (.I0(\Ki[6] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4592));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i351_2_lut (.I0(\Ki[7] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4591));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i21_rep_182_2_lut (.I0(n353[10]), .I1(n379[10]), 
            .I2(GND_net), .I3(GND_net), .O(n70667));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i21_rep_182_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52420_4_lut (.I0(n353[11]), .I1(n70667), .I2(n379[11]), .I3(n68152), 
            .O(n68146));
    defparam i52420_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_22_i25_rep_177_2_lut (.I0(n353[12]), .I1(n379[12]), 
            .I2(GND_net), .I3(GND_net), .O(n70662));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i25_rep_177_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i16_3_lut (.I0(n379[9]), .I1(n379[21]), .I2(n353[21]), 
            .I3(GND_net), .O(n16_adj_4602));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51555_4_lut (.I0(n353[21]), .I1(n353[9]), .I2(n379[21]), 
            .I3(n379[9]), .O(n67281));
    defparam i51555_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_22_i8_3_lut (.I0(n379[4]), .I1(n379[8]), .I2(n353[8]), 
            .I3(GND_net), .O(n8_adj_4603));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_22_i24_3_lut (.I0(n16_adj_4602), .I1(n379[22]), .I2(n353[22]), 
            .I3(GND_net), .O(n24_adj_4604));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51603_4_lut (.I0(n353[3]), .I1(n353[2]), .I2(n379[3]), .I3(n379[2]), 
            .O(n67329));
    defparam i51603_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_22_i9_rep_175_2_lut (.I0(n353[4]), .I1(n379[4]), .I2(GND_net), 
            .I3(GND_net), .O(n70660));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i9_rep_175_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51600_4_lut (.I0(n353[5]), .I1(n70660), .I2(n379[5]), .I3(n67329), 
            .O(n67326));
    defparam i51600_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_22_i13_rep_203_2_lut (.I0(n353[6]), .I1(n379[6]), .I2(GND_net), 
            .I3(GND_net), .O(n70688));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i13_rep_203_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52787_4_lut (.I0(n353[7]), .I1(n70688), .I2(n379[7]), .I3(n67326), 
            .O(n68513));
    defparam i52787_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_18_i400_2_lut (.I0(\Ki[8] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4583));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6163_17_lut (.I0(GND_net), .I1(n16053[14]), .I2(GND_net), 
            .I3(n51924), .O(n15335[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i449_2_lut (.I0(\Ki[9] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4582));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n51[7]), 
            .I3(n50462), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_9 (.CI(n50462), .I0(GND_net), .I1(n51[7]), 
            .CO(n50463));
    SB_CARRY add_10_4 (.CI(n50364), .I0(\PID_CONTROLLER.integral [2]), .I1(n105[6]), 
            .CO(n50365));
    SB_CARRY add_6163_17 (.CI(n51924), .I0(n16053[14]), .I1(GND_net), 
            .CO(n51925));
    SB_LUT4 LessThan_22_i17_rep_200_2_lut (.I0(n353[8]), .I1(n379[8]), .I2(GND_net), 
            .I3(GND_net), .O(n70685));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i17_rep_200_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_14_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[8]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_14_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[9]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_14_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n51[6]), 
            .I3(n50461), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_8 (.CI(n50461), .I0(GND_net), .I1(n51[6]), 
            .CO(n50462));
    SB_LUT4 unary_minus_14_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n51[5]), 
            .I3(n50460), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_10_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n105[5]), .I3(n50363), .O(n48[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_7 (.CI(n50460), .I0(GND_net), .I1(n51[5]), 
            .CO(n50461));
    SB_LUT4 unary_minus_14_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n51[4]), 
            .I3(n50459), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_3 (.CI(n50363), .I0(\PID_CONTROLLER.integral [1]), .I1(n105[5]), 
            .CO(n50364));
    SB_CARRY unary_minus_14_add_3_6 (.CI(n50459), .I0(GND_net), .I1(n51[4]), 
            .CO(n50460));
    SB_LUT4 unary_minus_14_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n51[3]), 
            .I3(n50458), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_16_lut (.I0(GND_net), .I1(n16053[13]), .I2(n1108), 
            .I3(n51923), .O(n15335[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52430_4_lut (.I0(n353[9]), .I1(n70685), .I2(n379[9]), .I3(n68513), 
            .O(n68156));
    defparam i52430_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i53053_4_lut (.I0(n353[11]), .I1(n70667), .I2(n379[11]), .I3(n68156), 
            .O(n68779));
    defparam i53053_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i51574_4_lut (.I0(n353[13]), .I1(n70662), .I2(n379[13]), .I3(n68779), 
            .O(n67300));
    defparam i51574_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Kp[1] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_10_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n105[4]), .I3(GND_net), .O(n48[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_10_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Kp[0] ), .I1(n105[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Kp[1] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4575));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_14_add_3_5 (.CI(n50458), .I0(GND_net), .I1(n51[3]), 
            .CO(n50459));
    SB_LUT4 mult_17_i26_2_lut (.I0(\Kp[0] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4574));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[10]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6163_16 (.CI(n51923), .I0(n16053[13]), .I1(n1108), .CO(n51924));
    SB_LUT4 add_6163_15_lut (.I0(GND_net), .I1(n16053[12]), .I2(n1035), 
            .I3(n51922), .O(n15335[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_15 (.CI(n51922), .I0(n16053[12]), .I1(n1035), .CO(n51923));
    SB_LUT4 LessThan_22_i29_rep_166_2_lut (.I0(n353[14]), .I1(n379[14]), 
            .I2(GND_net), .I3(GND_net), .O(n70651));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i29_rep_166_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6163_14_lut (.I0(GND_net), .I1(n16053[11]), .I2(n962), 
            .I3(n51921), .O(n15335[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52781_4_lut (.I0(n353[15]), .I1(n70651), .I2(n379[15]), .I3(n67300), 
            .O(n68507));
    defparam i52781_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_22_i33_rep_192_2_lut (.I0(n353[16]), .I1(n379[16]), 
            .I2(GND_net), .I3(GND_net), .O(n70677));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i33_rep_192_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53292_4_lut (.I0(n353[17]), .I1(n70677), .I2(n379[17]), .I3(n68507), 
            .O(n69018));
    defparam i53292_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_6163_14 (.CI(n51921), .I0(n16053[11]), .I1(n962), .CO(n51922));
    SB_LUT4 add_6163_13_lut (.I0(GND_net), .I1(n16053[10]), .I2(n889), 
            .I3(n51920), .O(n15335[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_10_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n105[4]), .CO(n50363));
    SB_CARRY add_6163_13 (.CI(n51920), .I0(n16053[10]), .I1(n889), .CO(n51921));
    SB_LUT4 mult_18_i498_2_lut (.I0(\Ki[10] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4572));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n51[2]), 
            .I3(n50457), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_9_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n50362), .O(n105[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Kp[2] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6163_12_lut (.I0(GND_net), .I1(n16053[9]), .I2(n816), 
            .I3(n51919), .O(n15335[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i37_rep_156_2_lut (.I0(n353[18]), .I1(n379[18]), 
            .I2(GND_net), .I3(GND_net), .O(n70641));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i37_rep_156_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Kp[3] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[11]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53501_4_lut (.I0(n353[19]), .I1(n70641), .I2(n379[19]), .I3(n69018), 
            .O(n69227));
    defparam i53501_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY unary_minus_14_add_3_4 (.CI(n50457), .I0(GND_net), .I1(n51[2]), 
            .CO(n50458));
    SB_LUT4 sub_9_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n50361), .O(n105[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n51[1]), 
            .I3(n50456), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Kp[2] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4570));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6163_12 (.CI(n51919), .I0(n16053[9]), .I1(n816), .CO(n51920));
    SB_LUT4 mult_17_i214_2_lut (.I0(\Kp[4] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Kp[5] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4567));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_9_add_2_24 (.CI(n50361), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n50362));
    SB_LUT4 LessThan_22_i41_rep_153_2_lut (.I0(n353[20]), .I1(n379[20]), 
            .I2(GND_net), .I3(GND_net), .O(n70638));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i41_rep_153_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6103_21_lut (.I0(GND_net), .I1(n14897[18]), .I2(GND_net), 
            .I3(n50964), .O(n14058[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51629_4_lut (.I0(n27), .I1(n15_adj_4595), .I2(n13_adj_4594), 
            .I3(n11_adj_4589), .O(n67355));
    defparam i51629_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_15_i14_3_lut (.I0(n48[13]), .I1(n49[13]), .I2(n182), .I3(GND_net), 
            .O(n219));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i12_3_lut (.I0(n353[7]), .I1(n353[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4606));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i75_2_lut (.I0(\Ki[1] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4560));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i171_2_lut (.I0(\Kp[3] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4559));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6103_20_lut (.I0(GND_net), .I1(n14897[17]), .I2(GND_net), 
            .I3(n50963), .O(n14058[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_11_lut (.I0(GND_net), .I1(n16053[8]), .I2(n743), 
            .I3(n51918), .O(n15335[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i10_3_lut (.I0(n353[5]), .I1(n353[6]), .I2(n13_adj_4594), 
            .I3(GND_net), .O(n10_adj_4607));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6163_11 (.CI(n51918), .I0(n16053[8]), .I1(n743), .CO(n51919));
    SB_CARRY add_6103_20 (.CI(n50963), .I0(n14897[17]), .I1(GND_net), 
            .CO(n50964));
    SB_LUT4 LessThan_20_i30_3_lut (.I0(n12_adj_4606), .I1(n353[17]), .I2(n35_adj_4588), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52469_4_lut (.I0(n13_adj_4594), .I1(n11_adj_4589), .I2(n9_adj_4587), 
            .I3(n67418), .O(n68195));
    defparam i52469_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52465_4_lut (.I0(n19_adj_4586), .I1(n17_adj_4581), .I2(n15_adj_4595), 
            .I3(n68195), .O(n68191));
    defparam i52465_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53346_4_lut (.I0(n25_adj_4576), .I1(n23_adj_4569), .I2(n21_adj_4568), 
            .I3(n68191), .O(n69072));
    defparam i53346_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52797_4_lut (.I0(n31), .I1(n29_adj_4580), .I2(n27), .I3(n69072), 
            .O(n68523));
    defparam i52797_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53417_4_lut (.I0(n37), .I1(n35_adj_4588), .I2(n33), .I3(n68523), 
            .O(n69143));
    defparam i53417_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_20_i16_3_lut (.I0(n353[9]), .I1(n353[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4608));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n353[4]), .I1(n353[8]), .I2(n17_adj_4581), 
            .I3(GND_net), .O(n8_adj_4609));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i24_3_lut (.I0(n16_adj_4608), .I1(n353[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4610));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52929_3_lut (.I0(n6_adj_4611), .I1(n353[10]), .I2(n21_adj_4568), 
            .I3(GND_net), .O(n68655));   // verilog/motorControl.v(56[16:33])
    defparam i52929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52930_3_lut (.I0(n68655), .I1(n353[11]), .I2(n23_adj_4569), 
            .I3(GND_net), .O(n68656));   // verilog/motorControl.v(56[16:33])
    defparam i52930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51673_4_lut (.I0(n21_adj_4568), .I1(n19_adj_4586), .I2(n17_adj_4581), 
            .I3(n9_adj_4587), .O(n67399));
    defparam i51673_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51608_4_lut (.I0(n43), .I1(n25_adj_4576), .I2(n23_adj_4569), 
            .I3(n67399), .O(n67334));
    defparam i51608_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52563_4_lut (.I0(n24_adj_4610), .I1(n8_adj_4609), .I2(n45), 
            .I3(n67332), .O(n68289));   // verilog/motorControl.v(56[16:33])
    defparam i52563_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51873_3_lut (.I0(n68656), .I1(n353[12]), .I2(n25_adj_4576), 
            .I3(GND_net), .O(n67599));   // verilog/motorControl.v(56[16:33])
    defparam i51873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i4_3_lut (.I0(n66320), .I1(n379[1]), .I2(n353[1]), 
            .I3(GND_net), .O(n4_adj_4612));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52919_3_lut (.I0(n4_adj_4612), .I1(n379[13]), .I2(n353[13]), 
            .I3(GND_net), .O(n68645));   // verilog/motorControl.v(56[37:57])
    defparam i52919_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52920_3_lut (.I0(n68645), .I1(n379[14]), .I2(n353[14]), .I3(GND_net), 
            .O(n68646));   // verilog/motorControl.v(56[37:57])
    defparam i52920_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_22_i12_3_lut (.I0(n379[7]), .I1(n379[16]), .I2(n353[16]), 
            .I3(GND_net), .O(n12_adj_4613));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51566_4_lut (.I0(n353[16]), .I1(n353[7]), .I2(n379[16]), 
            .I3(n379[7]), .O(n67292));
    defparam i51566_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_22_i35_rep_188_2_lut (.I0(n353[17]), .I1(n379[17]), 
            .I2(GND_net), .I3(GND_net), .O(n70673));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i35_rep_188_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i10_3_lut (.I0(n379[5]), .I1(n379[6]), .I2(n353[6]), 
            .I3(GND_net), .O(n10_adj_4614));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_22_i30_3_lut (.I0(n12_adj_4613), .I1(n379[17]), .I2(n353[17]), 
            .I3(GND_net), .O(n30_adj_4615));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51568_4_lut (.I0(n353[16]), .I1(n70647), .I2(n379[16]), .I3(n68140), 
            .O(n67294));
    defparam i51568_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i53308_4_lut (.I0(n30_adj_4615), .I1(n10_adj_4614), .I2(n70673), 
            .I3(n67292), .O(n69034));   // verilog/motorControl.v(56[37:57])
    defparam i53308_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51885_3_lut (.I0(n68646), .I1(n379[15]), .I2(n353[15]), .I3(GND_net), 
            .O(n67611));   // verilog/motorControl.v(56[37:57])
    defparam i51885_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53488_4_lut (.I0(n67611), .I1(n69034), .I2(n70673), .I3(n67294), 
            .O(n69214));   // verilog/motorControl.v(56[37:57])
    defparam i53488_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53489_3_lut (.I0(n69214), .I1(n379[18]), .I2(n353[18]), .I3(GND_net), 
            .O(n69215));   // verilog/motorControl.v(56[37:57])
    defparam i53489_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53446_3_lut (.I0(n69215), .I1(n379[19]), .I2(n353[19]), .I3(GND_net), 
            .O(n69172));   // verilog/motorControl.v(56[37:57])
    defparam i53446_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_22_i6_3_lut (.I0(n379[2]), .I1(n379[3]), .I2(n353[3]), 
            .I3(GND_net), .O(n6_adj_4616));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52921_3_lut (.I0(n6_adj_4616), .I1(n379[10]), .I2(n353[10]), 
            .I3(GND_net), .O(n68647));   // verilog/motorControl.v(56[37:57])
    defparam i52921_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52922_3_lut (.I0(n68647), .I1(n379[11]), .I2(n353[11]), .I3(GND_net), 
            .O(n68648));   // verilog/motorControl.v(56[37:57])
    defparam i52922_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51557_4_lut (.I0(n353[21]), .I1(n70662), .I2(n379[21]), .I3(n68146), 
            .O(n67283));
    defparam i51557_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_18_i547_2_lut (.I0(\Ki[11] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4558));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52565_4_lut (.I0(n24_adj_4604), .I1(n8_adj_4603), .I2(n70636), 
            .I3(n67281), .O(n68291));   // verilog/motorControl.v(56[37:57])
    defparam i52565_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51883_3_lut (.I0(n68648), .I1(n379[12]), .I2(n353[12]), .I3(GND_net), 
            .O(n67609));   // verilog/motorControl.v(56[37:57])
    defparam i51883_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51559_4_lut (.I0(n353[21]), .I1(n70638), .I2(n379[21]), .I3(n69227), 
            .O(n67285));
    defparam i51559_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_22_i45_rep_151_2_lut (.I0(n353[22]), .I1(n379[22]), 
            .I2(GND_net), .I3(GND_net), .O(n70636));   // verilog/motorControl.v(56[37:57])
    defparam LessThan_22_i45_rep_151_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_18_i596_2_lut (.I0(\Ki[12] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4557));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53173_4_lut (.I0(n67609), .I1(n68291), .I2(n70636), .I3(n67283), 
            .O(n68899));   // verilog/motorControl.v(56[37:57])
    defparam i53173_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51891_3_lut (.I0(n69172), .I1(n379[20]), .I2(n353[20]), .I3(GND_net), 
            .O(n67617));   // verilog/motorControl.v(56[37:57])
    defparam i51891_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6103_19_lut (.I0(GND_net), .I1(n14897[16]), .I2(GND_net), 
            .I3(n50962), .O(n14058[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53364_4_lut (.I0(n67617), .I1(n68899), .I2(n70636), .I3(n67285), 
            .O(n69090));   // verilog/motorControl.v(56[37:57])
    defparam i53364_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6163_10_lut (.I0(GND_net), .I1(n16053[7]), .I2(n670_adj_4471), 
            .I3(n51917), .O(n15335[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Kp[6] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i645_2_lut (.I0(\Ki[13] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4556));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Kp[7] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i124_2_lut (.I0(\Ki[2] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Kp[8] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i4_4_lut (.I0(deadband[0]), .I1(n353[1]), .I2(deadband[1]), 
            .I3(n353[0]), .O(n4_adj_4617));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52927_3_lut (.I0(n4_adj_4617), .I1(n353[13]), .I2(n27), .I3(GND_net), 
            .O(n68653));   // verilog/motorControl.v(56[16:33])
    defparam i52927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52928_3_lut (.I0(n68653), .I1(n353[14]), .I2(n29_adj_4580), 
            .I3(GND_net), .O(n68654));   // verilog/motorControl.v(56[16:33])
    defparam i52928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51619_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4580), .I3(n67355), 
            .O(n67345));
    defparam i51619_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53374_4_lut (.I0(n30), .I1(n10_adj_4607), .I2(n35_adj_4588), 
            .I3(n67342), .O(n69100));   // verilog/motorControl.v(56[16:33])
    defparam i53374_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51875_3_lut (.I0(n68654), .I1(n353[15]), .I2(n31), .I3(GND_net), 
            .O(n67601));   // verilog/motorControl.v(56[16:33])
    defparam i51875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53486_4_lut (.I0(n67601), .I1(n69100), .I2(n35_adj_4588), 
            .I3(n67345), .O(n69212));   // verilog/motorControl.v(56[16:33])
    defparam i53486_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53487_3_lut (.I0(n69212), .I1(n353[18]), .I2(n37), .I3(GND_net), 
            .O(n69213));   // verilog/motorControl.v(56[16:33])
    defparam i53487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53450_3_lut (.I0(n69213), .I1(n353[19]), .I2(n39), .I3(GND_net), 
            .O(n69176));   // verilog/motorControl.v(56[16:33])
    defparam i53450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51610_4_lut (.I0(n43), .I1(n41_adj_4561), .I2(n39), .I3(n69143), 
            .O(n67336));
    defparam i51610_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Kp[9] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i694_2_lut (.I0(\Ki[14] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4552));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6307_15_lut (.I0(GND_net), .I1(n18391[12]), .I2(n1050), 
            .I3(n50733), .O(n17972[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_14_lut (.I0(GND_net), .I1(n18391[11]), .I2(n977), 
            .I3(n50732), .O(n17972[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_3 (.CI(n50456), .I0(GND_net), .I1(n51[1]), 
            .CO(n50457));
    SB_CARRY add_6103_19 (.CI(n50962), .I0(n14897[16]), .I1(GND_net), 
            .CO(n50963));
    SB_CARRY add_6307_14 (.CI(n50732), .I0(n18391[11]), .I1(n977), .CO(n50733));
    SB_LUT4 add_6307_13_lut (.I0(GND_net), .I1(n18391[10]), .I2(n904), 
            .I3(n50731), .O(n17972[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n51[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_14_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_13 (.CI(n50731), .I0(n18391[10]), .I1(n904), .CO(n50732));
    SB_LUT4 i53171_4_lut (.I0(n67599), .I1(n68289), .I2(n45), .I3(n67334), 
            .O(n68897));   // verilog/motorControl.v(56[16:33])
    defparam i53171_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51881_3_lut (.I0(n69176), .I1(n353[20]), .I2(n41_adj_4561), 
            .I3(GND_net), .O(n67607));   // verilog/motorControl.v(56[16:33])
    defparam i51881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6103_18_lut (.I0(GND_net), .I1(n14897[15]), .I2(GND_net), 
            .I3(n50961), .O(n14058[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_12_lut (.I0(GND_net), .I1(n18391[9]), .I2(n831), 
            .I3(n50730), .O(n17972[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_10 (.CI(n51917), .I0(n16053[7]), .I1(n670_adj_4471), 
            .CO(n51918));
    SB_LUT4 add_6163_9_lut (.I0(GND_net), .I1(n16053[6]), .I2(n597_adj_4458), 
            .I3(n51916), .O(n15335[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_9 (.CI(n51916), .I0(n16053[6]), .I1(n597_adj_4458), 
            .CO(n51917));
    SB_CARRY add_6103_18 (.CI(n50961), .I0(n14897[15]), .I1(GND_net), 
            .CO(n50962));
    SB_CARRY add_6307_12 (.CI(n50730), .I0(n18391[9]), .I1(n831), .CO(n50731));
    SB_LUT4 add_6103_17_lut (.I0(GND_net), .I1(n14897[14]), .I2(GND_net), 
            .I3(n50960), .O(n14058[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_8_lut (.I0(GND_net), .I1(n16053[5]), .I2(n524_adj_4454), 
            .I3(n51915), .O(n15335[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_11_lut (.I0(GND_net), .I1(n18391[8]), .I2(n758), 
            .I3(n50729), .O(n17972[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_14_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n51[0]), 
            .CO(n50456));
    SB_LUT4 sub_9_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n50360), .O(n105[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_17 (.CI(n50960), .I0(n14897[14]), .I1(GND_net), 
            .CO(n50961));
    SB_LUT4 add_6103_16_lut (.I0(GND_net), .I1(n14897[13]), .I2(n1105), 
            .I3(n50959), .O(n14058[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_8 (.CI(n51915), .I0(n16053[5]), .I1(n524_adj_4454), 
            .CO(n51916));
    SB_CARRY add_6307_11 (.CI(n50729), .I0(n18391[8]), .I1(n758), .CO(n50730));
    SB_CARRY sub_9_add_2_23 (.CI(n50360), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n50361));
    SB_LUT4 i53365_3_lut (.I0(n69090), .I1(n353[23]), .I2(n47), .I3(GND_net), 
            .O(n69091));   // verilog/motorControl.v(56[37:57])
    defparam i53365_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6103_16 (.CI(n50959), .I0(n14897[13]), .I1(n1105), .CO(n50960));
    SB_LUT4 add_6307_10_lut (.I0(GND_net), .I1(n18391[7]), .I2(n685), 
            .I3(n50728), .O(n17972[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53362_4_lut (.I0(n67607), .I1(n68897), .I2(n45), .I3(n67336), 
            .O(n69088));   // verilog/motorControl.v(56[16:33])
    defparam i53362_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24_4_lut (.I0(n69088), .I1(n69091), .I2(deadband[23]), .I3(n353[23]), 
            .O(n405));   // verilog/motorControl.v(56[16:57])
    defparam i24_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Kp[8] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6307_10 (.CI(n50728), .I0(n18391[7]), .I1(n685), .CO(n50729));
    SB_LUT4 add_6103_15_lut (.I0(GND_net), .I1(n14897[12]), .I2(n1032), 
            .I3(n50958), .O(n14058[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_9_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n50359), .O(n105[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_15 (.CI(n50958), .I0(n14897[12]), .I1(n1032), .CO(n50959));
    SB_LUT4 add_6307_9_lut (.I0(GND_net), .I1(n18391[6]), .I2(n612), .I3(n50727), 
            .O(n17972[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6103_14_lut (.I0(GND_net), .I1(n14897[11]), .I2(n959), 
            .I3(n50957), .O(n14058[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_9 (.CI(n50727), .I0(n18391[6]), .I1(n612), .CO(n50728));
    SB_LUT4 add_6307_8_lut (.I0(GND_net), .I1(n18391[5]), .I2(n539), .I3(n50726), 
            .O(n17972[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_8 (.CI(n50726), .I0(n18391[5]), .I1(n539), .CO(n50727));
    SB_LUT4 add_6307_7_lut (.I0(GND_net), .I1(n18391[4]), .I2(n466), .I3(n50725), 
            .O(n17972[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_22 (.CI(n50359), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n50360));
    SB_LUT4 add_6163_7_lut (.I0(GND_net), .I1(n16053[4]), .I2(n451_adj_4447), 
            .I3(n51914), .O(n15335[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_14 (.CI(n50957), .I0(n14897[11]), .I1(n959), .CO(n50958));
    SB_LUT4 mult_18_i743_2_lut (.I0(\Ki[15] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4547));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Kp[4] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4546));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_9_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n50358), .O(n105[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_7 (.CI(n50725), .I0(n18391[4]), .I1(n466), .CO(n50726));
    SB_LUT4 add_6307_6_lut (.I0(GND_net), .I1(n18391[3]), .I2(n393), .I3(n50724), 
            .O(n17972[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_7 (.CI(n51914), .I0(n16053[4]), .I1(n451_adj_4447), 
            .CO(n51915));
    SB_LUT4 mult_17_i508_2_lut (.I0(\Kp[10] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6103_13_lut (.I0(GND_net), .I1(n14897[10]), .I2(n886), 
            .I3(n50956), .O(n14058[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_13 (.CI(n50956), .I0(n14897[10]), .I1(n886), .CO(n50957));
    SB_LUT4 mult_17_i269_2_lut (.I0(\Kp[5] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4545));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Kp[11] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Kp[12] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i85_2_lut (.I0(\Kp[1] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4544));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i38_2_lut (.I0(\Kp[0] ), .I1(n105[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i38_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6307_6 (.CI(n50724), .I0(n18391[3]), .I1(n393), .CO(n50725));
    SB_LUT4 add_6307_5_lut (.I0(GND_net), .I1(n18391[2]), .I2(n320), .I3(n50723), 
            .O(n17972[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6103_12_lut (.I0(GND_net), .I1(n14897[9]), .I2(n813), 
            .I3(n50955), .O(n14058[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_5 (.CI(n50723), .I0(n18391[2]), .I1(n320), .CO(n50724));
    SB_CARRY add_6103_12 (.CI(n50955), .I0(n14897[9]), .I1(n813), .CO(n50956));
    SB_LUT4 add_6163_6_lut (.I0(GND_net), .I1(n16053[3]), .I2(n378), .I3(n51913), 
            .O(n15335[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_4_lut (.I0(GND_net), .I1(n18391[1]), .I2(n247), .I3(n50722), 
            .O(n17972[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_6 (.CI(n51913), .I0(n16053[3]), .I1(n378), .CO(n51914));
    SB_LUT4 add_6103_11_lut (.I0(GND_net), .I1(n14897[8]), .I2(n740), 
            .I3(n50954), .O(n14058[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_4 (.CI(n50722), .I0(n18391[1]), .I1(n247), .CO(n50723));
    SB_LUT4 add_6307_3_lut (.I0(GND_net), .I1(n18391[0]), .I2(n174), .I3(n50721), 
            .O(n17972[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i318_2_lut (.I0(\Kp[6] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4543));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Kp[7] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4542));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6163_5_lut (.I0(GND_net), .I1(n16053[2]), .I2(n305), .I3(n51912), 
            .O(n15335[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(IntegralLimit[4]), .I1(n48[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4618));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(IntegralLimit[6]), .I1(n48[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4619));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Kp[13] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i173_2_lut (.I0(\Ki[3] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4541));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(IntegralLimit[7]), .I1(n48[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4620));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_9_add_2_21 (.CI(n50358), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n50359));
    SB_CARRY add_6163_5 (.CI(n51912), .I0(n16053[2]), .I1(n305), .CO(n51913));
    SB_CARRY add_6307_3 (.CI(n50721), .I0(n18391[0]), .I1(n174), .CO(n50722));
    SB_LUT4 add_6307_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17972[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_11 (.CI(n50954), .I0(n14897[8]), .I1(n740), .CO(n50955));
    SB_LUT4 add_6103_10_lut (.I0(GND_net), .I1(n14897[7]), .I2(n667), 
            .I3(n50953), .O(n14058[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n50721));
    SB_LUT4 sub_9_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n50357), .O(n105[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_4_lut (.I0(GND_net), .I1(n16053[1]), .I2(n232), .I3(n51911), 
            .O(n15335[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i134_2_lut (.I0(\Kp[2] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4540));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[12]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i222_2_lut (.I0(\Ki[4] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(IntegralLimit[10]), .I1(n48[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4621));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6163_4 (.CI(n51911), .I0(n16053[1]), .I1(n232), .CO(n51912));
    SB_CARRY add_6103_10 (.CI(n50953), .I0(n14897[7]), .I1(n667), .CO(n50954));
    SB_LUT4 add_6475_7_lut (.I0(GND_net), .I1(n60827), .I2(n490), .I3(n50720), 
            .O(n20041[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_6_lut (.I0(GND_net), .I1(n20109[3]), .I2(n417), .I3(n50719), 
            .O(n20041[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(IntegralLimit[9]), .I1(n48[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4622));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(IntegralLimit[8]), .I1(n48[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4623));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6163_3_lut (.I0(GND_net), .I1(n16053[0]), .I2(n159), .I3(n51910), 
            .O(n15335[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6103_9_lut (.I0(GND_net), .I1(n14897[6]), .I2(n594), .I3(n50952), 
            .O(n14058[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_20 (.CI(n50357), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n50358));
    SB_CARRY add_6475_6 (.CI(n50719), .I0(n20109[3]), .I1(n417), .CO(n50720));
    SB_LUT4 sub_9_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n50356), .O(n105[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_9 (.CI(n50952), .I0(n14897[6]), .I1(n594), .CO(n50953));
    SB_LUT4 LessThan_13_i9_2_lut (.I0(n48[4]), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4624));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6163_3 (.CI(n51910), .I0(n16053[0]), .I1(n159), .CO(n51911));
    SB_LUT4 mult_17_i183_2_lut (.I0(\Kp[3] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4537));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_13_i11_2_lut (.I0(n150), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4625));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n105[23]), .I1(\Kp[2] ), .I2(n50049), 
            .I3(n105[22]), .O(n62910));   // verilog/motorControl.v(55[22:28])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'h6ca0;
    SB_LUT4 LessThan_13_i13_2_lut (.I0(n48[6]), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4626));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6475_5_lut (.I0(GND_net), .I1(n20112), .I2(n344), .I3(n50718), 
            .O(n20041[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_2_lut (.I0(GND_net), .I1(n17), .I2(n86), .I3(GND_net), 
            .O(n15335[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_2 (.CI(GND_net), .I0(n17), .I1(n86), .CO(n51910));
    SB_LUT4 LessThan_13_i15_2_lut (.I0(n48[7]), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4627));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6103_8_lut (.I0(GND_net), .I1(n14897[5]), .I2(n521), .I3(n50951), 
            .O(n14058[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_5 (.CI(n50718), .I0(n20112), .I1(n344), .CO(n50719));
    SB_CARRY add_6103_8 (.CI(n50951), .I0(n14897[5]), .I1(n521), .CO(n50952));
    SB_CARRY sub_9_add_2_19 (.CI(n50356), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n50357));
    SB_LUT4 add_6475_4_lut (.I0(GND_net), .I1(n20113), .I2(n271), .I3(n50717), 
            .O(n20041[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_4 (.CI(n50717), .I0(n20113), .I1(n271), .CO(n50718));
    SB_LUT4 add_6103_7_lut (.I0(GND_net), .I1(n14897[4]), .I2(n448), .I3(n50950), 
            .O(n14058[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_3_lut (.I0(GND_net), .I1(n20109[0]), .I2(n198), .I3(n50716), 
            .O(n20041[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_3 (.CI(n50716), .I0(n20109[0]), .I1(n198), .CO(n50717));
    SB_LUT4 sub_9_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(n7), 
            .I3(n50355), .O(n105[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_13_i21_2_lut (.I0(n48[10]), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4629));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6403_11_lut (.I0(GND_net), .I1(n19547[8]), .I2(n770), 
            .I3(n51909), .O(n19328[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_13_i19_2_lut (.I0(n48[9]), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4630));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6403_10_lut (.I0(GND_net), .I1(n19547[7]), .I2(n697), 
            .I3(n51908), .O(n19328[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6403_10 (.CI(n51908), .I0(n19547[7]), .I1(n697), .CO(n51909));
    SB_LUT4 add_6403_9_lut (.I0(GND_net), .I1(n19547[6]), .I2(n624_c), 
            .I3(n51907), .O(n19328[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i271_2_lut (.I0(\Ki[5] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4535));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6103_7 (.CI(n50950), .I0(n14897[4]), .I1(n448), .CO(n50951));
    SB_LUT4 add_6475_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20041[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n50716));
    SB_LUT4 add_6103_6_lut (.I0(GND_net), .I1(n14897[3]), .I2(n375_adj_4432), 
            .I3(n50949), .O(n14058[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_6 (.CI(n50949), .I0(n14897[3]), .I1(n375_adj_4432), 
            .CO(n50950));
    SB_LUT4 add_6103_5_lut (.I0(GND_net), .I1(n14897[2]), .I2(n302), .I3(n50948), 
            .O(n14058[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_13_i17_2_lut (.I0(n48[8]), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4632));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_18_i702_2_lut (.I0(\Ki[14] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4633));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i320_2_lut (.I0(\Ki[6] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4534));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Kp[14] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Kp[15] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_9_add_2_18 (.CI(n50355), .I0(setpoint[16]), .I1(n7), 
            .CO(n50356));
    SB_CARRY add_6103_5 (.CI(n50948), .I0(n14897[2]), .I1(n302), .CO(n50949));
    SB_LUT4 sub_9_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n50354), .O(n105[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6103_4_lut (.I0(GND_net), .I1(n14897[1]), .I2(n229), .I3(n50947), 
            .O(n14058[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i751_2_lut (.I0(\Ki[15] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4634));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i232_2_lut (.I0(\Kp[4] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4532));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_952 (.I0(n105[22]), .I1(n20122[1]), .I2(n4_adj_4635), 
            .I3(\Kp[3] ), .O(n20063[2]));   // verilog/motorControl.v(55[22:28])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'hc66c;
    SB_LUT4 mult_18_i369_2_lut (.I0(\Ki[7] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[13]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i416_2_lut (.I0(\Kp[8] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4529));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_9_add_2_17 (.CI(n50354), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n50355));
    SB_CARRY add_6103_4 (.CI(n50947), .I0(n14897[1]), .I1(n229), .CO(n50948));
    SB_LUT4 add_6103_3_lut (.I0(GND_net), .I1(n14897[0]), .I2(n156_adj_4431), 
            .I3(n50946), .O(n14058[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_3 (.CI(n50946), .I0(n14897[0]), .I1(n156_adj_4431), 
            .CO(n50947));
    SB_LUT4 sub_9_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n50353), .O(n105[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_16 (.CI(n50353), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n50354));
    SB_LUT4 mult_17_i465_2_lut (.I0(\Kp[9] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4528));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i4_3_lut (.I0(n48[3]), .I1(n49[3]), .I2(n182), .I3(GND_net), 
            .O(n208[3]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i4_3_lut (.I0(n208[3]), .I1(IntegralLimit[3]), .I2(n156), 
            .I3(GND_net), .O(n233[3]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i55_2_lut (.I0(\Ki[1] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4527));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i8_2_lut (.I0(\Ki[0] ), .I1(n233[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4526));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i418_2_lut (.I0(\Ki[8] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_9_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n50352), .O(n105[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n29696), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_CARRY add_6403_9 (.CI(n51907), .I0(n19547[6]), .I1(n624_c), .CO(n51908));
    SB_LUT4 add_6103_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n14058[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6103_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6103_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n50946));
    SB_LUT4 add_6433_10_lut (.I0(GND_net), .I1(n19823[7]), .I2(n700), 
            .I3(n50945), .O(n19665[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_15 (.CI(n50352), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n50353));
    SB_LUT4 add_6403_8_lut (.I0(GND_net), .I1(n19547[5]), .I2(n551_c), 
            .I3(n51906), .O(n19328[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6403_8 (.CI(n51906), .I0(n19547[5]), .I1(n551_c), .CO(n51907));
    SB_LUT4 add_6403_7_lut (.I0(GND_net), .I1(n19547[4]), .I2(n478_c), 
            .I3(n51905), .O(n19328[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6433_9_lut (.I0(GND_net), .I1(n19823[6]), .I2(n627), .I3(n50944), 
            .O(n19665[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6433_9 (.CI(n50944), .I0(n19823[6]), .I1(n627), .CO(n50945));
    SB_CARRY add_6403_7 (.CI(n51905), .I0(n19547[4]), .I1(n478_c), .CO(n51906));
    SB_LUT4 add_6403_6_lut (.I0(GND_net), .I1(n19547[3]), .I2(n405_c), 
            .I3(n51904), .O(n19328[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6403_6 (.CI(n51904), .I0(n19547[3]), .I1(n405_c), .CO(n51905));
    SB_LUT4 add_6403_5_lut (.I0(GND_net), .I1(n19547[2]), .I2(n332_c), 
            .I3(n51903), .O(n19328[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6403_5 (.CI(n51903), .I0(n19547[2]), .I1(n332_c), .CO(n51904));
    SB_LUT4 add_6403_4_lut (.I0(GND_net), .I1(n19547[1]), .I2(n259_c), 
            .I3(n51902), .O(n19328[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6433_8_lut (.I0(GND_net), .I1(n19823[5]), .I2(n554), .I3(n50943), 
            .O(n19665[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_9_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n50351), .O(n105[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_14 (.CI(n50351), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n50352));
    SB_CARRY add_6403_4 (.CI(n51902), .I0(n19547[1]), .I1(n259_c), .CO(n51903));
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n29668), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n29667), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n29665), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_LUT4 add_6403_3_lut (.I0(GND_net), .I1(n19547[0]), .I2(n186_c), 
            .I3(n51901), .O(n19328[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6403_3 (.CI(n51901), .I0(n19547[0]), .I1(n186_c), .CO(n51902));
    SB_LUT4 add_6403_2_lut (.I0(GND_net), .I1(n44), .I2(n113_c), .I3(GND_net), 
            .O(n19328[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6403_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n29663), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_CARRY add_6403_2 (.CI(GND_net), .I0(n44), .I1(n113_c), .CO(n51901));
    SB_LUT4 add_6199_19_lut (.I0(GND_net), .I1(n16697[16]), .I2(GND_net), 
            .I3(n51900), .O(n16053[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6199_18_lut (.I0(GND_net), .I1(n16697[15]), .I2(GND_net), 
            .I3(n51899), .O(n16053[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_18 (.CI(n51899), .I0(n16697[15]), .I1(GND_net), 
            .CO(n51900));
    SB_LUT4 add_6199_17_lut (.I0(GND_net), .I1(n16697[14]), .I2(GND_net), 
            .I3(n51898), .O(n16053[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n29662), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n29661), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n29660), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_CARRY add_6199_17 (.CI(n51898), .I0(n16697[14]), .I1(GND_net), 
            .CO(n51899));
    SB_CARRY add_6433_8 (.CI(n50943), .I0(n19823[5]), .I1(n554), .CO(n50944));
    SB_LUT4 add_6433_7_lut (.I0(GND_net), .I1(n19823[4]), .I2(n481_adj_4637), 
            .I3(n50942), .O(n19665[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6433_7 (.CI(n50942), .I0(n19823[4]), .I1(n481_adj_4637), 
            .CO(n50943));
    SB_LUT4 add_6433_6_lut (.I0(GND_net), .I1(n19823[3]), .I2(n408), .I3(n50941), 
            .O(n19665[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6199_16_lut (.I0(GND_net), .I1(n16697[13]), .I2(n1111), 
            .I3(n51897), .O(n16053[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_16 (.CI(n51897), .I0(n16697[13]), .I1(n1111), .CO(n51898));
    SB_CARRY add_6433_6 (.CI(n50941), .I0(n19823[3]), .I1(n408), .CO(n50942));
    SB_LUT4 sub_9_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n50350), .O(n105[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_24_i45_2_lut (.I0(PWMLimit[22]), .I1(n353[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4638));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6433_5_lut (.I0(GND_net), .I1(n19823[2]), .I2(n335), .I3(n50940), 
            .O(n19665[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6433_5 (.CI(n50940), .I0(n19823[2]), .I1(n335), .CO(n50941));
    SB_CARRY sub_9_add_2_13 (.CI(n50350), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n50351));
    SB_LUT4 sub_9_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n50349), .O(n105[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_24_i25_2_lut (.I0(PWMLimit[12]), .I1(n353[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4639));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_24_i31_2_lut (.I0(PWMLimit[15]), .I1(n353[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4640));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_24_i27_2_lut (.I0(PWMLimit[13]), .I1(n353[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4641));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_24_i29_2_lut (.I0(PWMLimit[14]), .I1(n353[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4642));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_24_i19_2_lut (.I0(PWMLimit[9]), .I1(n353[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4643));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_24_i21_2_lut (.I0(PWMLimit[10]), .I1(n353[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4644));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i21_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n29632), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_LUT4 add_6199_15_lut (.I0(GND_net), .I1(n16697[12]), .I2(n1038), 
            .I3(n51896), .O(n16053[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_15 (.CI(n51896), .I0(n16697[12]), .I1(n1038), .CO(n51897));
    SB_LUT4 add_6199_14_lut (.I0(GND_net), .I1(n16697[11]), .I2(n965), 
            .I3(n51895), .O(n16053[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_12 (.CI(n50349), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n50350));
    SB_LUT4 LessThan_24_i23_2_lut (.I0(PWMLimit[11]), .I1(n353[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4645));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_9_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n50348), .O(n105[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_24_i15_2_lut (.I0(PWMLimit[7]), .I1(n353[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4646));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_24_i17_2_lut (.I0(PWMLimit[8]), .I1(n353[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4647));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6433_4_lut (.I0(GND_net), .I1(n19823[1]), .I2(n262), .I3(n50939), 
            .O(n19665[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6433_4 (.CI(n50939), .I0(n19823[1]), .I1(n262), .CO(n50940));
    SB_LUT4 add_6334_14_lut (.I0(GND_net), .I1(n18754[11]), .I2(n980), 
            .I3(n50700), .O(n18391[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6334_13_lut (.I0(GND_net), .I1(n18754[10]), .I2(n907), 
            .I3(n50699), .O(n18391[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_14 (.CI(n51895), .I0(n16697[11]), .I1(n965), .CO(n51896));
    SB_CARRY add_6334_13 (.CI(n50699), .I0(n18754[10]), .I1(n907), .CO(n50700));
    SB_LUT4 add_6433_3_lut (.I0(GND_net), .I1(n19823[0]), .I2(n189_adj_4648), 
            .I3(n50938), .O(n19665[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_11 (.CI(n50348), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n50349));
    SB_LUT4 sub_9_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(n10), 
            .I3(n50347), .O(n105[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_10 (.CI(n50347), .I0(setpoint[8]), .I1(n10), 
            .CO(n50348));
    SB_LUT4 LessThan_24_i7_2_lut (.I0(PWMLimit[3]), .I1(n353[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4650));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6433_3 (.CI(n50938), .I0(n19823[0]), .I1(n189_adj_4648), 
            .CO(n50939));
    SB_LUT4 add_6433_2_lut (.I0(GND_net), .I1(n47_adj_4651), .I2(n116_adj_4652), 
            .I3(GND_net), .O(n19665[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6433_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6433_2 (.CI(GND_net), .I0(n47_adj_4651), .I1(n116_adj_4652), 
            .CO(n50938));
    SB_LUT4 add_6334_12_lut (.I0(GND_net), .I1(n18754[9]), .I2(n834_adj_4653), 
            .I3(n50698), .O(n18391[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_24_i9_2_lut (.I0(PWMLimit[4]), .I1(n353[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4654));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6334_12 (.CI(n50698), .I0(n18754[9]), .I1(n834_adj_4653), 
            .CO(n50699));
    SB_LUT4 add_6199_13_lut (.I0(GND_net), .I1(n16697[10]), .I2(n892), 
            .I3(n51894), .O(n16053[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6334_11_lut (.I0(GND_net), .I1(n18754[8]), .I2(n761_adj_4655), 
            .I3(n50697), .O(n18391[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6334_11 (.CI(n50697), .I0(n18754[8]), .I1(n761_adj_4655), 
            .CO(n50698));
    SB_LUT4 LessThan_24_i11_2_lut (.I0(PWMLimit[5]), .I1(n353[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4656));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6199_13 (.CI(n51894), .I0(n16697[10]), .I1(n892), .CO(n51895));
    SB_LUT4 add_6199_12_lut (.I0(GND_net), .I1(n16697[9]), .I2(n819), 
            .I3(n51893), .O(n16053[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_12 (.CI(n51893), .I0(n16697[9]), .I1(n819), .CO(n51894));
    SB_LUT4 LessThan_24_i13_2_lut (.I0(PWMLimit[6]), .I1(n353[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4657));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6199_11_lut (.I0(GND_net), .I1(n16697[8]), .I2(n746), 
            .I3(n51892), .O(n16053[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_11 (.CI(n51892), .I0(n16697[8]), .I1(n746), .CO(n51893));
    SB_LUT4 add_6199_10_lut (.I0(GND_net), .I1(n16697[7]), .I2(n673), 
            .I3(n51891), .O(n16053[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_10 (.CI(n51891), .I0(n16697[7]), .I1(n673), .CO(n51892));
    SB_LUT4 add_6199_9_lut (.I0(GND_net), .I1(n16697[6]), .I2(n600), .I3(n51890), 
            .O(n16053[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_2_lut (.I0(PWMLimit[2]), .I1(n353[2]), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_4658));
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51551_4_lut (.I0(n11_adj_4656), .I1(n9_adj_4654), .I2(n7_adj_4650), 
            .I3(n5_adj_4658), .O(n67277));
    defparam i51551_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51547_4_lut (.I0(n17_adj_4647), .I1(n15_adj_4646), .I2(n13_adj_4657), 
            .I3(n67277), .O(n67273));
    defparam i51547_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6199_9 (.CI(n51890), .I0(n16697[6]), .I1(n600), .CO(n51891));
    SB_LUT4 i53047_4_lut (.I0(n23_adj_4645), .I1(n21_adj_4644), .I2(n19_adj_4643), 
            .I3(n67273), .O(n68773));
    defparam i53047_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_24_i4_4_lut (.I0(PWMLimit[0]), .I1(n353[1]), .I2(PWMLimit[1]), 
            .I3(n353[0]), .O(n4_adj_4659));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52909_3_lut (.I0(n4_adj_4659), .I1(n353[13]), .I2(n27_adj_4641), 
            .I3(GND_net), .O(n68635));   // verilog/motorControl.v(57[18:33])
    defparam i52909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52910_3_lut (.I0(n68635), .I1(n353[14]), .I2(n29_adj_4642), 
            .I3(GND_net), .O(n68636));   // verilog/motorControl.v(57[18:33])
    defparam i52910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_24_i10_3_lut (.I0(n353[5]), .I1(n353[6]), .I2(n13_adj_4657), 
            .I3(GND_net), .O(n10_adj_4660));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52370_4_lut (.I0(n29_adj_4642), .I1(n27_adj_4641), .I2(n15_adj_4646), 
            .I3(n67275), .O(n68096));
    defparam i52370_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_24_i12_3_lut (.I0(n10_adj_4660), .I1(n353[7]), .I2(n15_adj_4646), 
            .I3(GND_net), .O(n12_adj_4661));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51897_3_lut (.I0(n68636), .I1(n353[15]), .I2(n31_adj_4640), 
            .I3(GND_net), .O(n67623));   // verilog/motorControl.v(57[18:33])
    defparam i51897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Kp[1] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4662));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Kp[0] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4663));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_9_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n50346), .O(n105[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_9 (.CI(n50346), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n50347));
    SB_LUT4 LessThan_24_i8_3_lut (.I0(n353[4]), .I1(n353[8]), .I2(n17_adj_4647), 
            .I3(GND_net), .O(n8_adj_4664));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6199_8_lut (.I0(GND_net), .I1(n16697[5]), .I2(n527), .I3(n51889), 
            .O(n16053[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_8 (.CI(n51889), .I0(n16697[5]), .I1(n527), .CO(n51890));
    SB_LUT4 LessThan_24_i6_3_lut (.I0(n353[2]), .I1(n353[3]), .I2(n7_adj_4650), 
            .I3(GND_net), .O(n6_adj_4665));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_24_i16_3_lut (.I0(n8_adj_4664), .I1(n353[9]), .I2(n19_adj_4643), 
            .I3(GND_net), .O(n16_adj_4666));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53312_4_lut (.I0(n16_adj_4666), .I1(n6_adj_4665), .I2(n19_adj_4643), 
            .I3(n67271), .O(n69038));   // verilog/motorControl.v(57[18:33])
    defparam i53312_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53313_3_lut (.I0(n69038), .I1(n353[10]), .I2(n21_adj_4644), 
            .I3(GND_net), .O(n69039));   // verilog/motorControl.v(57[18:33])
    defparam i53313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53200_3_lut (.I0(n69039), .I1(n353[11]), .I2(n23_adj_4645), 
            .I3(GND_net), .O(n68926));   // verilog/motorControl.v(57[18:33])
    defparam i53200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52372_4_lut (.I0(n29_adj_4642), .I1(n27_adj_4641), .I2(n25_adj_4639), 
            .I3(n68773), .O(n68098));
    defparam i52372_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52876_4_lut (.I0(n67623), .I1(n12_adj_4661), .I2(n31_adj_4640), 
            .I3(n68096), .O(n68602));   // verilog/motorControl.v(57[18:33])
    defparam i52876_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51895_3_lut (.I0(n68926), .I1(n353[12]), .I2(n25_adj_4639), 
            .I3(GND_net), .O(n67621));   // verilog/motorControl.v(57[18:33])
    defparam i51895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52878_4_lut (.I0(n67621), .I1(n68602), .I2(n31_adj_4640), 
            .I3(n68098), .O(n68604));   // verilog/motorControl.v(57[18:33])
    defparam i52878_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_24_i34_3_lut (.I0(n68604), .I1(n353[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n34));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6199_7_lut (.I0(GND_net), .I1(n16697[4]), .I2(n454_adj_4667), 
            .I3(n51888), .O(n16053[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_7 (.CI(n51888), .I0(n16697[4]), .I1(n454_adj_4667), 
            .CO(n51889));
    SB_LUT4 i22405_3_lut (.I0(n34), .I1(PWMLimit[17]), .I2(n353[17]), 
            .I3(GND_net), .O(n36));
    defparam i22405_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 add_6199_6_lut (.I0(GND_net), .I1(n16697[3]), .I2(n381_adj_4668), 
            .I3(n51887), .O(n16053[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_6 (.CI(n51887), .I0(n16697[3]), .I1(n381_adj_4668), 
            .CO(n51888));
    SB_LUT4 add_6199_5_lut (.I0(GND_net), .I1(n16697[2]), .I2(n308), .I3(n51886), 
            .O(n16053[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_5 (.CI(n51886), .I0(n16697[2]), .I1(n308), .CO(n51887));
    SB_LUT4 LessThan_24_i38_3_lut (.I0(n36), .I1(n353[18]), .I2(PWMLimit[18]), 
            .I3(GND_net), .O(n38_adj_4669));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6199_4_lut (.I0(GND_net), .I1(n16697[1]), .I2(n235_adj_4670), 
            .I3(n51885), .O(n16053[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_4 (.CI(n51885), .I0(n16697[1]), .I1(n235_adj_4670), 
            .CO(n51886));
    SB_LUT4 counter_1944_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n51645), .O(n52[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6334_10_lut (.I0(GND_net), .I1(n18754[7]), .I2(n688_adj_4672), 
            .I3(n50696), .O(n18391[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23382_3_lut (.I0(n38_adj_4669), .I1(PWMLimit[19]), .I2(n353[19]), 
            .I3(GND_net), .O(n40));
    defparam i23382_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 LessThan_24_i44_3_lut (.I0(n42), .I1(n353[22]), .I2(n45_adj_4638), 
            .I3(GND_net), .O(n44_adj_4673));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i44_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52879_4_lut (.I0(n44_adj_4673), .I1(n40), .I2(n45_adj_4638), 
            .I3(n67242), .O(n68605));   // verilog/motorControl.v(57[18:33])
    defparam i52879_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52880_3_lut (.I0(n68605), .I1(PWMLimit[23]), .I2(n353[23]), 
            .I3(GND_net), .O(n406));   // verilog/motorControl.v(57[18:33])
    defparam i52880_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(n353[20]), .I1(n433[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4674));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(n353[13]), .I1(n433[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4675));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i25_2_lut (.I0(n353[12]), .I1(n433[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4676));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(n353[11]), .I1(n433[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4677));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6199_3_lut (.I0(GND_net), .I1(n16697[0]), .I2(n162), .I3(n51884), 
            .O(n16053[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_3 (.CI(n51884), .I0(n16697[0]), .I1(n162), .CO(n51885));
    SB_CARRY add_6334_10 (.CI(n50696), .I0(n18754[7]), .I1(n688_adj_4672), 
            .CO(n50697));
    SB_LUT4 counter_1944_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n51644), .O(n52[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6199_2_lut (.I0(GND_net), .I1(n20_adj_4679), .I2(n89), 
            .I3(GND_net), .O(n16053[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6199_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6199_2 (.CI(GND_net), .I0(n20_adj_4679), .I1(n89), .CO(n51884));
    SB_LUT4 add_6334_9_lut (.I0(GND_net), .I1(n18754[6]), .I2(n615_adj_4680), 
            .I3(n50695), .O(n18391[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6334_9 (.CI(n50695), .I0(n18754[6]), .I1(n615_adj_4680), 
            .CO(n50696));
    SB_LUT4 LessThan_26_i21_2_lut (.I0(n353[10]), .I1(n433[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4681));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(n433[0]), .I1(n433[1]), .I2(n353[1]), 
            .I3(n353[0]), .O(n4_adj_4683));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(n353[7]), .I1(n433[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4684));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(n353[8]), .I1(n433[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4685));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(n353[9]), .I1(n433[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4686));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i9_2_lut (.I0(n353[4]), .I1(n433[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4687));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6233_18_lut (.I0(GND_net), .I1(n17271[15]), .I2(GND_net), 
            .I3(n51883), .O(n16697[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(n353[5]), .I1(n433[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4688));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(n353[6]), .I1(n433[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4689));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i7_2_lut (.I0(n353[3]), .I1(n433[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4690));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51510_4_lut (.I0(n13_adj_4689), .I1(n11_adj_4688), .I2(n9_adj_4687), 
            .I3(n7_adj_4690), .O(n67236));
    defparam i51510_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51505_4_lut (.I0(n19_adj_4686), .I1(n17_adj_4685), .I2(n15_adj_4684), 
            .I3(n67236), .O(n67231));
    defparam i51505_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n433[6]), .I1(n433[7]), .I2(n15_adj_4684), 
            .I3(GND_net), .O(n12_adj_4691));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27592_3_lut (.I0(n4_adj_4683), .I1(n353[2]), .I2(n433[2]), 
            .I3(GND_net), .O(n6_adj_4692));
    defparam i27592_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 LessThan_26_i14_3_lut (.I0(n12_adj_4691), .I1(n433[8]), .I2(n17_adj_4685), 
            .I3(GND_net), .O(n14_adj_4693));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i10_3_lut (.I0(n433[5]), .I1(n433[9]), .I2(n19_adj_4686), 
            .I3(GND_net), .O(n10_adj_4694));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i8_3_lut (.I0(n433[3]), .I1(n433[4]), .I2(n9_adj_4687), 
            .I3(GND_net), .O(n8_adj_4695));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i18_3_lut (.I0(n10_adj_4694), .I1(n433[10]), .I2(n21_adj_4681), 
            .I3(GND_net), .O(n18_adj_4696));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53314_4_lut (.I0(n18_adj_4696), .I1(n8_adj_4695), .I2(n21_adj_4681), 
            .I3(n67229), .O(n69040));   // verilog/motorControl.v(59[27:43])
    defparam i53314_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53315_3_lut (.I0(n69040), .I1(n433[11]), .I2(n23_adj_4677), 
            .I3(GND_net), .O(n69041));   // verilog/motorControl.v(59[27:43])
    defparam i53315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53198_3_lut (.I0(n69041), .I1(n433[12]), .I2(n25_adj_4676), 
            .I3(GND_net), .O(n68924));   // verilog/motorControl.v(59[27:43])
    defparam i53198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53043_4_lut (.I0(n25_adj_4676), .I1(n23_adj_4677), .I2(n21_adj_4681), 
            .I3(n67231), .O(n68769));
    defparam i53043_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53395_4_lut (.I0(n14_adj_4693), .I1(n6_adj_4692), .I2(n17_adj_4685), 
            .I3(n67234), .O(n69121));   // verilog/motorControl.v(59[27:43])
    defparam i53395_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51901_3_lut (.I0(n68924), .I1(n433[13]), .I2(n27_adj_4675), 
            .I3(GND_net), .O(n67627));   // verilog/motorControl.v(59[27:43])
    defparam i51901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53472_4_lut (.I0(n67627), .I1(n69121), .I2(n27_adj_4675), 
            .I3(n68769), .O(n69198));   // verilog/motorControl.v(59[27:43])
    defparam i53472_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53473_3_lut (.I0(n69198), .I1(n433[14]), .I2(n353[14]), .I3(GND_net), 
            .O(n69199));   // verilog/motorControl.v(59[27:43])
    defparam i53473_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29619), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_LUT4 add_6233_17_lut (.I0(GND_net), .I1(n17271[14]), .I2(GND_net), 
            .I3(n51882), .O(n16697[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53392_3_lut (.I0(n69199), .I1(n433[15]), .I2(n353[15]), .I3(GND_net), 
            .O(n69118));   // verilog/motorControl.v(59[27:43])
    defparam i53392_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6233_17 (.CI(n51882), .I0(n17271[14]), .I1(GND_net), 
            .CO(n51883));
    SB_LUT4 i53367_3_lut (.I0(n69118), .I1(n433[16]), .I2(n353[16]), .I3(GND_net), 
            .O(n34_adj_4697));   // verilog/motorControl.v(59[27:43])
    defparam i53367_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i22409_3_lut (.I0(n34_adj_4697), .I1(n353[17]), .I2(n433[17]), 
            .I3(GND_net), .O(n36_adj_4698));
    defparam i22409_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 LessThan_26_i40_3_lut (.I0(n38_adj_4699), .I1(n433[20]), .I2(n41_adj_4674), 
            .I3(GND_net), .O(n40_adj_4700));   // verilog/motorControl.v(59[27:43])
    defparam LessThan_26_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53316_4_lut (.I0(n40_adj_4700), .I1(n36_adj_4698), .I2(n41_adj_4674), 
            .I3(n67216), .O(n69042));   // verilog/motorControl.v(59[27:43])
    defparam i53316_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53317_3_lut (.I0(n69042), .I1(n433[21]), .I2(n353[21]), .I3(GND_net), 
            .O(n69043));   // verilog/motorControl.v(59[27:43])
    defparam i53317_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53194_3_lut (.I0(n69043), .I1(n433[22]), .I2(n353[22]), .I3(GND_net), 
            .O(n68920));   // verilog/motorControl.v(59[27:43])
    defparam i53194_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51905_3_lut (.I0(n68920), .I1(n353[23]), .I2(n433[23]), .I3(GND_net), 
            .O(n432));   // verilog/motorControl.v(59[27:43])
    defparam i51905_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut (.I0(control_update), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n27916));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY counter_1944_add_4_32 (.CI(n51644), .I0(GND_net), .I1(counter[30]), 
            .CO(n51645));
    SB_LUT4 mux_28_i1_3_lut (.I0(n353[0]), .I1(n433[0]), .I2(n432), .I3(GND_net), 
            .O(n458[0]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_28_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_29_i1_3_lut (.I0(n458[0]), .I1(PWMLimit[0]), .I2(n406), 
            .I3(GND_net), .O(n483[0]));   // verilog/motorControl.v(59[24] 61[18])
    defparam mux_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_4_lut (.I0(setpoint[0]), .I1(n483[0]), .I2(n15), 
            .I3(n405), .O(duty_23__N_3602[0]));   // verilog/motorControl.v(45[18] 66[12])
    defparam duty_23__I_0_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_953 (.I0(counter[2]), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4701));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12_adj_4702));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6233_16_lut (.I0(GND_net), .I1(n17271[13]), .I2(n1114), 
            .I3(n51881), .O(n16697[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4909_4_lut (.I0(counter[5]), .I1(counter[7]), .I2(n12_adj_4702), 
            .I3(n8_adj_4701), .O(n16_adj_4703));
    defparam i4909_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_4704));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut (.I0(counter[23]), .I1(counter[25]), .I2(counter[26]), 
            .I3(counter[15]), .O(n61067));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(counter[22]), .I1(n61067), .I2(counter[17]), 
            .I3(GND_net), .O(n8_adj_4705));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_954 (.I0(counter[12]), .I1(n10_adj_4704), .I2(n16_adj_4703), 
            .I3(counter[8]), .O(n60808));
    defparam i5_4_lut_adj_954.LUT_INIT = 16'h8880;
    SB_LUT4 i1_4_lut_adj_955 (.I0(counter[21]), .I1(n60808), .I2(n8_adj_4705), 
            .I3(counter[18]), .O(n10_adj_4706));
    defparam i1_4_lut_adj_955.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_956 (.I0(counter[16]), .I1(counter[19]), .I2(counter[28]), 
            .I3(counter[27]), .O(n12_adj_4707));
    defparam i3_4_lut_adj_956.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(counter[20]), .I1(counter[14]), .I2(counter[30]), 
            .I3(n10_adj_4706), .O(n16_adj_4708));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(counter[24]), .I1(counter[29]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4709));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28476_4_lut (.I0(n11_adj_4709), .I1(counter[31]), .I2(n16_adj_4708), 
            .I3(n12_adj_4707), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:41])
    defparam i28476_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Kp[5] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6334_8_lut (.I0(GND_net), .I1(n18754[5]), .I2(n542_adj_4710), 
            .I3(n50694), .O(n18391[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i396_2_lut (.I0(\Ki[8] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i396_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6334_8 (.CI(n50694), .I0(n18754[5]), .I1(n542_adj_4710), 
            .CO(n50695));
    SB_LUT4 sub_9_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n50345), .O(n105[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6334_7_lut (.I0(GND_net), .I1(n18754[4]), .I2(n469_adj_4711), 
            .I3(n50693), .O(n18391[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6334_7 (.CI(n50693), .I0(n18754[4]), .I1(n469_adj_4711), 
            .CO(n50694));
    SB_CARRY add_6233_16 (.CI(n51881), .I0(n17271[13]), .I1(n1114), .CO(n51882));
    SB_LUT4 add_6334_6_lut (.I0(GND_net), .I1(n18754[3]), .I2(n396_adj_4712), 
            .I3(n50692), .O(n18391[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6233_15_lut (.I0(GND_net), .I1(n17271[12]), .I2(n1041), 
            .I3(n51880), .O(n16697[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n51643), .O(n52[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1944__i0 (.Q(counter[0]), .C(clk16MHz), .D(n52[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_CARRY add_6233_15 (.CI(n51880), .I0(n17271[12]), .I1(n1041), .CO(n51881));
    SB_CARRY counter_1944_add_4_31 (.CI(n51643), .I0(GND_net), .I1(counter[29]), 
            .CO(n51644));
    SB_LUT4 counter_1944_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n51642), .O(n52[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6233_14_lut (.I0(GND_net), .I1(n17271[11]), .I2(n968), 
            .I3(n51879), .O(n16697[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_30 (.CI(n51642), .I0(GND_net), .I1(counter[28]), 
            .CO(n51643));
    SB_CARRY add_6233_14 (.CI(n51879), .I0(n17271[11]), .I1(n968), .CO(n51880));
    SB_LUT4 counter_1944_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n51641), .O(n52[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6233_13_lut (.I0(GND_net), .I1(n17271[10]), .I2(n895), 
            .I3(n51878), .O(n16697[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_13 (.CI(n51878), .I0(n17271[10]), .I1(n895), .CO(n51879));
    SB_CARRY counter_1944_add_4_29 (.CI(n51641), .I0(GND_net), .I1(counter[27]), 
            .CO(n51642));
    SB_LUT4 add_6233_12_lut (.I0(GND_net), .I1(n17271[9]), .I2(n822), 
            .I3(n51877), .O(n16697[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_12 (.CI(n51877), .I0(n17271[9]), .I1(n822), .CO(n51878));
    SB_LUT4 counter_1944_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n51640), .O(n52[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_28 (.CI(n51640), .I0(GND_net), .I1(counter[26]), 
            .CO(n51641));
    SB_LUT4 add_6233_11_lut (.I0(GND_net), .I1(n17271[8]), .I2(n749), 
            .I3(n51876), .O(n16697[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_11 (.CI(n51876), .I0(n17271[8]), .I1(n749), .CO(n51877));
    SB_LUT4 add_6233_10_lut (.I0(GND_net), .I1(n17271[7]), .I2(n676), 
            .I3(n51875), .O(n16697[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_10 (.CI(n51875), .I0(n17271[7]), .I1(n676), .CO(n51876));
    SB_LUT4 add_6233_9_lut (.I0(GND_net), .I1(n17271[6]), .I2(n603_adj_4718), 
            .I3(n51874), .O(n16697[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1944__i31 (.Q(counter[31]), .C(clk16MHz), .D(n52[31]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i30 (.Q(counter[30]), .C(clk16MHz), .D(n52[30]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i29 (.Q(counter[29]), .C(clk16MHz), .D(n52[29]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i28 (.Q(counter[28]), .C(clk16MHz), .D(n52[28]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i27 (.Q(counter[27]), .C(clk16MHz), .D(n52[27]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i26 (.Q(counter[26]), .C(clk16MHz), .D(n52[26]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i25 (.Q(counter[25]), .C(clk16MHz), .D(n52[25]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i24 (.Q(counter[24]), .C(clk16MHz), .D(n52[24]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i23 (.Q(counter[23]), .C(clk16MHz), .D(n52[23]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i22 (.Q(counter[22]), .C(clk16MHz), .D(n52[22]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i21 (.Q(counter[21]), .C(clk16MHz), .D(n52[21]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i20 (.Q(counter[20]), .C(clk16MHz), .D(n52[20]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i19 (.Q(counter[19]), .C(clk16MHz), .D(n52[19]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i18 (.Q(counter[18]), .C(clk16MHz), .D(n52[18]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i17 (.Q(counter[17]), .C(clk16MHz), .D(n52[17]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i16 (.Q(counter[16]), .C(clk16MHz), .D(n52[16]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i15 (.Q(counter[15]), .C(clk16MHz), .D(n52[15]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i14 (.Q(counter[14]), .C(clk16MHz), .D(n52[14]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i13 (.Q(counter[13]), .C(clk16MHz), .D(n52[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i12 (.Q(counter[12]), .C(clk16MHz), .D(n52[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i11 (.Q(counter[11]), .C(clk16MHz), .D(n52[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i10 (.Q(counter[10]), .C(clk16MHz), .D(n52[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i9 (.Q(counter[9]), .C(clk16MHz), .D(n52[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i8 (.Q(counter[8]), .C(clk16MHz), .D(n52[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i7 (.Q(counter[7]), .C(clk16MHz), .D(n52[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i6 (.Q(counter[6]), .C(clk16MHz), .D(n52[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i5 (.Q(counter[5]), .C(clk16MHz), .D(n52[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i4 (.Q(counter[4]), .C(clk16MHz), .D(n52[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i3 (.Q(counter[3]), .C(clk16MHz), .D(n52[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i2 (.Q(counter[2]), .C(clk16MHz), .D(n52[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_1944__i1 (.Q(counter[1]), .C(clk16MHz), .D(n52[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_CARRY add_6334_6 (.CI(n50692), .I0(n18754[3]), .I1(n396_adj_4712), 
            .CO(n50693));
    SB_LUT4 mult_18_i445_2_lut (.I0(\Ki[9] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i445_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6233_9 (.CI(n51874), .I0(n17271[6]), .I1(n603_adj_4718), 
            .CO(n51875));
    SB_LUT4 counter_1944_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n51639), .O(n52[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i267_2_lut (.I0(\Ki[5] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i494_2_lut (.I0(\Ki[10] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6334_5_lut (.I0(GND_net), .I1(n18754[2]), .I2(n323_adj_4738), 
            .I3(n50691), .O(n18391[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_8 (.CI(n50345), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n50346));
    SB_CARRY add_6334_5 (.CI(n50691), .I0(n18754[2]), .I1(n323_adj_4738), 
            .CO(n50692));
    SB_LUT4 add_6334_4_lut (.I0(GND_net), .I1(n18754[1]), .I2(n250_adj_4739), 
            .I3(n50690), .O(n18391[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i543_2_lut (.I0(\Ki[11] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i592_2_lut (.I0(\Ki[12] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i316_2_lut (.I0(\Ki[6] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_9_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n50344), .O(n105[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6233_8_lut (.I0(GND_net), .I1(n17271[5]), .I2(n530_adj_4740), 
            .I3(n51873), .O(n16697[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_7 (.CI(n50344), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n50345));
    SB_LUT4 sub_9_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n50343), .O(n105[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_9_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6334_4 (.CI(n50690), .I0(n18754[1]), .I1(n250_adj_4739), 
            .CO(n50691));
    SB_LUT4 mult_17_i308_2_lut (.I0(\Kp[6] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6233_8 (.CI(n51873), .I0(n17271[5]), .I1(n530_adj_4740), 
            .CO(n51874));
    SB_LUT4 mult_18_i641_2_lut (.I0(\Ki[13] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i690_2_lut (.I0(\Ki[14] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6233_7_lut (.I0(GND_net), .I1(n17271[4]), .I2(n457_adj_4741), 
            .I3(n51872), .O(n16697[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i365_2_lut (.I0(\Ki[7] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i414_2_lut (.I0(\Ki[8] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i2_3_lut (.I0(n48[1]), .I1(n49[1]), .I2(n182), .I3(GND_net), 
            .O(n208[1]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6334_3_lut (.I0(GND_net), .I1(n18754[0]), .I2(n177_adj_4742), 
            .I3(n50689), .O(n18391[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6334_3 (.CI(n50689), .I0(n18754[0]), .I1(n177_adj_4742), 
            .CO(n50690));
    SB_LUT4 mux_16_i2_3_lut (.I0(n208[1]), .I1(IntegralLimit[1]), .I2(n156), 
            .I3(GND_net), .O(n233[1]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i739_2_lut (.I0(\Ki[15] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i739_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6233_7 (.CI(n51872), .I0(n17271[4]), .I1(n457_adj_4741), 
            .CO(n51873));
    SB_LUT4 mult_18_i463_2_lut (.I0(\Ki[9] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i512_2_lut (.I0(\Ki[10] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6334_2_lut (.I0(GND_net), .I1(n35_adj_4743), .I2(n104_adj_4744), 
            .I3(GND_net), .O(n18391[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6334_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6334_2 (.CI(GND_net), .I0(n35_adj_4743), .I1(n104_adj_4744), 
            .CO(n50689));
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30459), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_CARRY sub_9_add_2_6 (.CI(n50343), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n50344));
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30458), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30457), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30456), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30450), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30449), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30447), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30446), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30444), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_CARRY counter_1944_add_4_27 (.CI(n51639), .I0(GND_net), .I1(counter[25]), 
            .CO(n51640));
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30411), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30410), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30407), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30406), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_LUT4 counter_1944_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n51638), .O(n52[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_26 (.CI(n51638), .I0(GND_net), .I1(counter[24]), 
            .CO(n51639));
    SB_CARRY sub_9_add_2_5 (.CI(n50342), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n50343));
    SB_LUT4 add_6233_6_lut (.I0(GND_net), .I1(n17271[3]), .I2(n384_adj_4745), 
            .I3(n51871), .O(n16697[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_6 (.CI(n51871), .I0(n17271[3]), .I1(n384_adj_4745), 
            .CO(n51872));
    SB_LUT4 add_6233_5_lut (.I0(GND_net), .I1(n17271[2]), .I2(n311_adj_4746), 
            .I3(n51870), .O(n16697[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n51637), .O(n52[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_5 (.CI(n51870), .I0(n17271[2]), .I1(n311_adj_4746), 
            .CO(n51871));
    SB_LUT4 add_6233_4_lut (.I0(GND_net), .I1(n17271[1]), .I2(n238_adj_4747), 
            .I3(n51869), .O(n16697[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_4 (.CI(n51869), .I0(n17271[1]), .I1(n238_adj_4747), 
            .CO(n51870));
    SB_CARRY sub_9_add_2_4 (.CI(n50341), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n50342));
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30227), .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_LUT4 add_6233_3_lut (.I0(GND_net), .I1(n17271[0]), .I2(n165_adj_4748), 
            .I3(n51868), .O(n16697[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6233_3 (.CI(n51868), .I0(n17271[0]), .I1(n165_adj_4748), 
            .CO(n51869));
    SB_LUT4 add_6233_2_lut (.I0(GND_net), .I1(n23_adj_4749), .I2(n92_adj_4750), 
            .I3(GND_net), .O(n16697[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6233_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_25 (.CI(n51637), .I0(GND_net), .I1(counter[23]), 
            .CO(n51638));
    SB_CARRY add_6233_2 (.CI(GND_net), .I0(n23_adj_4749), .I1(n92_adj_4750), 
            .CO(n51868));
    SB_LUT4 mult_18_i104_2_lut (.I0(\Ki[2] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4525));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6422_10_lut (.I0(GND_net), .I1(n19726[7]), .I2(n700_adj_4751), 
            .I3(n51867), .O(n19547[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i281_2_lut (.I0(\Kp[5] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4524));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i234_2_lut (.I0(\Kp[4] ), .I1(n105[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_957 (.I0(n20122[1]), .I1(n6_adj_4752), .I2(n347), 
            .I3(n58043), .O(n20063[3]));   // verilog/motorControl.v(55[22:28])
    defparam i1_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 mult_18_i153_2_lut (.I0(\Ki[3] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4523));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6422_9_lut (.I0(GND_net), .I1(n19726[6]), .I2(n627_adj_4753), 
            .I3(n51866), .O(n19547[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Kp[1] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Kp[0] ), .I1(n105[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4522));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_958 (.I0(n62906), .I1(n105[23]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4635));   // verilog/motorControl.v(55[22:28])
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h8888;
    SB_LUT4 i36212_4_lut (.I0(n20122[1]), .I1(\Kp[3] ), .I2(n4_adj_4635), 
            .I3(n105[22]), .O(n6_adj_4752));   // verilog/motorControl.v(55[22:28])
    defparam i36212_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 mult_17_i40_2_lut (.I0(\Kp[0] ), .I1(n105[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62_c));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i40_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6422_9 (.CI(n51866), .I0(n19726[6]), .I1(n627_adj_4753), 
            .CO(n51867));
    SB_LUT4 counter_1944_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n51636), .O(n52[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_24 (.CI(n51636), .I0(GND_net), .I1(counter[22]), 
            .CO(n51637));
    SB_LUT4 counter_1944_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n51635), .O(n52[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6422_8_lut (.I0(GND_net), .I1(n19726[5]), .I2(n554_adj_4754), 
            .I3(n51865), .O(n19547[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6422_8 (.CI(n51865), .I0(n19726[5]), .I1(n554_adj_4754), 
            .CO(n51866));
    SB_CARRY counter_1944_add_4_23 (.CI(n51635), .I0(GND_net), .I1(counter[21]), 
            .CO(n51636));
    SB_LUT4 i36151_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n50049));   // verilog/motorControl.v(55[22:28])
    defparam i36151_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(\Kp[1] ), .I1(\Kp[2] ), .I2(\Kp[0] ), .I3(GND_net), 
            .O(n62906));   // verilog/motorControl.v(55[22:28])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i47763_3_lut (.I0(n105[23]), .I1(n62906), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n58043));   // verilog/motorControl.v(55[22:28])
    defparam i47763_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 add_6422_7_lut (.I0(GND_net), .I1(n19726[4]), .I2(n481_adj_4755), 
            .I3(n51864), .O(n19547[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6422_7 (.CI(n51864), .I0(n19726[4]), .I1(n481_adj_4755), 
            .CO(n51865));
    SB_LUT4 add_6422_6_lut (.I0(GND_net), .I1(n19726[3]), .I2(n408_adj_4756), 
            .I3(n51863), .O(n19547[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6422_6 (.CI(n51863), .I0(n19726[3]), .I1(n408_adj_4756), 
            .CO(n51864));
    SB_LUT4 counter_1944_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n51634), .O(n52[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6422_5_lut (.I0(GND_net), .I1(n19726[2]), .I2(n335_adj_4757), 
            .I3(n51862), .O(n19547[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Kp[2] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4758));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6422_5 (.CI(n51862), .I0(n19726[2]), .I1(n335_adj_4757), 
            .CO(n51863));
    SB_LUT4 add_6422_4_lut (.I0(GND_net), .I1(n19726[1]), .I2(n262_adj_4759), 
            .I3(n51861), .O(n19547[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36160_3_lut (.I0(n105[23]), .I1(n50063), .I2(n50278), .I3(GND_net), 
            .O(n20122[1]));   // verilog/motorControl.v(55[22:28])
    defparam i36160_3_lut.LUT_INIT = 16'h6c6c;
    SB_CARRY add_6422_4 (.CI(n51861), .I0(n19726[1]), .I1(n262_adj_4759), 
            .CO(n51862));
    SB_LUT4 add_6422_3_lut (.I0(GND_net), .I1(n19726[0]), .I2(n189_adj_4758), 
            .I3(n51860), .O(n19547[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i330_2_lut (.I0(\Kp[6] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4521));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_22 (.CI(n51634), .I0(GND_net), .I1(counter[20]), 
            .CO(n51635));
    SB_LUT4 i1_4_lut_adj_959 (.I0(n105[23]), .I1(\Kp[5] ), .I2(n50278), 
            .I3(n105[22]), .O(n62896));   // verilog/motorControl.v(55[22:28])
    defparam i1_4_lut_adj_959.LUT_INIT = 16'hc60a;
    SB_CARRY add_6422_3 (.CI(n51860), .I0(n19726[0]), .I1(n189_adj_4758), 
            .CO(n51861));
    SB_LUT4 i1_rep_256_2_lut (.I0(n20122[1]), .I1(n58043), .I2(GND_net), 
            .I3(GND_net), .O(n70741));   // verilog/motorControl.v(55[22:28])
    defparam i1_rep_256_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_960 (.I0(n50063), .I1(n62896), .I2(\Kp[4] ), 
            .I3(n105[23]), .O(n62900));   // verilog/motorControl.v(55[22:28])
    defparam i1_4_lut_adj_960.LUT_INIT = 16'h9666;
    SB_LUT4 i36220_4_lut (.I0(n70741), .I1(\Kp[4] ), .I2(n6_adj_4752), 
            .I3(n105[22]), .O(n8_adj_4760));   // verilog/motorControl.v(55[22:28])
    defparam i36220_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_17_add_1221_24_lut (.I0(n105[23]), .I1(n12072[21]), .I2(GND_net), 
            .I3(n51105), .O(n11613[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6422_2_lut (.I0(GND_net), .I1(n47_adj_4663), .I2(n116_adj_4662), 
            .I3(GND_net), .O(n19547[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6422_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_9_add_2_3 (.CI(n50340), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n50341));
    SB_LUT4 mult_17_i177_2_lut (.I0(\Kp[3] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4759));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6422_2 (.CI(GND_net), .I0(n47_adj_4663), .I1(n116_adj_4662), 
            .CO(n51860));
    SB_LUT4 add_6265_17_lut (.I0(GND_net), .I1(n17779[14]), .I2(GND_net), 
            .I3(n51859), .O(n17271[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n51633), .O(n52[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Kp[4] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4757));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36173_4_lut (.I0(n20122[1]), .I1(\Kp[3] ), .I2(n62906), .I3(n105[23]), 
            .O(n6_adj_4761));   // verilog/motorControl.v(55[22:28])
    defparam i36173_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_961 (.I0(n6_adj_4761), .I1(n8_adj_4760), .I2(n62900), 
            .I3(n58043), .O(n60191));   // verilog/motorControl.v(55[22:28])
    defparam i1_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Kp[5] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4756));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_23_lut (.I0(GND_net), .I1(n12072[20]), .I2(GND_net), 
            .I3(n51104), .O(n258[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_23 (.CI(n51104), .I0(n12072[20]), .I1(GND_net), 
            .CO(n51105));
    SB_LUT4 mult_18_i467_2_lut (.I0(\Ki[9] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_21 (.CI(n51633), .I0(GND_net), .I1(counter[19]), 
            .CO(n51634));
    SB_LUT4 counter_1944_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n51632), .O(n52[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_20 (.CI(n51632), .I0(GND_net), .I1(counter[18]), 
            .CO(n51633));
    SB_LUT4 counter_1944_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n51631), .O(n52[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Kp[10] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4519));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i563_2_lut (.I0(\Kp[11] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4518));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_9_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(n18), 
            .CO(n50340));
    SB_LUT4 mult_17_add_1221_22_lut (.I0(GND_net), .I1(n12072[19]), .I2(GND_net), 
            .I3(n51103), .O(n258[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_22 (.CI(n51103), .I0(n12072[19]), .I1(GND_net), 
            .CO(n51104));
    SB_LUT4 mult_17_add_1221_21_lut (.I0(GND_net), .I1(n12072[18]), .I2(GND_net), 
            .I3(n51102), .O(n258[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_19 (.CI(n51631), .I0(GND_net), .I1(counter[17]), 
            .CO(n51632));
    SB_LUT4 mult_17_i324_2_lut (.I0(\Kp[6] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4755));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1221_21 (.CI(n51102), .I0(n12072[18]), .I1(GND_net), 
            .CO(n51103));
    SB_LUT4 mult_17_i373_2_lut (.I0(\Kp[7] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4754));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Kp[12] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4517));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[14]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Kp[2] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[15]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_14_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[16]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Kp[3] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4511));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Kp[4] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4510));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Kp[5] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4508));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i202_2_lut (.I0(\Ki[4] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4507));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_20_lut (.I0(GND_net), .I1(n12072[17]), .I2(GND_net), 
            .I3(n51101), .O(n258[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Kp[6] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4506));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i251_2_lut (.I0(\Ki[5] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4505));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Kp[7] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4504));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[17]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Kp[8] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4753));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Kp[8] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4501));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i516_2_lut (.I0(\Ki[10] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i300_2_lut (.I0(\Ki[6] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4500));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1944_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n51630), .O(n52[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_18 (.CI(n51630), .I0(GND_net), .I1(counter[16]), 
            .CO(n51631));
    SB_LUT4 counter_1944_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n51629), .O(n52[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_17 (.CI(n51629), .I0(GND_net), .I1(counter[15]), 
            .CO(n51630));
    SB_LUT4 counter_1944_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n51628), .O(n52[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i565_2_lut (.I0(\Ki[11] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_16 (.CI(n51628), .I0(GND_net), .I1(counter[14]), 
            .CO(n51629));
    SB_LUT4 counter_1944_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n51627), .O(n52[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6265_16_lut (.I0(GND_net), .I1(n17779[13]), .I2(n1117_adj_4634), 
            .I3(n51858), .O(n17271[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_16 (.CI(n51858), .I0(n17779[13]), .I1(n1117_adj_4634), 
            .CO(n51859));
    SB_LUT4 unary_minus_14_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[18]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Kp[9] ), .I1(n105[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4751));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Kp[9] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4498));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_15 (.CI(n51627), .I0(GND_net), .I1(counter[13]), 
            .CO(n51628));
    SB_LUT4 add_6265_15_lut (.I0(GND_net), .I1(n17779[12]), .I2(n1044_adj_4633), 
            .I3(n51857), .O(n17271[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6142_20_lut (.I0(GND_net), .I1(n15656[17]), .I2(GND_net), 
            .I3(n50916), .O(n14897[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i13_3_lut (.I0(n48[12]), .I1(n49[12]), .I2(n182), .I3(GND_net), 
            .O(n208[12]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i13_3_lut (.I0(n208[12]), .I1(IntegralLimit[12]), .I2(n156), 
            .I3(GND_net), .O(n233[12]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i73_2_lut (.I0(\Ki[1] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4497));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i26_2_lut (.I0(\Ki[0] ), .I1(n233[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i63_2_lut (.I0(\Ki[1] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4750));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i16_2_lut (.I0(\Ki[0] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4749));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[19]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i349_2_lut (.I0(\Ki[7] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[20]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_15_i18_3_lut (.I0(n48[17]), .I1(n49[17]), .I2(n182), .I3(GND_net), 
            .O(n208[17]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i18_3_lut (.I0(n208[17]), .I1(IntegralLimit[17]), .I2(n156), 
            .I3(GND_net), .O(n233[17]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6265_15 (.CI(n51857), .I0(n17779[12]), .I1(n1044_adj_4633), 
            .CO(n51858));
    SB_LUT4 add_6265_14_lut (.I0(GND_net), .I1(n17779[11]), .I2(n971_adj_4601), 
            .I3(n51856), .O(n17271[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i83_2_lut (.I0(\Ki[1] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4494));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i36_2_lut (.I0(\Ki[0] ), .I1(n233[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4493));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Kp[10] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4492));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i398_2_lut (.I0(\Ki[8] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i132_2_lut (.I0(\Ki[2] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4491));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Kp[11] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4490));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1221_20 (.CI(n51101), .I0(n12072[17]), .I1(GND_net), 
            .CO(n51102));
    SB_CARRY add_6265_14 (.CI(n51856), .I0(n17779[11]), .I1(n971_adj_4601), 
            .CO(n51857));
    SB_LUT4 add_6142_19_lut (.I0(GND_net), .I1(n15656[16]), .I2(GND_net), 
            .I3(n50915), .O(n14897[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n51626), .O(n52[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_19 (.CI(n50915), .I0(n15656[16]), .I1(GND_net), 
            .CO(n50916));
    SB_LUT4 add_6265_13_lut (.I0(GND_net), .I1(n17779[10]), .I2(n898_adj_4590), 
            .I3(n51855), .O(n17271[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_14 (.CI(n51626), .I0(GND_net), .I1(counter[12]), 
            .CO(n51627));
    SB_LUT4 unary_minus_14_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[21]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Kp[12] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4488));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i181_2_lut (.I0(\Ki[3] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4487));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i122_2_lut (.I0(\Ki[2] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_19_lut (.I0(GND_net), .I1(n12072[16]), .I2(GND_net), 
            .I3(n51100), .O(n258[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6142_18_lut (.I0(GND_net), .I1(n15656[15]), .I2(GND_net), 
            .I3(n50914), .O(n14897[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_14_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[22]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6142_18 (.CI(n50914), .I0(n15656[15]), .I1(GND_net), 
            .CO(n50915));
    SB_LUT4 mult_18_i447_2_lut (.I0(\Ki[9] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i230_2_lut (.I0(\Ki[4] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4485));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1221_19 (.CI(n51100), .I0(n12072[16]), .I1(GND_net), 
            .CO(n51101));
    SB_LUT4 add_6142_17_lut (.I0(GND_net), .I1(n15656[14]), .I2(GND_net), 
            .I3(n50913), .O(n14897[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_17 (.CI(n50913), .I0(n15656[14]), .I1(GND_net), 
            .CO(n50914));
    SB_LUT4 mult_18_i171_2_lut (.I0(\Ki[3] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4483));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_14_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n51[23]));   // verilog/motorControl.v(53[26:40])
    defparam unary_minus_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i279_2_lut (.I0(\Ki[5] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4482));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_18_lut (.I0(GND_net), .I1(n12072[15]), .I2(GND_net), 
            .I3(n51099), .O(n258[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Kp[13] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4481));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i328_2_lut (.I0(\Ki[6] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4480));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6142_16_lut (.I0(GND_net), .I1(n15656[13]), .I2(n1108_adj_4562), 
            .I3(n50912), .O(n14897[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Kp[14] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4479));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6142_16 (.CI(n50912), .I0(n15656[13]), .I1(n1108_adj_4562), 
            .CO(n50913));
    SB_LUT4 mux_15_i17_3_lut (.I0(n48[16]), .I1(n49[16]), .I2(n182), .I3(GND_net), 
            .O(n208[16]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i17_3_lut (.I0(n208[16]), .I1(IntegralLimit[16]), .I2(n156), 
            .I3(GND_net), .O(n233[16]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_17_add_1221_18 (.CI(n51099), .I0(n12072[15]), .I1(GND_net), 
            .CO(n51100));
    SB_LUT4 add_6142_15_lut (.I0(GND_net), .I1(n15656[12]), .I2(n1035_adj_4555), 
            .I3(n50911), .O(n14897[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_15 (.CI(n50911), .I0(n15656[12]), .I1(n1035_adj_4555), 
            .CO(n50912));
    SB_LUT4 mult_18_i377_2_lut (.I0(\Ki[7] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4478));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_17_lut (.I0(GND_net), .I1(n12072[14]), .I2(GND_net), 
            .I3(n51098), .O(n258[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i496_2_lut (.I0(\Ki[10] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6142_14_lut (.I0(GND_net), .I1(n15656[11]), .I2(n962_adj_4554), 
            .I3(n50910), .O(n14897[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_14 (.CI(n50910), .I0(n15656[11]), .I1(n962_adj_4554), 
            .CO(n50911));
    SB_LUT4 mult_17_i741_2_lut (.I0(\Kp[15] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4477));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1221_17 (.CI(n51098), .I0(n12072[14]), .I1(GND_net), 
            .CO(n51099));
    SB_LUT4 add_6142_13_lut (.I0(GND_net), .I1(n15656[10]), .I2(n889_adj_4553), 
            .I3(n50909), .O(n14897[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_13 (.CI(n50909), .I0(n15656[10]), .I1(n889_adj_4553), 
            .CO(n50910));
    SB_LUT4 counter_1944_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n51625), .O(n52[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Kp[1] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Kp[0] ), .I1(n105[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i38_3_lut_3_lut (.I0(n433[19]), .I1(n353[19]), .I2(n433[18]), 
            .I3(GND_net), .O(n38_adj_4699));
    defparam LessThan_26_i38_3_lut_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 mult_18_i220_2_lut (.I0(\Ki[4] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[20]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6142_12_lut (.I0(GND_net), .I1(n15656[9]), .I2(n816_adj_4550), 
            .I3(n50908), .O(n14897[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51490_3_lut_4_lut (.I0(n433[19]), .I1(n353[19]), .I2(n433[18]), 
            .I3(n353[18]), .O(n67216));
    defparam i51490_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_6265_13 (.CI(n51855), .I0(n17779[10]), .I1(n898_adj_4590), 
            .CO(n51856));
    SB_LUT4 mult_17_add_1221_16_lut (.I0(GND_net), .I1(n12072[13]), .I2(n1096), 
            .I3(n51097), .O(n258[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6265_12_lut (.I0(GND_net), .I1(n17779[9]), .I2(n825_adj_4549), 
            .I3(n51854), .O(n17271[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_12 (.CI(n50908), .I0(n15656[9]), .I1(n816_adj_4550), 
            .CO(n50909));
    SB_LUT4 mult_18_i112_2_lut (.I0(\Ki[2] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4748));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6265_12 (.CI(n51854), .I0(n17779[9]), .I1(n825_adj_4549), 
            .CO(n51855));
    SB_CARRY mult_17_add_1221_16 (.CI(n51097), .I0(n12072[13]), .I1(n1096), 
            .CO(n51098));
    SB_LUT4 add_6265_11_lut (.I0(GND_net), .I1(n17779[8]), .I2(n752_adj_4548), 
            .I3(n51853), .O(n17271[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6142_11_lut (.I0(GND_net), .I1(n15656[8]), .I2(n743_adj_4533), 
            .I3(n50907), .O(n14897[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28972_1_lut (.I0(n353[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n42898));   // verilog/motorControl.v(55[22:42])
    defparam i28972_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6142_11 (.CI(n50907), .I0(n15656[8]), .I1(n743_adj_4533), 
            .CO(n50908));
    SB_LUT4 unary_minus_21_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[0]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i269_2_lut (.I0(\Ki[5] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4473));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i545_2_lut (.I0(\Ki[11] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_24_i42_3_lut_3_lut (.I0(PWMLimit[21]), .I1(n353[21]), 
            .I2(n353[20]), .I3(GND_net), .O(n42));   // verilog/motorControl.v(57[18:33])
    defparam LessThan_24_i42_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_DFFER result_i23 (.Q(duty[23]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[23]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i22 (.Q(duty[22]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[22]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i21 (.Q(duty[21]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[21]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i20 (.Q(duty[20]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[20]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i19 (.Q(duty[19]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[19]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i18 (.Q(duty[18]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[18]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i17 (.Q(duty[17]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[17]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i16 (.Q(duty[16]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[16]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i15 (.Q(duty[15]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[15]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i14 (.Q(duty[14]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[14]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i13 (.Q(duty[13]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[13]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i12 (.Q(duty[12]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[12]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i11 (.Q(duty[11]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[11]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i10 (.Q(duty[10]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[10]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i9 (.Q(duty[9]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[9]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i8 (.Q(duty[8]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[8]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i7 (.Q(duty[7]), .C(clk16MHz), .E(n27916), .D(\duty_23__N_3602[7] ), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i6 (.Q(duty[6]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[6]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i5 (.Q(duty[5]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[5]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i4 (.Q(duty[4]), .C(clk16MHz), .E(n27916), .D(\duty_23__N_3602[4] ), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i3 (.Q(duty[3]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[3]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i2 (.Q(duty[2]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[2]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_DFFER result_i1 (.Q(duty[1]), .C(clk16MHz), .E(n27916), .D(duty_23__N_3602[1]), 
            .R(reset));   // verilog/motorControl.v(42[14] 67[8])
    SB_CARRY add_6265_11 (.CI(n51853), .I0(n17779[8]), .I1(n752_adj_4548), 
            .CO(n51854));
    SB_LUT4 add_6265_10_lut (.I0(GND_net), .I1(n17779[7]), .I2(n679), 
            .I3(n51852), .O(n17271[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_10 (.CI(n51852), .I0(n17779[7]), .I1(n679), .CO(n51853));
    SB_LUT4 add_6142_10_lut (.I0(GND_net), .I1(n15656[7]), .I2(n670), 
            .I3(n50906), .O(n14897[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6265_9_lut (.I0(GND_net), .I1(n17779[6]), .I2(n606), .I3(n51851), 
            .O(n17271[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51516_3_lut_4_lut (.I0(PWMLimit[21]), .I1(n353[21]), .I2(n353[20]), 
            .I3(PWMLimit[20]), .O(n67242));   // verilog/motorControl.v(57[18:33])
    defparam i51516_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Kp[2] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i594_2_lut (.I0(\Ki[12] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i594_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6265_9 (.CI(n51851), .I0(n17779[6]), .I1(n606), .CO(n51852));
    SB_LUT4 add_6265_8_lut (.I0(GND_net), .I1(n17779[5]), .I2(n533), .I3(n51850), 
            .O(n17271[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i643_2_lut (.I0(\Ki[13] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i318_2_lut (.I0(\Ki[6] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4470));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[1]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Kp[3] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_15_lut (.I0(GND_net), .I1(n12072[12]), .I2(n1023), 
            .I3(n51096), .O(n258[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_8 (.CI(n51850), .I0(n17779[5]), .I1(n533), .CO(n51851));
    SB_LUT4 add_6265_7_lut (.I0(GND_net), .I1(n17779[4]), .I2(n460), .I3(n51849), 
            .O(n17271[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_13 (.CI(n51625), .I0(GND_net), .I1(counter[11]), 
            .CO(n51626));
    SB_CARRY add_6142_10 (.CI(n50906), .I0(n15656[7]), .I1(n670), .CO(n50907));
    SB_LUT4 add_6142_9_lut (.I0(GND_net), .I1(n15656[6]), .I2(n597), .I3(n50905), 
            .O(n14897[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i367_2_lut (.I0(\Ki[7] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[2]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Kp[4] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4467));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Kp[5] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4466));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1221_15 (.CI(n51096), .I0(n12072[12]), .I1(n1023), 
            .CO(n51097));
    SB_CARRY add_6142_9 (.CI(n50905), .I0(n15656[6]), .I1(n597), .CO(n50906));
    SB_LUT4 unary_minus_21_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[3]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6142_8_lut (.I0(GND_net), .I1(n15656[5]), .I2(n524), .I3(n50904), 
            .O(n14897[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_7 (.CI(n51849), .I0(n17779[4]), .I1(n460), .CO(n51850));
    SB_LUT4 add_6265_6_lut (.I0(GND_net), .I1(n17779[3]), .I2(n387), .I3(n51848), 
            .O(n17271[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1221_14_lut (.I0(GND_net), .I1(n12072[11]), .I2(n950), 
            .I3(n51095), .O(n258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_8 (.CI(n50904), .I0(n15656[5]), .I1(n524), .CO(n50905));
    SB_LUT4 add_6142_7_lut (.I0(GND_net), .I1(n15656[4]), .I2(n451), .I3(n50903), 
            .O(n14897[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_6 (.CI(n51848), .I0(n17779[3]), .I1(n387), .CO(n51849));
    SB_LUT4 mult_18_i692_2_lut (.I0(\Ki[14] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i692_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6142_7 (.CI(n50903), .I0(n15656[4]), .I1(n451), .CO(n50904));
    SB_LUT4 mult_17_i310_2_lut (.I0(\Kp[6] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4465));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1944_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n51624), .O(n52[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6265_5_lut (.I0(GND_net), .I1(n17779[2]), .I2(n314), .I3(n51847), 
            .O(n17271[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i741_2_lut (.I0(\Ki[15] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Kp[7] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4464));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i416_2_lut (.I0(\Ki[8] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i465_2_lut (.I0(\Ki[9] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6265_5 (.CI(n51847), .I0(n17779[2]), .I1(n314), .CO(n51848));
    SB_CARRY mult_17_add_1221_14 (.CI(n51095), .I0(n12072[11]), .I1(n950), 
            .CO(n51096));
    SB_LUT4 add_6142_6_lut (.I0(GND_net), .I1(n15656[3]), .I2(n378_adj_4764), 
            .I3(n50902), .O(n14897[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1221_13_lut (.I0(GND_net), .I1(n12072[10]), .I2(n877), 
            .I3(n51094), .O(n258[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Kp[8] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4463));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i514_2_lut (.I0(\Ki[10] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[4]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6142_6 (.CI(n50902), .I0(n15656[3]), .I1(n378_adj_4764), 
            .CO(n50903));
    SB_LUT4 add_6142_5_lut (.I0(GND_net), .I1(n15656[2]), .I2(n305_adj_4765), 
            .I3(n50901), .O(n14897[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_5 (.CI(n50901), .I0(n15656[2]), .I1(n305_adj_4765), 
            .CO(n50902));
    SB_LUT4 add_6142_4_lut (.I0(GND_net), .I1(n15656[1]), .I2(n232_adj_4766), 
            .I3(n50900), .O(n14897[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_4 (.CI(n50900), .I0(n15656[1]), .I1(n232_adj_4766), 
            .CO(n50901));
    SB_CARRY mult_17_add_1221_13 (.CI(n51094), .I0(n12072[10]), .I1(n877), 
            .CO(n51095));
    SB_LUT4 mult_17_add_1221_12_lut (.I0(GND_net), .I1(n12072[9]), .I2(n804), 
            .I3(n51093), .O(n258[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6142_3_lut (.I0(GND_net), .I1(n15656[0]), .I2(n159_adj_4767), 
            .I3(n50899), .O(n14897[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_3 (.CI(n50899), .I0(n15656[0]), .I1(n159_adj_4767), 
            .CO(n50900));
    SB_CARRY mult_17_add_1221_12 (.CI(n51093), .I0(n12072[9]), .I1(n804), 
            .CO(n51094));
    SB_LUT4 mult_17_add_1221_11_lut (.I0(GND_net), .I1(n12072[8]), .I2(n731), 
            .I3(n51092), .O(n258[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_11 (.CI(n51092), .I0(n12072[8]), .I1(n731), 
            .CO(n51093));
    SB_LUT4 mult_17_add_1221_10_lut (.I0(GND_net), .I1(n12072[7]), .I2(n658), 
            .I3(n51091), .O(n258[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6142_2_lut (.I0(GND_net), .I1(n17_adj_4768), .I2(n86_adj_4769), 
            .I3(GND_net), .O(n14897[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6142_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6142_2 (.CI(GND_net), .I0(n17_adj_4768), .I1(n86_adj_4769), 
            .CO(n50899));
    SB_CARRY mult_17_add_1221_10 (.CI(n51091), .I0(n12072[7]), .I1(n658), 
            .CO(n51092));
    SB_LUT4 mult_17_add_1221_9_lut (.I0(GND_net), .I1(n12072[6]), .I2(n585), 
            .I3(n51090), .O(n258[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_9 (.CI(n51090), .I0(n12072[6]), .I1(n585), 
            .CO(n51091));
    SB_LUT4 mult_17_i457_2_lut (.I0(\Kp[9] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4462));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_12 (.CI(n51624), .I0(GND_net), .I1(counter[10]), 
            .CO(n51625));
    SB_LUT4 mult_17_i506_2_lut (.I0(\Kp[10] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1221_8_lut (.I0(GND_net), .I1(n12072[5]), .I2(n512), 
            .I3(n51089), .O(n258[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_8 (.CI(n51089), .I0(n12072[5]), .I1(n512), 
            .CO(n51090));
    SB_LUT4 mult_17_add_1221_7_lut (.I0(GND_net), .I1(n12072[4]), .I2(n439_adj_4771), 
            .I3(n51088), .O(n258[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6265_4_lut (.I0(GND_net), .I1(n17779[1]), .I2(n241_adj_4772), 
            .I3(n51846), .O(n17271[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_4 (.CI(n51846), .I0(n17779[1]), .I1(n241_adj_4772), 
            .CO(n51847));
    SB_LUT4 counter_1944_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n51623), .O(n52[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_7 (.CI(n51088), .I0(n12072[4]), .I1(n439_adj_4771), 
            .CO(n51089));
    SB_LUT4 mult_17_add_1221_6_lut (.I0(GND_net), .I1(n12072[3]), .I2(n366_adj_4773), 
            .I3(n51087), .O(n258[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_6 (.CI(n51087), .I0(n12072[3]), .I1(n366_adj_4773), 
            .CO(n51088));
    SB_LUT4 add_6265_3_lut (.I0(GND_net), .I1(n17779[0]), .I2(n168_adj_4774), 
            .I3(n51845), .O(n17271[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1221_5_lut (.I0(GND_net), .I1(n12072[2]), .I2(n293_adj_4775), 
            .I3(n51086), .O(n258[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_3 (.CI(n51845), .I0(n17779[0]), .I1(n168_adj_4774), 
            .CO(n51846));
    SB_CARRY mult_17_add_1221_5 (.CI(n51086), .I0(n12072[2]), .I1(n293_adj_4775), 
            .CO(n51087));
    SB_LUT4 mult_17_add_1221_4_lut (.I0(GND_net), .I1(n12072[1]), .I2(n220_adj_4776), 
            .I3(n51085), .O(n258[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6265_2_lut (.I0(GND_net), .I1(n26_adj_4777), .I2(n95_adj_4778), 
            .I3(GND_net), .O(n17271[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6265_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_4 (.CI(n51085), .I0(n12072[1]), .I1(n220_adj_4776), 
            .CO(n51086));
    SB_LUT4 mult_17_add_1221_3_lut (.I0(GND_net), .I1(n12072[0]), .I2(n147_adj_4779), 
            .I3(n51084), .O(n258[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6265_2 (.CI(GND_net), .I0(n26_adj_4777), .I1(n95_adj_4778), 
            .CO(n51845));
    SB_LUT4 add_6295_16_lut (.I0(GND_net), .I1(n18225[13]), .I2(n1120_adj_4780), 
            .I3(n51844), .O(n17779[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_3 (.CI(n51084), .I0(n12072[0]), .I1(n147_adj_4779), 
            .CO(n51085));
    SB_LUT4 mult_17_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_4781), .I2(n74), 
            .I3(GND_net), .O(n258[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1221_2 (.CI(GND_net), .I0(n5_adj_4781), .I1(n74), 
            .CO(n51084));
    SB_LUT4 add_6295_15_lut (.I0(GND_net), .I1(n18225[12]), .I2(n1047_adj_4782), 
            .I3(n51843), .O(n17779[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_15 (.CI(n51843), .I0(n18225[12]), .I1(n1047_adj_4782), 
            .CO(n51844));
    SB_LUT4 add_6179_19_lut (.I0(GND_net), .I1(n16339[16]), .I2(GND_net), 
            .I3(n50878), .O(n15656[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6179_18_lut (.I0(GND_net), .I1(n16339[15]), .I2(GND_net), 
            .I3(n50877), .O(n15656[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_18 (.CI(n50877), .I0(n16339[15]), .I1(GND_net), 
            .CO(n50878));
    SB_LUT4 add_6179_17_lut (.I0(GND_net), .I1(n16339[14]), .I2(GND_net), 
            .I3(n50876), .O(n15656[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Kp[1] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4783));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6179_17 (.CI(n50876), .I0(n16339[14]), .I1(GND_net), 
            .CO(n50877));
    SB_LUT4 add_6179_16_lut (.I0(GND_net), .I1(n16339[13]), .I2(n1111_adj_4784), 
            .I3(n50875), .O(n15656[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_16 (.CI(n50875), .I0(n16339[13]), .I1(n1111_adj_4784), 
            .CO(n50876));
    SB_LUT4 add_6295_14_lut (.I0(GND_net), .I1(n18225[11]), .I2(n974_adj_4785), 
            .I3(n51842), .O(n17779[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_11 (.CI(n51623), .I0(GND_net), .I1(counter[9]), 
            .CO(n51624));
    SB_LUT4 add_6179_15_lut (.I0(GND_net), .I1(n16339[12]), .I2(n1038_adj_4786), 
            .I3(n50874), .O(n15656[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Kp[0] ), .I1(n105[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4787));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6179_15 (.CI(n50874), .I0(n16339[12]), .I1(n1038_adj_4786), 
            .CO(n50875));
    SB_LUT4 add_6179_14_lut (.I0(GND_net), .I1(n16339[11]), .I2(n965_adj_4788), 
            .I3(n50873), .O(n15656[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_14 (.CI(n50873), .I0(n16339[11]), .I1(n965_adj_4788), 
            .CO(n50874));
    SB_LUT4 counter_1944_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n51622), .O(n52[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6179_13_lut (.I0(GND_net), .I1(n16339[10]), .I2(n892_adj_4789), 
            .I3(n50872), .O(n15656[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_13 (.CI(n50872), .I0(n16339[10]), .I1(n892_adj_4789), 
            .CO(n50873));
    SB_CARRY counter_1944_add_4_10 (.CI(n51622), .I0(GND_net), .I1(counter[8]), 
            .CO(n51623));
    SB_LUT4 add_6179_12_lut (.I0(GND_net), .I1(n16339[9]), .I2(n819_adj_4790), 
            .I3(n50871), .O(n15656[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_12 (.CI(n50871), .I0(n16339[9]), .I1(n819_adj_4790), 
            .CO(n50872));
    SB_LUT4 add_6179_11_lut (.I0(GND_net), .I1(n16339[8]), .I2(n746_adj_4791), 
            .I3(n50870), .O(n15656[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_11 (.CI(n50870), .I0(n16339[8]), .I1(n746_adj_4791), 
            .CO(n50871));
    SB_LUT4 add_6179_10_lut (.I0(GND_net), .I1(n16339[7]), .I2(n673_adj_4792), 
            .I3(n50869), .O(n15656[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_10 (.CI(n50869), .I0(n16339[7]), .I1(n673_adj_4792), 
            .CO(n50870));
    SB_LUT4 add_6179_9_lut (.I0(GND_net), .I1(n16339[6]), .I2(n600_adj_4793), 
            .I3(n50868), .O(n15656[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_14 (.CI(n51842), .I0(n18225[11]), .I1(n974_adj_4785), 
            .CO(n51843));
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n54[23]), 
            .I3(n50524), .O(n433[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n54[22]), 
            .I3(n50523), .O(n433[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_9 (.CI(n50868), .I0(n16339[6]), .I1(n600_adj_4793), 
            .CO(n50869));
    SB_LUT4 add_6179_8_lut (.I0(GND_net), .I1(n16339[5]), .I2(n527_adj_4796), 
            .I3(n50867), .O(n15656[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_8 (.CI(n50867), .I0(n16339[5]), .I1(n527_adj_4796), 
            .CO(n50868));
    SB_LUT4 add_6295_13_lut (.I0(GND_net), .I1(n18225[10]), .I2(n901_adj_4797), 
            .I3(n51841), .O(n17779[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6179_7_lut (.I0(GND_net), .I1(n16339[4]), .I2(n454_adj_4798), 
            .I3(n50866), .O(n15656[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_13 (.CI(n51841), .I0(n18225[10]), .I1(n901_adj_4797), 
            .CO(n51842));
    SB_LUT4 counter_1944_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n51621), .O(n52[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_7 (.CI(n50866), .I0(n16339[4]), .I1(n454_adj_4798), 
            .CO(n50867));
    SB_LUT4 add_6179_6_lut (.I0(GND_net), .I1(n16339[3]), .I2(n381_adj_4799), 
            .I3(n50865), .O(n15656[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6295_12_lut (.I0(GND_net), .I1(n18225[9]), .I2(n828_adj_4800), 
            .I3(n51840), .O(n17779[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_24 (.CI(n50523), .I0(GND_net), .I1(n54[22]), 
            .CO(n50524));
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n54[21]), 
            .I3(n50522), .O(n433[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_9 (.CI(n51621), .I0(GND_net), .I1(counter[7]), 
            .CO(n51622));
    SB_LUT4 add_19_25_lut (.I0(GND_net), .I1(n11613[0]), .I2(n12188[0]), 
            .I3(n50408), .O(n353[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n50522), .I0(GND_net), .I1(n54[21]), 
            .CO(n50523));
    SB_LUT4 add_19_24_lut (.I0(GND_net), .I1(n258[22]), .I2(n303[22]), 
            .I3(n50407), .O(n353[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n54[20]), 
            .I3(n50521), .O(n433[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n51620), .O(n52[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_6 (.CI(n50865), .I0(n16339[3]), .I1(n381_adj_4799), 
            .CO(n50866));
    SB_LUT4 add_6179_5_lut (.I0(GND_net), .I1(n16339[2]), .I2(n308_adj_4804), 
            .I3(n50864), .O(n15656[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_12 (.CI(n51840), .I0(n18225[9]), .I1(n828_adj_4800), 
            .CO(n51841));
    SB_LUT4 add_6295_11_lut (.I0(GND_net), .I1(n18225[8]), .I2(n755_adj_4805), 
            .I3(n51839), .O(n17779[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_5 (.CI(n50864), .I0(n16339[2]), .I1(n308_adj_4804), 
            .CO(n50865));
    SB_LUT4 add_6179_4_lut (.I0(GND_net), .I1(n16339[1]), .I2(n235_adj_4806), 
            .I3(n50863), .O(n15656[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_8 (.CI(n51620), .I0(GND_net), .I1(counter[6]), 
            .CO(n51621));
    SB_CARRY add_19_24 (.CI(n50407), .I0(n258[22]), .I1(n303[22]), .CO(n50408));
    SB_CARRY add_6179_4 (.CI(n50863), .I0(n16339[1]), .I1(n235_adj_4806), 
            .CO(n50864));
    SB_LUT4 add_6179_3_lut (.I0(GND_net), .I1(n16339[0]), .I2(n162_adj_4807), 
            .I3(n50862), .O(n15656[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_3 (.CI(n50862), .I0(n16339[0]), .I1(n162_adj_4807), 
            .CO(n50863));
    SB_LUT4 add_6179_2_lut (.I0(GND_net), .I1(n20_adj_4808), .I2(n89_adj_4809), 
            .I3(GND_net), .O(n15656[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6179_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_19_23_lut (.I0(GND_net), .I1(n258[21]), .I2(n303[21]), 
            .I3(n50406), .O(n353[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6179_2 (.CI(GND_net), .I0(n20_adj_4808), .I1(n89_adj_4809), 
            .CO(n50862));
    SB_LUT4 add_6449_9_lut (.I0(GND_net), .I1(n19947[6]), .I2(n630), .I3(n50861), 
            .O(n19823[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_8_lut (.I0(GND_net), .I1(n19947[5]), .I2(n557), .I3(n50860), 
            .O(n19823[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_8 (.CI(n50860), .I0(n19947[5]), .I1(n557), .CO(n50861));
    SB_LUT4 add_6449_7_lut (.I0(GND_net), .I1(n19947[4]), .I2(n484_adj_4810), 
            .I3(n50859), .O(n19823[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_11 (.CI(n51839), .I0(n18225[8]), .I1(n755_adj_4805), 
            .CO(n51840));
    SB_LUT4 counter_1944_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n51619), .O(n52[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_7 (.CI(n51619), .I0(GND_net), .I1(counter[5]), 
            .CO(n51620));
    SB_CARRY add_19_23 (.CI(n50406), .I0(n258[21]), .I1(n303[21]), .CO(n50407));
    SB_CARRY unary_minus_27_add_3_22 (.CI(n50521), .I0(GND_net), .I1(n54[20]), 
            .CO(n50522));
    SB_LUT4 add_19_22_lut (.I0(GND_net), .I1(n258[20]), .I2(n303[20]), 
            .I3(n50405), .O(n353[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n54[19]), 
            .I3(n50520), .O(n433[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_22 (.CI(n50405), .I0(n258[20]), .I1(n303[20]), .CO(n50406));
    SB_LUT4 add_19_21_lut (.I0(GND_net), .I1(n258[19]), .I2(n303[19]), 
            .I3(n50404), .O(n353[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_7 (.CI(n50859), .I0(n19947[4]), .I1(n484_adj_4810), 
            .CO(n50860));
    SB_LUT4 add_6295_10_lut (.I0(GND_net), .I1(n18225[7]), .I2(n682_adj_4813), 
            .I3(n51838), .O(n17779[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_6_lut (.I0(GND_net), .I1(n19947[3]), .I2(n411), .I3(n50858), 
            .O(n19823[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_10 (.CI(n51838), .I0(n18225[7]), .I1(n682_adj_4813), 
            .CO(n51839));
    SB_CARRY add_6449_6 (.CI(n50858), .I0(n19947[3]), .I1(n411), .CO(n50859));
    SB_CARRY unary_minus_27_add_3_21 (.CI(n50520), .I0(GND_net), .I1(n54[19]), 
            .CO(n50521));
    SB_LUT4 add_6449_5_lut (.I0(GND_net), .I1(n19947[2]), .I2(n338), .I3(n50857), 
            .O(n19823[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_21 (.CI(n50404), .I0(n258[19]), .I1(n303[19]), .CO(n50405));
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n54[18]), 
            .I3(n50519), .O(n433[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_5 (.CI(n50857), .I0(n19947[2]), .I1(n338), .CO(n50858));
    SB_LUT4 add_6449_4_lut (.I0(GND_net), .I1(n19947[1]), .I2(n265), .I3(n50856), 
            .O(n19823[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_4 (.CI(n50856), .I0(n19947[1]), .I1(n265), .CO(n50857));
    SB_LUT4 add_6295_9_lut (.I0(GND_net), .I1(n18225[6]), .I2(n609_adj_4815), 
            .I3(n51837), .O(n17779[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n51618), .O(n52[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_6 (.CI(n51618), .I0(GND_net), .I1(counter[4]), 
            .CO(n51619));
    SB_LUT4 add_19_20_lut (.I0(GND_net), .I1(n258[18]), .I2(n303[18]), 
            .I3(n50403), .O(n353[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_3_lut (.I0(GND_net), .I1(n19947[0]), .I2(n192_adj_4816), 
            .I3(n50855), .O(n19823[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_20 (.CI(n50403), .I0(n258[18]), .I1(n303[18]), .CO(n50404));
    SB_CARRY add_6449_3 (.CI(n50855), .I0(n19947[0]), .I1(n192_adj_4816), 
            .CO(n50856));
    SB_CARRY unary_minus_27_add_3_20 (.CI(n50519), .I0(GND_net), .I1(n54[18]), 
            .CO(n50520));
    SB_LUT4 add_6449_2_lut (.I0(GND_net), .I1(n50), .I2(n119_adj_4817), 
            .I3(GND_net), .O(n19823[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_19_19_lut (.I0(GND_net), .I1(n258[17]), .I2(n303[17]), 
            .I3(n50402), .O(n353[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n54[17]), 
            .I3(n50518), .O(n433[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_19 (.CI(n50402), .I0(n258[17]), .I1(n303[17]), .CO(n50403));
    SB_CARRY unary_minus_27_add_3_19 (.CI(n50518), .I0(GND_net), .I1(n54[17]), 
            .CO(n50519));
    SB_LUT4 mult_17_i555_2_lut (.I0(\Kp[11] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6295_9 (.CI(n51837), .I0(n18225[6]), .I1(n609_adj_4815), 
            .CO(n51838));
    SB_LUT4 mult_17_i604_2_lut (.I0(\Kp[12] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_19_18_lut (.I0(GND_net), .I1(n258[16]), .I2(n303[16]), 
            .I3(n50401), .O(n353[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n54[16]), 
            .I3(n50517), .O(n433[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_18 (.CI(n50401), .I0(n258[16]), .I1(n303[16]), .CO(n50402));
    SB_LUT4 add_19_17_lut (.I0(GND_net), .I1(n258[15]), .I2(n303[15]), 
            .I3(n50400), .O(n353[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_2 (.CI(GND_net), .I0(n50), .I1(n119_adj_4817), .CO(n50855));
    SB_CARRY add_19_17 (.CI(n50400), .I0(n258[15]), .I1(n303[15]), .CO(n50401));
    SB_LUT4 add_19_16_lut (.I0(GND_net), .I1(n258[14]), .I2(n303[14]), 
            .I3(n50399), .O(n353[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i563_2_lut (.I0(\Ki[11] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1944_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n51617), .O(n52[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_16 (.CI(n50399), .I0(n258[14]), .I1(n303[14]), .CO(n50400));
    SB_CARRY unary_minus_27_add_3_18 (.CI(n50517), .I0(GND_net), .I1(n54[16]), 
            .CO(n50518));
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n54[15]), 
            .I3(n50516), .O(n433[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6415_11_lut (.I0(GND_net), .I1(n19665[8]), .I2(n770_adj_4822), 
            .I3(n51059), .O(n19469[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_17 (.CI(n50516), .I0(GND_net), .I1(n54[15]), 
            .CO(n50517));
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n54[14]), 
            .I3(n50515), .O(n433[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6415_10_lut (.I0(GND_net), .I1(n19665[7]), .I2(n697_adj_4824), 
            .I3(n51058), .O(n19469[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6295_8_lut (.I0(GND_net), .I1(n18225[5]), .I2(n536_adj_4825), 
            .I3(n51836), .O(n17779[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_5 (.CI(n51617), .I0(GND_net), .I1(counter[3]), 
            .CO(n51618));
    SB_CARRY add_6295_8 (.CI(n51836), .I0(n18225[5]), .I1(n536_adj_4825), 
            .CO(n51837));
    SB_LUT4 add_6295_7_lut (.I0(GND_net), .I1(n18225[4]), .I2(n463_adj_4826), 
            .I3(n51835), .O(n17779[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_7 (.CI(n51835), .I0(n18225[4]), .I1(n463_adj_4826), 
            .CO(n51836));
    SB_LUT4 add_6295_6_lut (.I0(GND_net), .I1(n18225[3]), .I2(n390_adj_4827), 
            .I3(n51834), .O(n17779[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_6 (.CI(n51834), .I0(n18225[3]), .I1(n390_adj_4827), 
            .CO(n51835));
    SB_LUT4 add_6295_5_lut (.I0(GND_net), .I1(n18225[2]), .I2(n317_adj_4828), 
            .I3(n51833), .O(n17779[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i610_2_lut (.I0(\Ki[12] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4829));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6295_5 (.CI(n51833), .I0(n18225[2]), .I1(n317_adj_4828), 
            .CO(n51834));
    SB_LUT4 counter_1944_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n51616), .O(n52[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Kp[13] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6295_4_lut (.I0(GND_net), .I1(n18225[1]), .I2(n244_adj_4830), 
            .I3(n51832), .O(n17779[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Kp[14] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_4 (.CI(n51616), .I0(GND_net), .I1(counter[2]), 
            .CO(n51617));
    SB_LUT4 counter_1944_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n51615), .O(n52[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_4 (.CI(n51832), .I0(n18225[1]), .I1(n244_adj_4830), 
            .CO(n51833));
    SB_LUT4 add_6295_3_lut (.I0(GND_net), .I1(n18225[0]), .I2(n171_adj_4831), 
            .I3(n51831), .O(n17779[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_3 (.CI(n51831), .I0(n18225[0]), .I1(n171_adj_4831), 
            .CO(n51832));
    SB_LUT4 add_6295_2_lut (.I0(GND_net), .I1(n29_adj_4832), .I2(n98_adj_4833), 
            .I3(GND_net), .O(n17779[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6295_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i659_2_lut (.I0(\Ki[13] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4834));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i659_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1944_add_4_3 (.CI(n51615), .I0(GND_net), .I1(counter[1]), 
            .CO(n51616));
    SB_LUT4 unary_minus_21_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[5]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6415_10 (.CI(n51058), .I0(n19665[7]), .I1(n697_adj_4824), 
            .CO(n51059));
    SB_LUT4 add_6415_9_lut (.I0(GND_net), .I1(n19665[6]), .I2(n624), .I3(n51057), 
            .O(n19469[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1944_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n52[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1944_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6415_9 (.CI(n51057), .I0(n19665[6]), .I1(n624), .CO(n51058));
    SB_LUT4 mult_18_i612_2_lut (.I0(\Ki[12] ), .I1(n233[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_19_15_lut (.I0(GND_net), .I1(n258[13]), .I2(n303[13]), 
            .I3(n50398), .O(n353[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6415_8_lut (.I0(GND_net), .I1(n19665[5]), .I2(n551), .I3(n51056), 
            .O(n19469[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_15 (.CI(n50398), .I0(n258[13]), .I1(n303[13]), .CO(n50399));
    SB_CARRY add_6415_8 (.CI(n51056), .I0(n19665[5]), .I1(n551), .CO(n51057));
    SB_LUT4 mult_17_i751_2_lut (.I0(\Kp[15] ), .I1(n105[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Kp[9] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4838));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Kp[10] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4839));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6415_7_lut (.I0(GND_net), .I1(n19665[4]), .I2(n478_adj_1), 
            .I3(n51055), .O(n19469[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6415_7 (.CI(n51055), .I0(n19665[4]), .I1(n478_adj_1), 
            .CO(n51056));
    SB_LUT4 unary_minus_21_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[6]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_19_14_lut (.I0(GND_net), .I1(n258[12]), .I2(n303[12]), 
            .I3(n50397), .O(n353[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1944_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n51615));
    SB_CARRY unary_minus_27_add_3_16 (.CI(n50515), .I0(GND_net), .I1(n54[14]), 
            .CO(n50516));
    SB_LUT4 add_6415_6_lut (.I0(GND_net), .I1(n19665[3]), .I2(n405_adj_2), 
            .I3(n51054), .O(n19469[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6295_2 (.CI(GND_net), .I0(n29_adj_4832), .I1(n98_adj_4833), 
            .CO(n51831));
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n54[13]), 
            .I3(n50514), .O(n433[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6439_9_lut (.I0(GND_net), .I1(n19869[6]), .I2(n630_adj_4843), 
            .I3(n51830), .O(n19726[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6439_8_lut (.I0(GND_net), .I1(n19869[5]), .I2(n557_adj_4844), 
            .I3(n51829), .O(n19726[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6439_8 (.CI(n51829), .I0(n19869[5]), .I1(n557_adj_4844), 
            .CO(n51830));
    SB_LUT4 add_6439_7_lut (.I0(GND_net), .I1(n19869[4]), .I2(n484_adj_4845), 
            .I3(n51828), .O(n19726[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6439_7 (.CI(n51828), .I0(n19869[4]), .I1(n484_adj_4845), 
            .CO(n51829));
    SB_LUT4 add_6439_6_lut (.I0(GND_net), .I1(n19869[3]), .I2(n411_adj_4846), 
            .I3(n51827), .O(n19726[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_14 (.CI(n50397), .I0(n258[12]), .I1(n303[12]), .CO(n50398));
    SB_LUT4 add_19_13_lut (.I0(GND_net), .I1(n258[11]), .I2(n303[11]), 
            .I3(n50396), .O(n353[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6439_6 (.CI(n51827), .I0(n19869[3]), .I1(n411_adj_4846), 
            .CO(n51828));
    SB_CARRY add_6415_6 (.CI(n51054), .I0(n19665[3]), .I1(n405_adj_2), 
            .CO(n51055));
    SB_LUT4 add_6415_5_lut (.I0(GND_net), .I1(n19665[2]), .I2(n332), .I3(n51053), 
            .O(n19469[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6415_5 (.CI(n51053), .I0(n19665[2]), .I1(n332), .CO(n51054));
    SB_LUT4 add_6439_5_lut (.I0(GND_net), .I1(n19869[2]), .I2(n338_adj_4848), 
            .I3(n51826), .O(n19726[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i69_2_lut (.I0(\Ki[1] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4849));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i22_2_lut (.I0(\Ki[0] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4850));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Kp[1] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4459));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50886_3_lut_4_lut (.I0(n48[3]), .I1(n49[3]), .I2(n49[2]), 
            .I3(n48[2]), .O(n66612));   // verilog/motorControl.v(52[25:48])
    defparam i50886_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_6439_5 (.CI(n51826), .I0(n19869[2]), .I1(n338_adj_4848), 
            .CO(n51827));
    SB_LUT4 add_6439_4_lut (.I0(GND_net), .I1(n19869[1]), .I2(n265_adj_4851), 
            .I3(n51825), .O(n19726[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6439_4 (.CI(n51825), .I0(n19869[1]), .I1(n265_adj_4851), 
            .CO(n51826));
    SB_LUT4 add_6439_3_lut (.I0(GND_net), .I1(n19869[0]), .I2(n192_adj_4852), 
            .I3(n51824), .O(n19726[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i118_2_lut (.I0(\Ki[2] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4853));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i36_2_lut (.I0(\Kp[0] ), .I1(n105[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i36_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6439_3 (.CI(n51824), .I0(n19869[0]), .I1(n192_adj_4852), 
            .CO(n51825));
    SB_LUT4 add_6439_2_lut (.I0(GND_net), .I1(n50_adj_4854), .I2(n119_adj_4855), 
            .I3(GND_net), .O(n19726[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6439_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6439_2 (.CI(GND_net), .I0(n50_adj_4854), .I1(n119_adj_4855), 
            .CO(n51824));
    SB_LUT4 add_6415_4_lut (.I0(GND_net), .I1(n19665[1]), .I2(n259), .I3(n51052), 
            .O(n19469[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_15 (.CI(n50514), .I0(GND_net), .I1(n54[13]), 
            .CO(n50515));
    SB_LUT4 mult_17_i102_2_lut (.I0(\Kp[2] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4857));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i167_2_lut (.I0(\Ki[3] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4858));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i51_2_lut (.I0(\Ki[1] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4859));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6323_15_lut (.I0(GND_net), .I1(n18613[12]), .I2(n1050_adj_4860), 
            .I3(n51823), .O(n18225[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i4_2_lut (.I0(\Ki[0] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4861));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[7]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[8]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6415_4 (.CI(n51052), .I0(n19665[1]), .I1(n259), .CO(n51053));
    SB_LUT4 add_6323_14_lut (.I0(GND_net), .I1(n18613[11]), .I2(n977_adj_4862), 
            .I3(n51822), .O(n18225[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_13_i6_3_lut_3_lut (.I0(n48[3]), .I1(n49[3]), .I2(n49[2]), 
            .I3(GND_net), .O(n6_adj_4863));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_21_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[23]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36191_2_lut_3_lut (.I0(\Kp[1] ), .I1(n105[22]), .I2(n62_c), 
            .I3(GND_net), .O(n20063[0]));   // verilog/motorControl.v(55[22:28])
    defparam i36191_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 add_6415_3_lut (.I0(GND_net), .I1(n19665[0]), .I2(n186), .I3(n51051), 
            .O(n19469[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n54[12]), 
            .I3(n50513), .O(n433[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6415_3 (.CI(n51051), .I0(n19665[0]), .I1(n186), .CO(n51052));
    SB_LUT4 add_6382_12_lut (.I0(GND_net), .I1(n19328[9]), .I2(n840_adj_4867), 
            .I3(n52019), .O(n19065[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6382_11_lut (.I0(GND_net), .I1(n19328[8]), .I2(n767_adj_4868), 
            .I3(n52018), .O(n19065[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_11 (.CI(n52018), .I0(n19328[8]), .I1(n767_adj_4868), 
            .CO(n52019));
    SB_LUT4 add_6382_10_lut (.I0(GND_net), .I1(n19328[7]), .I2(n694_adj_4869), 
            .I3(n52017), .O(n19065[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_10 (.CI(n52017), .I0(n19328[7]), .I1(n694_adj_4869), 
            .CO(n52018));
    SB_LUT4 add_6382_9_lut (.I0(GND_net), .I1(n19328[6]), .I2(n621_adj_4870), 
            .I3(n52016), .O(n19065[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_9 (.CI(n52016), .I0(n19328[6]), .I1(n621_adj_4870), 
            .CO(n52017));
    SB_LUT4 add_6382_8_lut (.I0(GND_net), .I1(n19328[5]), .I2(n548_adj_4871), 
            .I3(n52015), .O(n19065[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_8 (.CI(n52015), .I0(n19328[5]), .I1(n548_adj_4871), 
            .CO(n52016));
    SB_LUT4 add_6382_7_lut (.I0(GND_net), .I1(n19328[4]), .I2(n475_adj_4872), 
            .I3(n52014), .O(n19065[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6415_2_lut (.I0(GND_net), .I1(n44_adj_4873), .I2(n113), 
            .I3(GND_net), .O(n19469[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6415_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_7 (.CI(n52014), .I0(n19328[4]), .I1(n475_adj_4872), 
            .CO(n52015));
    SB_LUT4 add_6382_6_lut (.I0(GND_net), .I1(n19328[3]), .I2(n402_adj_4875), 
            .I3(n52013), .O(n19065[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_6 (.CI(n52013), .I0(n19328[3]), .I1(n402_adj_4875), 
            .CO(n52014));
    SB_LUT4 mult_18_i100_2_lut (.I0(\Ki[2] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4876));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6382_5_lut (.I0(GND_net), .I1(n19328[2]), .I2(n329_adj_4877), 
            .I3(n52012), .O(n19065[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[0]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n50513), .I0(GND_net), .I1(n54[12]), 
            .CO(n50514));
    SB_CARRY add_6323_14 (.CI(n51822), .I0(n18613[11]), .I1(n977_adj_4862), 
            .CO(n51823));
    SB_CARRY add_6382_5 (.CI(n52012), .I0(n19328[2]), .I1(n329_adj_4877), 
            .CO(n52013));
    SB_LUT4 add_6382_4_lut (.I0(GND_net), .I1(n19328[1]), .I2(n256_adj_4879), 
            .I3(n52011), .O(n19065[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_13_lut (.I0(GND_net), .I1(n18613[10]), .I2(n904_adj_4880), 
            .I3(n51821), .O(n18225[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_4 (.CI(n52011), .I0(n19328[1]), .I1(n256_adj_4879), 
            .CO(n52012));
    SB_LUT4 add_6382_3_lut (.I0(GND_net), .I1(n19328[0]), .I2(n183_adj_4881), 
            .I3(n52010), .O(n19065[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_3 (.CI(n52010), .I0(n19328[0]), .I1(n183_adj_4881), 
            .CO(n52011));
    SB_LUT4 add_6382_2_lut (.I0(GND_net), .I1(n41_adj_4882), .I2(n110_adj_4883), 
            .I3(GND_net), .O(n19065[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6382_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6382_2 (.CI(GND_net), .I0(n41_adj_4882), .I1(n110_adj_4883), 
            .CO(n52010));
    SB_LUT4 mult_18_add_1225_24_lut (.I0(n233[23]), .I1(n12695[21]), .I2(GND_net), 
            .I3(n52009), .O(n12188[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6415_2 (.CI(GND_net), .I0(n44_adj_4873), .I1(n113), .CO(n51051));
    SB_LUT4 add_5992_23_lut (.I0(GND_net), .I1(n13134[20]), .I2(GND_net), 
            .I3(n51050), .O(n12072[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_22_lut (.I0(GND_net), .I1(n13134[19]), .I2(GND_net), 
            .I3(n51049), .O(n12072[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_22 (.CI(n51049), .I0(n13134[19]), .I1(GND_net), 
            .CO(n51050));
    SB_LUT4 add_5992_21_lut (.I0(GND_net), .I1(n13134[18]), .I2(GND_net), 
            .I3(n51048), .O(n12072[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_13 (.CI(n51821), .I0(n18613[10]), .I1(n904_adj_4880), 
            .CO(n51822));
    SB_LUT4 add_6323_12_lut (.I0(GND_net), .I1(n18613[9]), .I2(n831_adj_4884), 
            .I3(n51820), .O(n18225[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_add_1225_23_lut (.I0(GND_net), .I1(n12695[20]), .I2(GND_net), 
            .I3(n52008), .O(n303[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Kp[3] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4885));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[1]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i149_2_lut (.I0(\Ki[3] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4887));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5992_21 (.CI(n51048), .I0(n13134[18]), .I1(GND_net), 
            .CO(n51049));
    SB_CARRY mult_18_add_1225_23 (.CI(n52008), .I0(n12695[20]), .I1(GND_net), 
            .CO(n52009));
    SB_LUT4 mult_18_add_1225_22_lut (.I0(GND_net), .I1(n12695[19]), .I2(GND_net), 
            .I3(n52007), .O(n303[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_20_lut (.I0(GND_net), .I1(n13134[17]), .I2(GND_net), 
            .I3(n51047), .O(n12072[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_22 (.CI(n52007), .I0(n12695[19]), .I1(GND_net), 
            .CO(n52008));
    SB_LUT4 mult_18_add_1225_21_lut (.I0(GND_net), .I1(n12695[18]), .I2(GND_net), 
            .I3(n52006), .O(n303[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_21 (.CI(n52006), .I0(n12695[18]), .I1(GND_net), 
            .CO(n52007));
    SB_LUT4 mult_18_add_1225_20_lut (.I0(GND_net), .I1(n12695[17]), .I2(GND_net), 
            .I3(n52005), .O(n303[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_20 (.CI(n52005), .I0(n12695[17]), .I1(GND_net), 
            .CO(n52006));
    SB_LUT4 mult_18_add_1225_19_lut (.I0(GND_net), .I1(n12695[16]), .I2(GND_net), 
            .I3(n52004), .O(n303[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_19 (.CI(n52004), .I0(n12695[16]), .I1(GND_net), 
            .CO(n52005));
    SB_LUT4 mult_18_add_1225_18_lut (.I0(GND_net), .I1(n12695[15]), .I2(GND_net), 
            .I3(n52003), .O(n303[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_18 (.CI(n52003), .I0(n12695[15]), .I1(GND_net), 
            .CO(n52004));
    SB_LUT4 mult_18_add_1225_17_lut (.I0(GND_net), .I1(n12695[14]), .I2(GND_net), 
            .I3(n52002), .O(n303[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_17 (.CI(n52002), .I0(n12695[14]), .I1(GND_net), 
            .CO(n52003));
    SB_LUT4 mult_18_add_1225_16_lut (.I0(GND_net), .I1(n12695[13]), .I2(n1096_adj_4888), 
            .I3(n52001), .O(n303[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n54[11]), 
            .I3(n50512), .O(n433[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_20 (.CI(n51047), .I0(n13134[17]), .I1(GND_net), 
            .CO(n51048));
    SB_LUT4 add_5992_19_lut (.I0(GND_net), .I1(n13134[16]), .I2(GND_net), 
            .I3(n51046), .O(n12072[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[1] ), .I1(n105[22]), .I2(n62_c), .I3(n62910), 
            .O(n20063[1]));   // verilog/motorControl.v(55[22:28])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_CARRY add_5992_19 (.CI(n51046), .I0(n13134[16]), .I1(GND_net), 
            .CO(n51047));
    SB_LUT4 add_5992_18_lut (.I0(GND_net), .I1(n13134[15]), .I2(GND_net), 
            .I3(n51045), .O(n12072[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i198_2_lut (.I0(\Ki[4] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4890));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i198_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5992_18 (.CI(n51045), .I0(n13134[15]), .I1(GND_net), 
            .CO(n51046));
    SB_CARRY add_19_13 (.CI(n50396), .I0(n258[11]), .I1(n303[11]), .CO(n50397));
    SB_LUT4 add_19_12_lut (.I0(GND_net), .I1(n258[10]), .I2(n303[10]), 
            .I3(n50395), .O(n353[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_13 (.CI(n50512), .I0(GND_net), .I1(n54[11]), 
            .CO(n50513));
    SB_CARRY add_6323_12 (.CI(n51820), .I0(n18613[9]), .I1(n831_adj_4884), 
            .CO(n51821));
    SB_LUT4 add_5992_17_lut (.I0(GND_net), .I1(n13134[14]), .I2(GND_net), 
            .I3(n51044), .O(n12072[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_12 (.CI(n50395), .I0(n258[10]), .I1(n303[10]), .CO(n50396));
    SB_CARRY add_5992_17 (.CI(n51044), .I0(n13134[14]), .I1(GND_net), 
            .CO(n51045));
    SB_LUT4 add_5992_16_lut (.I0(GND_net), .I1(n13134[13]), .I2(n1099_adj_4892), 
            .I3(n51043), .O(n12072[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_11_lut (.I0(GND_net), .I1(n18613[8]), .I2(n758_adj_4893), 
            .I3(n51819), .O(n18225[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_16 (.CI(n51043), .I0(n13134[13]), .I1(n1099_adj_4892), 
            .CO(n51044));
    SB_LUT4 add_5992_15_lut (.I0(GND_net), .I1(n13134[12]), .I2(n1026_adj_4894), 
            .I3(n51042), .O(n12072[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_15 (.CI(n51042), .I0(n13134[12]), .I1(n1026_adj_4894), 
            .CO(n51043));
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n54[10]), 
            .I3(n50511), .O(n433[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_11 (.CI(n51819), .I0(n18613[8]), .I1(n758_adj_4893), 
            .CO(n51820));
    SB_LUT4 add_5992_14_lut (.I0(GND_net), .I1(n13134[11]), .I2(n953_adj_4896), 
            .I3(n51041), .O(n12072[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n50511), .I0(GND_net), .I1(n54[10]), 
            .CO(n50512));
    SB_LUT4 add_19_11_lut (.I0(GND_net), .I1(n258[9]), .I2(n303[9]), .I3(n50394), 
            .O(n353[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_14 (.CI(n51041), .I0(n13134[11]), .I1(n953_adj_4896), 
            .CO(n51042));
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n54[9]), 
            .I3(n50510), .O(n433[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_11 (.CI(n50394), .I0(n258[9]), .I1(n303[9]), .CO(n50395));
    SB_LUT4 add_19_10_lut (.I0(GND_net), .I1(n258[8]), .I2(n303[8]), .I3(n50393), 
            .O(n353[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_i247_2_lut (.I0(\Ki[5] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4898));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_18_add_1225_16 (.CI(n52001), .I0(n12695[13]), .I1(n1096_adj_4888), 
            .CO(n52002));
    SB_LUT4 mult_18_add_1225_15_lut (.I0(GND_net), .I1(n12695[12]), .I2(n1023_adj_4899), 
            .I3(n52000), .O(n303[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51043_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n48[3]), .I2(n48[2]), 
            .I3(IntegralLimit[2]), .O(n66769));   // verilog/motorControl.v(50[16:38])
    defparam i51043_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_19_10 (.CI(n50393), .I0(n258[8]), .I1(n303[8]), .CO(n50394));
    SB_CARRY unary_minus_27_add_3_11 (.CI(n50510), .I0(GND_net), .I1(n54[9]), 
            .CO(n50511));
    SB_LUT4 add_19_9_lut (.I0(GND_net), .I1(n258[7]), .I2(n303[7]), .I3(n50392), 
            .O(n353[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n54[8]), 
            .I3(n50509), .O(n433[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_13_lut (.I0(GND_net), .I1(n13134[10]), .I2(n880_adj_4902), 
            .I3(n51040), .O(n12072[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_10 (.CI(n50509), .I0(GND_net), .I1(n54[8]), 
            .CO(n50510));
    SB_CARRY add_19_9 (.CI(n50392), .I0(n258[7]), .I1(n303[7]), .CO(n50393));
    SB_CARRY add_5992_13 (.CI(n51040), .I0(n13134[10]), .I1(n880_adj_4902), 
            .CO(n51041));
    SB_LUT4 add_5992_12_lut (.I0(GND_net), .I1(n13134[9]), .I2(n807_adj_4903), 
            .I3(n51039), .O(n12072[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n54[7]), 
            .I3(n50508), .O(n433[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n50508), .I0(GND_net), .I1(n54[7]), 
            .CO(n50509));
    SB_LUT4 add_6214_18_lut (.I0(GND_net), .I1(n16950[15]), .I2(GND_net), 
            .I3(n50835), .O(n16339[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_19_8_lut (.I0(GND_net), .I1(n258[6]), .I2(n303[6]), .I3(n50391), 
            .O(n353[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_12 (.CI(n51039), .I0(n13134[9]), .I1(n807_adj_4903), 
            .CO(n51040));
    SB_LUT4 add_6214_17_lut (.I0(GND_net), .I1(n16950[14]), .I2(GND_net), 
            .I3(n50834), .O(n16339[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_17 (.CI(n50834), .I0(n16950[14]), .I1(GND_net), 
            .CO(n50835));
    SB_LUT4 add_5992_11_lut (.I0(GND_net), .I1(n13134[8]), .I2(n734_adj_4905), 
            .I3(n51038), .O(n12072[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_8 (.CI(n50391), .I0(n258[6]), .I1(n303[6]), .CO(n50392));
    SB_LUT4 add_19_7_lut (.I0(GND_net), .I1(n258[5]), .I2(n303[5]), .I3(n50390), 
            .O(n353[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_19_7 (.CI(n50390), .I0(n258[5]), .I1(n303[5]), .CO(n50391));
    SB_CARRY add_5992_11 (.CI(n51038), .I0(n13134[8]), .I1(n734_adj_4905), 
            .CO(n51039));
    SB_LUT4 add_5992_10_lut (.I0(GND_net), .I1(n13134[7]), .I2(n661_adj_4906), 
            .I3(n51037), .O(n12072[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6214_16_lut (.I0(GND_net), .I1(n16950[13]), .I2(n1114_adj_4907), 
            .I3(n50833), .O(n16339[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_16 (.CI(n50833), .I0(n16950[13]), .I1(n1114_adj_4907), 
            .CO(n50834));
    SB_CARRY add_5992_10 (.CI(n51037), .I0(n13134[7]), .I1(n661_adj_4906), 
            .CO(n51038));
    SB_LUT4 add_6214_15_lut (.I0(GND_net), .I1(n16950[12]), .I2(n1041_adj_4908), 
            .I3(n50832), .O(n16339[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_9_lut (.I0(GND_net), .I1(n13134[6]), .I2(n588_adj_4909), 
            .I3(n51036), .O(n12072[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_15 (.CI(n50832), .I0(n16950[12]), .I1(n1041_adj_4908), 
            .CO(n50833));
    SB_LUT4 add_19_6_lut (.I0(GND_net), .I1(n258[4]), .I2(n303[4]), .I3(n50389), 
            .O(n353[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_9 (.CI(n51036), .I0(n13134[6]), .I1(n588_adj_4909), 
            .CO(n51037));
    SB_LUT4 add_6214_14_lut (.I0(GND_net), .I1(n16950[11]), .I2(n968_adj_4911), 
            .I3(n50831), .O(n16339[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_14 (.CI(n50831), .I0(n16950[11]), .I1(n968_adj_4911), 
            .CO(n50832));
    SB_LUT4 add_6214_13_lut (.I0(GND_net), .I1(n16950[10]), .I2(n895_adj_4912), 
            .I3(n50830), .O(n16339[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_8_lut (.I0(GND_net), .I1(n13134[5]), .I2(n515_adj_4913), 
            .I3(n51035), .O(n12072[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_8 (.CI(n51035), .I0(n13134[5]), .I1(n515_adj_4913), 
            .CO(n51036));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n54[6]), 
            .I3(n50507), .O(n433[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_10_lut (.I0(GND_net), .I1(n18613[7]), .I2(n685_adj_4915), 
            .I3(n51818), .O(n18225[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_10 (.CI(n51818), .I0(n18613[7]), .I1(n685_adj_4915), 
            .CO(n51819));
    SB_LUT4 add_6323_9_lut (.I0(GND_net), .I1(n18613[6]), .I2(n612_adj_4916), 
            .I3(n51817), .O(n18225[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_8 (.CI(n50507), .I0(GND_net), .I1(n54[6]), 
            .CO(n50508));
    SB_CARRY add_6323_9 (.CI(n51817), .I0(n18613[6]), .I1(n612_adj_4916), 
            .CO(n51818));
    SB_LUT4 add_6323_8_lut (.I0(GND_net), .I1(n18613[5]), .I2(n539_adj_4917), 
            .I3(n51816), .O(n18225[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_7_lut (.I0(GND_net), .I1(n13134[4]), .I2(n442_adj_4918), 
            .I3(n51034), .O(n12072[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_7 (.CI(n51034), .I0(n13134[4]), .I1(n442_adj_4918), 
            .CO(n51035));
    SB_CARRY add_6214_13 (.CI(n50830), .I0(n16950[10]), .I1(n895_adj_4912), 
            .CO(n50831));
    SB_CARRY add_6323_8 (.CI(n51816), .I0(n18613[5]), .I1(n539_adj_4917), 
            .CO(n51817));
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n54[5]), 
            .I3(n50506), .O(n433[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_7 (.CI(n50506), .I0(GND_net), .I1(n54[5]), 
            .CO(n50507));
    SB_CARRY add_19_6 (.CI(n50389), .I0(n258[4]), .I1(n303[4]), .CO(n50390));
    SB_LUT4 add_5992_6_lut (.I0(GND_net), .I1(n13134[3]), .I2(n369_adj_4920), 
            .I3(n51033), .O(n12072[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n54[4]), 
            .I3(n50505), .O(n433[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_7_lut (.I0(GND_net), .I1(n18613[4]), .I2(n466_adj_4922), 
            .I3(n51815), .O(n18225[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_15 (.CI(n52000), .I0(n12695[12]), .I1(n1023_adj_4899), 
            .CO(n52001));
    SB_LUT4 mult_18_add_1225_14_lut (.I0(GND_net), .I1(n12695[11]), .I2(n950_adj_4923), 
            .I3(n51999), .O(n303[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_6 (.CI(n51033), .I0(n13134[3]), .I1(n369_adj_4920), 
            .CO(n51034));
    SB_CARRY mult_18_add_1225_14 (.CI(n51999), .I0(n12695[11]), .I1(n950_adj_4923), 
            .CO(n52000));
    SB_CARRY add_6323_7 (.CI(n51815), .I0(n18613[4]), .I1(n466_adj_4922), 
            .CO(n51816));
    SB_CARRY unary_minus_27_add_3_6 (.CI(n50505), .I0(GND_net), .I1(n54[4]), 
            .CO(n50506));
    SB_LUT4 mult_18_add_1225_13_lut (.I0(GND_net), .I1(n12695[10]), .I2(n877_adj_4924), 
            .I3(n51998), .O(n303[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_13 (.CI(n51998), .I0(n12695[10]), .I1(n877_adj_4924), 
            .CO(n51999));
    SB_LUT4 mult_18_add_1225_12_lut (.I0(GND_net), .I1(n12695[9]), .I2(n804_adj_4925), 
            .I3(n51997), .O(n303[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_12 (.CI(n51997), .I0(n12695[9]), .I1(n804_adj_4925), 
            .CO(n51998));
    SB_LUT4 add_6323_6_lut (.I0(GND_net), .I1(n18613[3]), .I2(n393_adj_4926), 
            .I3(n51814), .O(n18225[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_add_1225_11_lut (.I0(GND_net), .I1(n12695[8]), .I2(n731_adj_4927), 
            .I3(n51996), .O(n303[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n48[3]), 
            .I2(n48[2]), .I3(GND_net), .O(n6_adj_4928));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n54[3]), 
            .I3(n50504), .O(n433[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6214_12_lut (.I0(GND_net), .I1(n16950[9]), .I2(n822_adj_4930), 
            .I3(n50829), .O(n16339[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_5_lut (.I0(GND_net), .I1(n13134[2]), .I2(n296_adj_4931), 
            .I3(n51032), .O(n12072[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n50504), .I0(GND_net), .I1(n54[3]), 
            .CO(n50505));
    SB_CARRY mult_18_add_1225_11 (.CI(n51996), .I0(n12695[8]), .I1(n731_adj_4927), 
            .CO(n51997));
    SB_CARRY add_6323_6 (.CI(n51814), .I0(n18613[3]), .I1(n393_adj_4926), 
            .CO(n51815));
    SB_CARRY add_6214_12 (.CI(n50829), .I0(n16950[9]), .I1(n822_adj_4930), 
            .CO(n50830));
    SB_LUT4 mult_18_add_1225_10_lut (.I0(GND_net), .I1(n12695[7]), .I2(n658_adj_4932), 
            .I3(n51995), .O(n303[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_10 (.CI(n51995), .I0(n12695[7]), .I1(n658_adj_4932), 
            .CO(n51996));
    SB_LUT4 mult_18_i296_2_lut (.I0(\Ki[6] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4933));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n54[2]), 
            .I3(n50503), .O(n433[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_18_add_1225_9_lut (.I0(GND_net), .I1(n12695[6]), .I2(n585_adj_4935), 
            .I3(n51994), .O(n303[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_5_lut (.I0(GND_net), .I1(n18613[2]), .I2(n320_adj_4936), 
            .I3(n51813), .O(n18225[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_9 (.CI(n51994), .I0(n12695[6]), .I1(n585_adj_4935), 
            .CO(n51995));
    SB_LUT4 mult_18_add_1225_8_lut (.I0(GND_net), .I1(n12695[5]), .I2(n512_adj_4937), 
            .I3(n51993), .O(n303[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_8 (.CI(n51993), .I0(n12695[5]), .I1(n512_adj_4937), 
            .CO(n51994));
    SB_CARRY add_6323_5 (.CI(n51813), .I0(n18613[2]), .I1(n320_adj_4936), 
            .CO(n51814));
    SB_LUT4 mult_18_add_1225_7_lut (.I0(GND_net), .I1(n12695[4]), .I2(n439_adj_4933), 
            .I3(n51992), .O(n303[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_5 (.CI(n51032), .I0(n13134[2]), .I1(n296_adj_4931), 
            .CO(n51033));
    SB_CARRY mult_18_add_1225_7 (.CI(n51992), .I0(n12695[4]), .I1(n439_adj_4933), 
            .CO(n51993));
    SB_CARRY unary_minus_27_add_3_4 (.CI(n50503), .I0(GND_net), .I1(n54[2]), 
            .CO(n50504));
    SB_LUT4 mult_18_add_1225_6_lut (.I0(GND_net), .I1(n12695[3]), .I2(n366_adj_4898), 
            .I3(n51991), .O(n303[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_6 (.CI(n51991), .I0(n12695[3]), .I1(n366_adj_4898), 
            .CO(n51992));
    SB_LUT4 mult_18_add_1225_5_lut (.I0(GND_net), .I1(n12695[2]), .I2(n293_adj_4890), 
            .I3(n51990), .O(n303[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_5 (.CI(n51990), .I0(n12695[2]), .I1(n293_adj_4890), 
            .CO(n51991));
    SB_LUT4 mult_18_i345_2_lut (.I0(\Ki[7] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4937));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_add_1225_4_lut (.I0(GND_net), .I1(n12695[1]), .I2(n220_adj_4887), 
            .I3(n51989), .O(n303[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_4 (.CI(n51989), .I0(n12695[1]), .I1(n220_adj_4887), 
            .CO(n51990));
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n54[1]), 
            .I3(n50502), .O(n433[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_4_lut (.I0(GND_net), .I1(n13134[1]), .I2(n223_adj_4885), 
            .I3(n51031), .O(n12072[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n50502), .I0(GND_net), .I1(n54[1]), 
            .CO(n50503));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n54[0]), 
            .I3(VCC_net), .O(n433[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n54[0]), 
            .CO(n50502));
    SB_LUT4 mult_18_add_1225_3_lut (.I0(GND_net), .I1(n12695[0]), .I2(n147_adj_4876), 
            .I3(n51988), .O(n303[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_3 (.CI(n51988), .I0(n12695[0]), .I1(n147_adj_4876), 
            .CO(n51989));
    SB_CARRY add_5992_4 (.CI(n51031), .I0(n13134[1]), .I1(n223_adj_4885), 
            .CO(n51032));
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(n353[23]), .I1(GND_net), .I2(n46[23]), 
            .I3(n50501), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_18_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4861), .I2(n74_adj_4859), 
            .I3(GND_net), .O(n303[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_18_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_18_add_1225_2 (.CI(GND_net), .I0(n5_adj_4861), .I1(n74_adj_4859), 
            .CO(n51988));
    SB_LUT4 add_6041_23_lut (.I0(GND_net), .I1(n13661[20]), .I2(GND_net), 
            .I3(n51987), .O(n12695[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_4_lut (.I0(GND_net), .I1(n18613[1]), .I2(n247_adj_4858), 
            .I3(n51812), .O(n18225[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_3_lut (.I0(GND_net), .I1(n13134[0]), .I2(n150_adj_4857), 
            .I3(n51030), .O(n12072[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n46[22]), 
            .I3(n50500), .O(n379[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_4 (.CI(n51812), .I0(n18613[1]), .I1(n247_adj_4858), 
            .CO(n51813));
    SB_LUT4 add_6323_3_lut (.I0(GND_net), .I1(n18613[0]), .I2(n174_adj_4853), 
            .I3(n51811), .O(n18225[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_3 (.CI(n51811), .I0(n18613[0]), .I1(n174_adj_4853), 
            .CO(n51812));
    SB_LUT4 add_6323_2_lut (.I0(GND_net), .I1(n32_adj_4850), .I2(n101_adj_4849), 
            .I3(GND_net), .O(n18225[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6214_11_lut (.I0(GND_net), .I1(n16950[8]), .I2(n749_adj_4839), 
            .I3(n50828), .O(n16339[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6214_11 (.CI(n50828), .I0(n16950[8]), .I1(n749_adj_4839), 
            .CO(n50829));
    SB_CARRY add_5992_3 (.CI(n51030), .I0(n13134[0]), .I1(n150_adj_4857), 
            .CO(n51031));
    SB_LUT4 add_6214_10_lut (.I0(GND_net), .I1(n16950[7]), .I2(n676_adj_4838), 
            .I3(n50827), .O(n16339[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_19_5_lut (.I0(GND_net), .I1(n258[3]), .I2(n303[3]), .I3(n50388), 
            .O(n353[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_19_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_2 (.CI(GND_net), .I0(n32_adj_4850), .I1(n101_adj_4849), 
            .CO(n51811));
    SB_CARRY add_6214_10 (.CI(n50827), .I0(n16950[7]), .I1(n676_adj_4838), 
            .CO(n50828));
    SB_LUT4 unary_minus_21_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[9]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i216_2_lut (.I0(\Ki[4] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4936));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i394_2_lut (.I0(\Ki[8] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4935));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[2]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i443_2_lut (.I0(\Ki[9] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4932));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Kp[4] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4931));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Kp[11] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4930));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6214_9_lut (.I0(GND_net), .I1(n16950[6]), .I2(n603), .I3(n50826), 
            .O(n16339[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6214_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6349_14_lut (.I0(GND_net), .I1(n18947[11]), .I2(n980_adj_4834), 
            .I3(n51810), .O(n18613[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6349_13_lut (.I0(GND_net), .I1(n18947[10]), .I2(n907_adj_4829), 
            .I3(n51809), .O(n18613[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6349_13 (.CI(n51809), .I0(n18947[10]), .I1(n907_adj_4829), 
            .CO(n51810));
    SB_LUT4 add_5992_2_lut (.I0(GND_net), .I1(n8_adj_4787), .I2(n77_adj_4783), 
            .I3(GND_net), .O(n12072[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[3]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i492_2_lut (.I0(\Ki[10] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4927));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i265_2_lut (.I0(\Ki[5] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4926));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6349_12_lut (.I0(GND_net), .I1(n18947[9]), .I2(n834), 
            .I3(n51808), .O(n18613[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6349_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_2 (.CI(GND_net), .I0(n8_adj_4787), .I1(n77_adj_4783), 
            .CO(n51030));
    SB_LUT4 mult_18_i541_2_lut (.I0(\Ki[11] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4925));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i590_2_lut (.I0(\Ki[12] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4924));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i639_2_lut (.I0(\Ki[13] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4923));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i314_2_lut (.I0(\Ki[6] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4922));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[4]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i161_2_lut (.I0(\Ki[3] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4747));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Kp[5] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4920));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[5]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Kp[6] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4918));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i363_2_lut (.I0(\Ki[7] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4917));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Kp[2] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i412_2_lut (.I0(\Ki[8] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4916));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[10]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[11]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i461_2_lut (.I0(\Ki[9] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4915));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[6]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Kp[7] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4913));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Kp[12] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4912));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Kp[13] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4911));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i210_2_lut (.I0(\Ki[4] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4746));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Kp[8] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4909));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Kp[14] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4908));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Kp[15] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4907));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Kp[9] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4906));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Kp[10] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4905));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[7]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Kp[11] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4903));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Kp[12] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4902));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[8]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i688_2_lut (.I0(\Ki[14] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4899));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[9]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Kp[13] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4896));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[10]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[12]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Kp[14] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4894));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i510_2_lut (.I0(\Ki[10] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4893));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Kp[15] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4892));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[11]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i737_2_lut (.I0(\Ki[15] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4888));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i559_2_lut (.I0(\Ki[11] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4884));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i75_2_lut (.I0(\Kp[1] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4883));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Kp[0] ), .I1(n105[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4882));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Kp[2] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4881));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i608_2_lut (.I0(\Ki[12] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4880));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Kp[3] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4879));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Kp[4] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4877));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[13]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[14]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Kp[5] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4875));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Kp[3] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i30_2_lut (.I0(\Ki[0] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4873));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Kp[6] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4872));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Kp[7] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4871));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Kp[8] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4870));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Kp[9] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4869));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51692_3_lut_4_lut (.I0(deadband[3]), .I1(n353[3]), .I2(n353[2]), 
            .I3(deadband[2]), .O(n67418));   // verilog/motorControl.v(56[16:33])
    defparam i51692_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Kp[10] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4868));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Kp[11] ), .I1(n105[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4867));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[12]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i657_2_lut (.I0(\Ki[13] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4862));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n353[3]), 
            .I2(n353[2]), .I3(GND_net), .O(n6_adj_4611));   // verilog/motorControl.v(56[16:33])
    defparam LessThan_20_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_18_i706_2_lut (.I0(\Ki[14] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4860));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Kp[1] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4855));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Kp[0] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4854));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Kp[2] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4852));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51694_2_lut_4_lut (.I0(n48[21]), .I1(n49[21]), .I2(n48[9]), 
            .I3(n49[9]), .O(n67420));
    defparam i51694_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Kp[3] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4851));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Kp[4] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4848));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Kp[5] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4846));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Kp[6] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4845));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51717_2_lut_4_lut (.I0(n48[16]), .I1(n49[16]), .I2(n48[7]), 
            .I3(n49[7]), .O(n67443));
    defparam i51717_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Kp[7] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4844));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Kp[8] ), .I1(n105[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4843));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[13]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50893_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n48[21]), .I2(IntegralLimit[9]), 
            .I3(n48[9]), .O(n66619));
    defparam i50893_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_15_i3_3_lut (.I0(n48[2]), .I1(n49[2]), .I2(n182), .I3(GND_net), 
            .O(n208[2]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i3_3_lut (.I0(n208[2]), .I1(IntegralLimit[2]), .I2(n156), 
            .I3(GND_net), .O(n233[2]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i53_2_lut (.I0(\Ki[1] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i6_2_lut (.I0(\Ki[0] ), .I1(n233[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4446));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[15]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i67_2_lut (.I0(\Ki[1] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4833));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i20_2_lut (.I0(\Ki[0] ), .I1(n233[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4832));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i116_2_lut (.I0(\Ki[2] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4831));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[16]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50927_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n48[16]), .I2(IntegralLimit[7]), 
            .I3(n48[7]), .O(n66653));
    defparam i50927_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Kp[4] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i102_2_lut (.I0(\Ki[2] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4444));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i165_2_lut (.I0(\Ki[3] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4830));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i214_2_lut (.I0(\Ki[4] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4828));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i263_2_lut (.I0(\Ki[5] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4827));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i312_2_lut (.I0(\Ki[6] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4826));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i361_2_lut (.I0(\Ki[7] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4825));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i469_2_lut (.I0(\Ki[9] ), .I1(n244), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4824));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[14]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i518_2_lut (.I0(\Ki[10] ), .I1(n244), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4822));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[15]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[16]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i259_2_lut (.I0(\Ki[5] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4745));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[17]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i81_2_lut (.I0(\Ki[1] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4817));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i34_2_lut (.I0(\Ki[0] ), .I1(n233[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i130_2_lut (.I0(\Ki[2] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4816));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i410_2_lut (.I0(\Ki[8] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4815));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i179_2_lut (.I0(\Ki[3] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[18]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i228_2_lut (.I0(\Ki[4] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i277_2_lut (.I0(\Ki[5] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i459_2_lut (.I0(\Ki[9] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4813));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[19]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i326_2_lut (.I0(\Ki[6] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4810));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i375_2_lut (.I0(\Ki[7] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i424_2_lut (.I0(\Ki[8] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Kp[1] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4809));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Kp[0] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4808));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Kp[2] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4807));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Kp[3] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4806));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i508_2_lut (.I0(\Ki[10] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4805));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Kp[4] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4804));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[20]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[21]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_18_i557_2_lut (.I0(\Ki[11] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4800));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Kp[5] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4799));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Kp[6] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4798));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i606_2_lut (.I0(\Ki[12] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4797));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Kp[7] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4796));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[22]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n54[23]));   // verilog/motorControl.v(60[26:35])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Kp[8] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4793));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Kp[9] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4792));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[17]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Kp[10] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4791));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Kp[11] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4790));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Kp[12] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4789));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Kp[13] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4788));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Kp[14] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4786));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i655_2_lut (.I0(\Ki[13] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4785));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Kp[15] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4784));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Kp[7] ), .I1(n105[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[21]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(IntegralLimit[18]), .I1(n48[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4939));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(IntegralLimit[19]), .I1(n48[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4940));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(IntegralLimit[20]), .I1(n135), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4941));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(IntegralLimit[17]), .I1(n48[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4942));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(IntegralLimit[16]), .I1(n48[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4943));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(IntegralLimit[14]), .I1(n48[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4944));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(IntegralLimit[13]), .I1(n48[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4945));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(IntegralLimit[15]), .I1(n48[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4946));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(IntegralLimit[11]), .I1(n48[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4947));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(IntegralLimit[12]), .I1(n48[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4948));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(IntegralLimit[21]), .I1(n48[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4949));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_18_i151_2_lut (.I0(\Ki[3] ), .I1(n233[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Kp[5] ), .I1(n105[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(IntegralLimit[22]), .I1(n48[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4950));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_21_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[18]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51022_4_lut (.I0(n21_adj_4621), .I1(n19_adj_4622), .I2(n17_adj_4623), 
            .I3(n9_adj_4618), .O(n66748));
    defparam i51022_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_15_i1_3_lut (.I0(n48[0]), .I1(n49[0]), .I2(n182), .I3(GND_net), 
            .O(n208[0]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i1_3_lut (.I0(n208[0]), .I1(IntegralLimit[0]), .I2(n156), 
            .I3(GND_net), .O(n233[0]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50990_4_lut (.I0(n27_adj_4945), .I1(n15_adj_4620), .I2(n13_adj_4619), 
            .I3(n36515), .O(n66716));
    defparam i50990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n48[7]), .I1(n48[16]), .I2(n33_adj_4943), 
            .I3(GND_net), .O(n12_adj_4952));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i2_2_lut (.I0(\Ki[0] ), .I1(n233[0]), .I2(GND_net), 
            .I3(GND_net), .O(n303[0]));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Kp[0] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n258[0]));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[19]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n150), .I1(n48[6]), .I2(n13_adj_4619), 
            .I3(GND_net), .O(n10_adj_4953));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4952), .I1(n48[17]), .I2(n35_adj_4942), 
            .I3(GND_net), .O(n30_adj_4954));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i704_2_lut (.I0(\Ki[14] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4782));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Kp[1] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Kp[0] ), .I1(n105[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4781));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51944_4_lut (.I0(n13_adj_4619), .I1(n36515), .I2(n9_adj_4618), 
            .I3(n66769), .O(n67670));
    defparam i51944_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51934_4_lut (.I0(n19_adj_4622), .I1(n17_adj_4623), .I2(n15_adj_4620), 
            .I3(n67670), .O(n67660));
    defparam i51934_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_18_i753_2_lut (.I0(\Ki[15] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4780));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53179_4_lut (.I0(n25_adj_4948), .I1(n23_adj_4947), .I2(n21_adj_4621), 
            .I3(n67660), .O(n68905));
    defparam i53179_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52567_4_lut (.I0(n31_adj_4946), .I1(n29_adj_4944), .I2(n27_adj_4945), 
            .I3(n68905), .O(n68293));
    defparam i52567_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Kp[2] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4779));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i65_2_lut (.I0(\Ki[1] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4778));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53354_4_lut (.I0(n37_adj_4939), .I1(n35_adj_4942), .I2(n33_adj_4943), 
            .I3(n68293), .O(n69080));
    defparam i53354_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_18_i18_2_lut (.I0(\Ki[0] ), .I1(n233[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4777));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n48[9]), .I1(n48[21]), .I2(n43_adj_4949), 
            .I3(GND_net), .O(n16_adj_4955));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52621_3_lut (.I0(n6_adj_4928), .I1(n48[10]), .I2(n21_adj_4621), 
            .I3(GND_net), .O(n68347));   // verilog/motorControl.v(50[16:38])
    defparam i52621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Kp[3] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4776));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52622_3_lut (.I0(n68347), .I1(n48[11]), .I2(n23_adj_4947), 
            .I3(GND_net), .O(n68348));   // verilog/motorControl.v(50[16:38])
    defparam i52622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n48[4]), .I1(n48[8]), .I2(n17_adj_4623), 
            .I3(GND_net), .O(n8_adj_4956));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_4955), .I1(n48[22]), .I2(n45_adj_4950), 
            .I3(GND_net), .O(n24_adj_4957));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50899_4_lut (.I0(n43_adj_4949), .I1(n25_adj_4948), .I2(n23_adj_4947), 
            .I3(n66748), .O(n66625));
    defparam i50899_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Kp[4] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4775));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52559_4_lut (.I0(n24_adj_4957), .I1(n8_adj_4956), .I2(n45_adj_4950), 
            .I3(n66619), .O(n68285));   // verilog/motorControl.v(50[16:38])
    defparam i52559_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_18_i114_2_lut (.I0(\Ki[2] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4774));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Kp[5] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4773));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51865_3_lut (.I0(n68348), .I1(n48[12]), .I2(n25_adj_4948), 
            .I3(GND_net), .O(n67591));   // verilog/motorControl.v(50[16:38])
    defparam i51865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(n48[0]), .I1(n48[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4958));   // verilog/motorControl.v(50[16:38])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i53159_3_lut (.I0(n4_adj_4958), .I1(n48[13]), .I2(n27_adj_4945), 
            .I3(GND_net), .O(n68885));   // verilog/motorControl.v(50[16:38])
    defparam i53159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53160_3_lut (.I0(n68885), .I1(n48[14]), .I2(n29_adj_4944), 
            .I3(GND_net), .O(n68886));   // verilog/motorControl.v(50[16:38])
    defparam i53160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i163_2_lut (.I0(\Ki[3] ), .I1(n233[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4772));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Kp[6] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4771));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50938_4_lut (.I0(n33_adj_4943), .I1(n31_adj_4946), .I2(n29_adj_4944), 
            .I3(n66716), .O(n66664));
    defparam i50938_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Kp[7] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Kp[8] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53393_4_lut (.I0(n30_adj_4954), .I1(n10_adj_4953), .I2(n35_adj_4942), 
            .I3(n66653), .O(n69119));   // verilog/motorControl.v(50[16:38])
    defparam i53393_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i71_2_lut (.I0(\Kp[1] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4744));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i24_2_lut (.I0(\Kp[0] ), .I1(n105[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4743));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52869_3_lut (.I0(n68886), .I1(n48[15]), .I2(n31_adj_4946), 
            .I3(GND_net), .O(n68595));   // verilog/motorControl.v(50[16:38])
    defparam i52869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Kp[2] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4742));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53522_4_lut (.I0(n68595), .I1(n69119), .I2(n35_adj_4942), 
            .I3(n66664), .O(n69248));   // verilog/motorControl.v(50[16:38])
    defparam i53522_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53523_3_lut (.I0(n69248), .I1(n48[18]), .I2(n37_adj_4939), 
            .I3(GND_net), .O(n69249));   // verilog/motorControl.v(50[16:38])
    defparam i53523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i308_2_lut (.I0(\Ki[6] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4741));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53491_3_lut (.I0(n69249), .I1(n48[19]), .I2(n39_adj_4940), 
            .I3(GND_net), .O(n69217));   // verilog/motorControl.v(50[16:38])
    defparam i53491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50902_4_lut (.I0(n43_adj_4949), .I1(n41_adj_4941), .I2(n39_adj_4940), 
            .I3(n69080), .O(n66628));
    defparam i50902_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53165_4_lut (.I0(n67591), .I1(n68285), .I2(n45_adj_4950), 
            .I3(n66625), .O(n68891));   // verilog/motorControl.v(50[16:38])
    defparam i53165_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Kp[1] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4769));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53438_3_lut (.I0(n69217), .I1(n135), .I2(n41_adj_4941), .I3(GND_net), 
            .O(n40_adj_4959));   // verilog/motorControl.v(50[16:38])
    defparam i53438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53167_4_lut (.I0(n40_adj_4959), .I1(n68891), .I2(n45_adj_4950), 
            .I3(n66628), .O(n68893));   // verilog/motorControl.v(50[16:38])
    defparam i53167_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_18_i357_2_lut (.I0(\Ki[7] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4740));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53168_3_lut (.I0(n68893), .I1(IntegralLimit[23]), .I2(n48[23]), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(50[16:38])
    defparam i53168_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Kp[0] ), .I1(n105[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4768));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_13_i37_2_lut (.I0(n48[18]), .I1(n49[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4960));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Kp[9] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_13_i39_2_lut (.I0(n48[19]), .I1(n49[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4961));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i35_2_lut (.I0(n48[17]), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4962));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i33_2_lut (.I0(n48[16]), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4963));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i29_2_lut (.I0(n48[14]), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4964));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i31_2_lut (.I0(n48[15]), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4965));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Kp[10] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Kp[2] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4767));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Kp[3] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4739));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Kp[4] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4738));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_13_i27_2_lut (.I0(n48[13]), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4966));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i45_2_lut (.I0(n48[22]), .I1(n49[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4967));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i23_2_lut (.I0(n48[11]), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4968));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i25_2_lut (.I0(n48[12]), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4969));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_13_i43_2_lut (.I0(n48[21]), .I1(n49[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4970));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50872_4_lut (.I0(n21_adj_4629), .I1(n19_adj_4630), .I2(n17_adj_4632), 
            .I3(n9_adj_4624), .O(n66598));
    defparam i50872_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50813_4_lut (.I0(n27_adj_4966), .I1(n15_adj_4627), .I2(n13_adj_4626), 
            .I3(n11_adj_4625), .O(n66539));
    defparam i50813_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Kp[11] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Kp[3] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4766));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_13_i12_3_lut (.I0(n49[7]), .I1(n49[16]), .I2(n33_adj_4963), 
            .I3(GND_net), .O(n12_adj_4971));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_13_i10_3_lut (.I0(n49[5]), .I1(n49[6]), .I2(n13_adj_4626), 
            .I3(GND_net), .O(n10_adj_4972));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Kp[4] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4765));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_13_i30_3_lut (.I0(n12_adj_4971), .I1(n49[17]), .I2(n35_adj_4962), 
            .I3(GND_net), .O(n30_adj_4973));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51774_4_lut (.I0(n13_adj_4626), .I1(n11_adj_4625), .I2(n9_adj_4624), 
            .I3(n66612), .O(n67500));
    defparam i51774_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51768_4_lut (.I0(n19_adj_4630), .I1(n17_adj_4632), .I2(n15_adj_4627), 
            .I3(n67500), .O(n67494));
    defparam i51768_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53123_4_lut (.I0(n25_adj_4969), .I1(n23_adj_4968), .I2(n21_adj_4629), 
            .I3(n67494), .O(n68849));
    defparam i53123_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Kp[12] ), .I1(n105[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Kp[5] ), .I1(n105[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4764));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36342_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n50278));   // verilog/motorControl.v(55[22:28])
    defparam i36342_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i36153_2_lut_3_lut (.I0(\Kp[0] ), .I1(n105[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n50063));   // verilog/motorControl.v(55[22:28])
    defparam i36153_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i52489_4_lut (.I0(n31_adj_4965), .I1(n29_adj_4964), .I2(n27_adj_4966), 
            .I3(n68849), .O(n68215));
    defparam i52489_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53348_4_lut (.I0(n37_adj_4960), .I1(n35_adj_4962), .I2(n33_adj_4963), 
            .I3(n68215), .O(n69074));
    defparam i53348_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_13_i16_3_lut (.I0(n49[9]), .I1(n49[21]), .I2(n43_adj_4970), 
            .I3(GND_net), .O(n16_adj_4974));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53109_3_lut (.I0(n6_adj_4863), .I1(n49[10]), .I2(n21_adj_4629), 
            .I3(GND_net), .O(n68835));   // verilog/motorControl.v(52[25:48])
    defparam i53109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53110_3_lut (.I0(n68835), .I1(n49[11]), .I2(n23_adj_4968), 
            .I3(GND_net), .O(n68836));   // verilog/motorControl.v(52[25:48])
    defparam i53110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_13_i8_3_lut (.I0(n49[4]), .I1(n49[8]), .I2(n17_adj_4632), 
            .I3(GND_net), .O(n8_adj_4975));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_13_i24_3_lut (.I0(n16_adj_4974), .I1(n49[22]), .I2(n45_adj_4967), 
            .I3(GND_net), .O(n24_adj_4976));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51696_4_lut (.I0(n43_adj_4970), .I1(n25_adj_4969), .I2(n23_adj_4968), 
            .I3(n66598), .O(n67422));
    defparam i51696_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52561_4_lut (.I0(n24_adj_4976), .I1(n8_adj_4975), .I2(n45_adj_4967), 
            .I3(n67420), .O(n68287));   // verilog/motorControl.v(52[25:48])
    defparam i52561_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52873_3_lut (.I0(n68836), .I1(n49[12]), .I2(n25_adj_4969), 
            .I3(GND_net), .O(n68599));   // verilog/motorControl.v(52[25:48])
    defparam i52873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_13_i4_4_lut (.I0(n48[0]), .I1(n49[1]), .I2(n48[1]), 
            .I3(n49[0]), .O(n4_adj_4977));   // verilog/motorControl.v(52[25:48])
    defparam LessThan_13_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53107_3_lut (.I0(n4_adj_4977), .I1(n49[13]), .I2(n27_adj_4966), 
            .I3(GND_net), .O(n68833));   // verilog/motorControl.v(52[25:48])
    defparam i53107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53108_3_lut (.I0(n68833), .I1(n49[14]), .I2(n29_adj_4964), 
            .I3(GND_net), .O(n68834));   // verilog/motorControl.v(52[25:48])
    defparam i53108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50779_4_lut (.I0(n33_adj_4963), .I1(n31_adj_4965), .I2(n29_adj_4964), 
            .I3(n66539), .O(n66505));
    defparam i50779_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53306_4_lut (.I0(n30_adj_4973), .I1(n10_adj_4972), .I2(n35_adj_4962), 
            .I3(n67443), .O(n69032));   // verilog/motorControl.v(52[25:48])
    defparam i53306_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52875_3_lut (.I0(n68834), .I1(n49[15]), .I2(n31_adj_4965), 
            .I3(GND_net), .O(n28));   // verilog/motorControl.v(52[25:48])
    defparam i52875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53451_4_lut (.I0(n28), .I1(n69032), .I2(n35_adj_4962), .I3(n66505), 
            .O(n69177));   // verilog/motorControl.v(52[25:48])
    defparam i53451_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53452_3_lut (.I0(n69177), .I1(n49[18]), .I2(n37_adj_4960), 
            .I3(GND_net), .O(n69178));   // verilog/motorControl.v(52[25:48])
    defparam i53452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53379_3_lut (.I0(n69178), .I1(n49[19]), .I2(n39_adj_4961), 
            .I3(GND_net), .O(n69105));   // verilog/motorControl.v(52[25:48])
    defparam i53379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51699_4_lut (.I0(n43_adj_4970), .I1(n41_adj_3), .I2(n39_adj_4961), 
            .I3(n69074), .O(n67425));
    defparam i51699_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53169_4_lut (.I0(n68599), .I1(n68287), .I2(n45_adj_4967), 
            .I3(n67422), .O(n68895));   // verilog/motorControl.v(52[25:48])
    defparam i53169_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51871_3_lut (.I0(n69105), .I1(n187), .I2(n41_adj_3), .I3(GND_net), 
            .O(n67597));   // verilog/motorControl.v(52[25:48])
    defparam i51871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53360_4_lut (.I0(n67597), .I1(n68895), .I2(n45_adj_4967), 
            .I3(n67425), .O(n69086));   // verilog/motorControl.v(52[25:48])
    defparam i53360_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53361_3_lut (.I0(n69086), .I1(n48[23]), .I2(n49[23]), .I3(GND_net), 
            .O(n182));   // verilog/motorControl.v(52[25:48])
    defparam i53361_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_15_i11_3_lut (.I0(n48[10]), .I1(n49[10]), .I2(n182), .I3(GND_net), 
            .O(n208[10]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_962 (.I0(\data_in_frame[9][7] ), .I1(\data_in_frame[6][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4979));   // verilog/coms.v(99[12:25])
    defparam i2_2_lut_adj_962.LUT_INIT = 16'h6666;
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[8][4] ), .I1(\data_in_frame[8][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4980));   // verilog/coms.v(99[12:25])
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut (.I0(n58520), .I1(\data_in_frame[4][2] ), .I2(\data_in_frame[8][6] ), 
            .I3(\data_in_frame[1][6] ), .O(n24_adj_4981));   // verilog/coms.v(99[12:25])
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(\data_in_frame[12][0] ), .I1(n16_adj_4979), .I2(n58075), 
            .I3(n58405), .O(n22_adj_4982));   // verilog/coms.v(99[12:25])
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut (.I0(n58556), .I1(n24_adj_4981), .I2(n18_adj_4980), 
            .I3(\data_in_frame[3][7] ), .O(n26_adj_4983));   // verilog/coms.v(99[12:25])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[4][1] ), .I1(n26_adj_4983), .I2(n22_adj_4982), 
            .I3(\data_in_frame[8][3] ), .O(n58766));   // verilog/coms.v(99[12:25])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_16_i11_3_lut (.I0(n208[10]), .I1(IntegralLimit[10]), .I2(n156), 
            .I3(GND_net), .O(n233[10]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i561_2_lut (.I0(\Ki[11] ), .I1(n233[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n46[22]));   // verilog/motorControl.v(56[47:56])
    defparam unary_minus_21_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51503_2_lut_4_lut (.I0(n353[9]), .I1(n433[9]), .I2(n353[5]), 
            .I3(n433[5]), .O(n67229));
    defparam i51503_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51508_2_lut_4_lut (.I0(n353[7]), .I1(n433[7]), .I2(n353[6]), 
            .I3(n433[6]), .O(n67234));
    defparam i51508_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51545_2_lut_4_lut (.I0(PWMLimit[8]), .I1(n353[8]), .I2(PWMLimit[4]), 
            .I3(n353[4]), .O(n67271));
    defparam i51545_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51549_2_lut_4_lut (.I0(PWMLimit[6]), .I1(n353[6]), .I2(PWMLimit[5]), 
            .I3(n353[5]), .O(n67275));
    defparam i51549_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_18_i406_2_lut (.I0(\Ki[8] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4718));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i455_2_lut (.I0(\Ki[9] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i504_2_lut (.I0(\Ki[10] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i553_2_lut (.I0(\Ki[11] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i602_2_lut (.I0(\Ki[12] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i651_2_lut (.I0(\Ki[13] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i700_2_lut (.I0(\Ki[14] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Kp[5] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4712));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Kp[6] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4711));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51606_2_lut_4_lut (.I0(deadband[21]), .I1(n353[21]), .I2(deadband[9]), 
            .I3(n353[9]), .O(n67332));
    defparam i51606_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Kp[7] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4710));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i749_2_lut (.I0(\Ki[15] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51616_2_lut_4_lut (.I0(deadband[16]), .I1(n353[16]), .I2(deadband[7]), 
            .I3(n353[7]), .O(n67342));
    defparam i51616_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i36280_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n233[21]), .I2(\Ki[1] ), 
            .I3(n37050), .O(n20183[0]));   // verilog/motorControl.v(55[31:42])
    defparam i36280_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36282_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n233[21]), .I2(\Ki[1] ), 
            .I3(n37050), .O(n50204));   // verilog/motorControl.v(55[31:42])
    defparam i36282_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i36096_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n233[19]), .I2(\Ki[1] ), 
            .I3(n37154), .O(n20109[0]));   // verilog/motorControl.v(55[31:42])
    defparam i36096_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36098_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n233[19]), .I2(\Ki[1] ), 
            .I3(n37154), .O(n50001));   // verilog/motorControl.v(55[31:42])
    defparam i36098_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i36316_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n20183[0]), 
            .O(n4_adj_4434));   // verilog/motorControl.v(55[31:42])
    defparam i36316_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_963 (.I0(n62), .I1(n131), .I2(n204), .I3(n20183[0]), 
            .O(n20158));   // verilog/motorControl.v(55[31:42])
    defparam i1_3_lut_4_lut_adj_963.LUT_INIT = 16'h8778;
    SB_LUT4 i36303_2_lut_4_lut (.I0(n37050), .I1(\Ki[0] ), .I2(\Ki[1] ), 
            .I3(n233[19]), .O(n20159));   // verilog/motorControl.v(55[31:42])
    defparam i36303_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Kp[8] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4680));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i61_2_lut (.I0(\Ki[1] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i14_2_lut (.I0(\Ki[0] ), .I1(n233[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4679));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i110_2_lut (.I0(\Ki[2] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Kp[9] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4672));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i159_2_lut (.I0(\Ki[3] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4670));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i208_2_lut (.I0(\Ki[4] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i257_2_lut (.I0(\Ki[5] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4668));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i306_2_lut (.I0(\Ki[6] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4667));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i355_2_lut (.I0(\Ki[7] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i404_2_lut (.I0(\Ki[8] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i453_2_lut (.I0(\Ki[9] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i502_2_lut (.I0(\Ki[10] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i551_2_lut (.I0(\Ki[11] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Kp[10] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4655));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i600_2_lut (.I0(\Ki[12] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Kp[11] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4653));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i16_3_lut (.I0(n48[15]), .I1(n49[15]), .I2(n182), .I3(GND_net), 
            .O(n208[15]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i16_3_lut (.I0(n208[15]), .I1(IntegralLimit[15]), .I2(n156), 
            .I3(GND_net), .O(n233[15]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_18_i79_2_lut (.I0(\Ki[1] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4652));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i32_2_lut (.I0(\Ki[0] ), .I1(n233[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4651));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i128_2_lut (.I0(\Ki[2] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4648));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Kp[12] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Kp[13] ), .I1(n105[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(55[22:28])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i177_2_lut (.I0(\Ki[3] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i649_2_lut (.I0(\Ki[13] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_18_i698_2_lut (.I0(\Ki[14] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28955_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n42880));   // verilog/motorControl.v(42[14] 67[8])
    defparam i28955_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15636_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[4]), 
            .I3(\PID_CONTROLLER.integral [4]), .O(n29667));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15636_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15634_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[5]), 
            .I3(\PID_CONTROLLER.integral [5]), .O(n29665));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15634_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15632_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[6]), 
            .I3(\PID_CONTROLLER.integral [6]), .O(n29663));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15632_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mult_18_i226_2_lut (.I0(\Ki[4] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16375_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[23]), 
            .I3(\PID_CONTROLLER.integral [23]), .O(n30406));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16376_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[22]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n30407));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16379_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[21]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n30410));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16379_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n37050), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n30411));   // verilog/motorControl.v(45[18] 66[12])
    defparam i8_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16413_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[19]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n30444));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16413_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23184_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n37154), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n30446));   // verilog/motorControl.v(45[18] 66[12])
    defparam i23184_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16416_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[17]), 
            .I3(\PID_CONTROLLER.integral [17]), .O(n30447));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16418_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[16]), 
            .I3(\PID_CONTROLLER.integral [16]), .O(n30449));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16418_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mult_18_i747_2_lut (.I0(\Ki[15] ), .I1(n233[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16419_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[15]), 
            .I3(\PID_CONTROLLER.integral [15]), .O(n30450));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16419_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16425_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[14]), 
            .I3(\PID_CONTROLLER.integral [14]), .O(n30456));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mult_18_i275_2_lut (.I0(\Ki[5] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n244), 
            .I3(\PID_CONTROLLER.integral [13]), .O(n30457));   // verilog/motorControl.v(45[18] 66[12])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16427_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[12]), 
            .I3(\PID_CONTROLLER.integral [12]), .O(n30458));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16428_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[11]), 
            .I3(\PID_CONTROLLER.integral [11]), .O(n30459));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15588_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[0]), 
            .I3(\PID_CONTROLLER.integral [0]), .O(n29619));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15588_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mult_18_i324_2_lut (.I0(\Ki[6] ), .I1(n233[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4637));   // verilog/motorControl.v(55[31:42])
    defparam mult_18_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15601_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[10]), 
            .I3(\PID_CONTROLLER.integral [10]), .O(n29632));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15601_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15629_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[9]), 
            .I3(\PID_CONTROLLER.integral [9]), .O(n29660));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15629_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15630_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[8]), 
            .I3(\PID_CONTROLLER.integral [8]), .O(n29661));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15630_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15631_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[7]), 
            .I3(\PID_CONTROLLER.integral [7]), .O(n29662));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15631_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15637_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[3]), 
            .I3(\PID_CONTROLLER.integral [3]), .O(n29668));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15637_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15665_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[2]), 
            .I3(\PID_CONTROLLER.integral [2]), .O(n29696));   // verilog/motorControl.v(45[18] 66[12])
    defparam i15665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16196_3_lut_4_lut (.I0(control_update), .I1(n15), .I2(n233[1]), 
            .I3(\PID_CONTROLLER.integral [1]), .O(n30227));   // verilog/motorControl.v(45[18] 66[12])
    defparam i16196_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_15_i10_3_lut (.I0(n48[9]), .I1(n49[9]), .I2(n182), .I3(GND_net), 
            .O(n208[9]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i10_3_lut (.I0(n208[9]), .I1(IntegralLimit[9]), .I2(n156), 
            .I3(GND_net), .O(n233[9]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i9_3_lut (.I0(n48[8]), .I1(n49[8]), .I2(n182), .I3(GND_net), 
            .O(n208[8]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i9_3_lut (.I0(n208[8]), .I1(IntegralLimit[8]), .I2(n156), 
            .I3(GND_net), .O(n233[8]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n48[7]), .I1(n49[7]), .I2(n182), .I3(GND_net), 
            .O(n208[7]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_16_i8_3_lut (.I0(n208[7]), .I1(IntegralLimit[7]), .I2(n156), 
            .I3(GND_net), .O(n233[7]));   // verilog/motorControl.v(52[22] 54[16])
    defparam mux_16_i8_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
