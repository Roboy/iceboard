// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Jan 28 22:25:46 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    output SCL;   // verilog/TinyFPGA_B.v(21[10:13])
    input SDA /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, CLK_c, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(42[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(88[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(89[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(123[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(125[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(126[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(127[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(128[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(130[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(131[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(132[22:35])
    
    wire n4;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(162[22:33])
    wire [22:0]pwm_setpoint_22__N_3;
    
    wire RX_N_2;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]motor_state_23__N_50;
    wire [23:0]displacement_23__N_26;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    wire [31:0]one_wire_N_399;
    
    wire n2252, n20822, n4141, n14886, n14885, n18789, n14884, 
        n14883, n14882, n14881, n14880, n14879, n14878, n14877, 
        n30126, n14876, n14875, n14874, n14873;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n3, n4_adj_4462, n5, n6, n7, n8, n9, n10, n11, n12, 
        n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
        n23, n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active, n14872;
    wire [31:0]\FRAME_MATCHER.state_31__N_2380 ;
    
    wire n14869, n14868, n14867, n1554, n14866, n14865, n14864, 
        n14863, n14862, n14861, n14860, n14859, n14858, n14857, 
        n14856, n14855, n14854, n14853, n14852, n14851, n14850, 
        n14849, n14848, n30820, n15_adj_4463, n10_adj_4464, n29356, 
        n29966, n29350, n29347, n29343, n29341, n13551, n22113, 
        n22112, n22111, n25063, n22110, n22109, n22108, n22107, 
        n22106, n22105, n22104, n22050, n22049, n22103, n12_adj_4465, 
        n22102, n22048, n14847, n14846, n22101, n13497, n26880, 
        n22047, n22046, n26858, n26856, n22100, n22045, n22099, 
        n22044, n22043, n22042, n22041, n26836, n22098, n22097, 
        n22096, n22040, n22039, n22095, n22094, n22038, n22093, 
        n22092, n22037, n26748, n30875, n22036, n22035, n22034, 
        n22033, n22091, n15348, n15347, n15346, n15342, n15337, 
        n15336, n15335, n15334, n15333, n15332, n15331, n15330, 
        n15329, n15328, n15327, n15326, n15325, n15324, n15323, 
        n15322, n15321, n15320, n15319, n15318, n15317, n15316, 
        n15315, n15314, n15313, n15312, n15311, n15310, n15309, 
        n15308, n1, n14845, n14844, n22032, n22031, n22030, n22029, 
        n15132, n15131, n15130, n15129, n15128, n15127, n15126, 
        n15125, n15124, n15123, n15122, n15121, n15120, n15119, 
        n15118, n15117, n15116, n15115, n15114, n15113, n15112, 
        n15111, n15110, n15109, n15108, n15107, n15106, n15105, 
        n15104, n7_adj_4466, n4_adj_4467, n15103, n15102, n63, n15101, 
        n15100, n15099, n15098, n15097, n15096, n15095, quadA_debounced, 
        quadB_debounced, n15094, n15093, quadA_debounced_adj_4468, quadB_debounced_adj_4469, 
        n15092, n15091, n15090, n15089, n15088, n15087, n15086, 
        n14766, n15085, n15084, n15083, n15082, n15081, n15080, 
        n14672, n15079, n15077, n15076, n15075, n15074, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n15073, n15072, n15071, n15070, n15069, n5_adj_4470, n4_adj_4471, 
        n4137, n15068, n15067, n15066, n15065, n15064, n15063, 
        n15062, n15061, n15060, n15059, n15058, n15057, n15056, 
        n3_adj_4472, n15055, n4_adj_4473, n15054, n15053;
    wire [2:0]r_SM_Main_2__N_3262;
    
    wire n15052, n15051, n15050, n14843, n15049, n15048, n15047, 
        n15046, n15045, n15044, n15043, n15042, n15041, n15040, 
        n15039, n15038;
    wire [2:0]r_SM_Main_adj_4567;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_4569;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3333;
    
    wire n15037, n15036, n15035, n15034, n15033, n15032, n15031, 
        n15030, n15029, n15028, n15027, n15026, n15025, n15024, 
        n15023, n15022, n15021, n15020, n15019, n15018, n15017, 
        n15016, n15015, n15014, n15013;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15012, n15011, n15_adj_4478, n15010, n15009;
    wire [1:0]reg_B_adj_4578;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15008, n15007, n15006, n15005, n2, n14641, n15004, n15003, 
        n15002, n15001, n15000, n14999, n14998, n14997, n14996, 
        n14995, n14994, n14993, n14992, n14991, n14990, n14621, 
        n14989, n14988, n14987, n14986, n14985, n14984, n14983, 
        n14982, n14981, n14980, n14979, n14978, n14977, n14976, 
        n14975, n14974, n14973, n14972, n14971, n4_adj_4481, n14970, 
        n30123, n14969, n14968, n14967, n14966, n14965, n14964, 
        n14963, n14962, n14961, n14960, n14959, n14958, n14957, 
        n14956, n14955, n14954, n14953, n14952, n14951, n6_adj_4482, 
        n7_adj_4483, n8_adj_4484, n9_adj_4485, n10_adj_4486, n11_adj_4487, 
        n12_adj_4488, n13_adj_4489, n14_adj_4490, n15_adj_4491, n16_adj_4492, 
        n17_adj_4493, n18_adj_4494, n19_adj_4495, n20_adj_4496, n21_adj_4497, 
        n22_adj_4498, n23_adj_4499, n24_adj_4500, n25_adj_4501, n14950, 
        n14842, n14841, n14840, n30127, n30055, n29873, n4_adj_4502, 
        n6_adj_4503, n7_adj_4504, n8_adj_4505, n9_adj_4506, n10_adj_4507, 
        n11_adj_4508, n12_adj_4509, n13_adj_4510, n15_adj_4511, n17_adj_4512, 
        n19_adj_4513, n21_adj_4514, n29972, n23_adj_4515, n25_adj_4516, 
        n27, n29970, n29, n30, n31, n33, n35, n30074, n30054, 
        n29973, n29971, n29954, n29948, n5_adj_4517, n7_adj_4518, 
        n29946, n14949, n14948, n14947, n14946, n14945, n14944, 
        n14943, n14942, n14941, n14940, n14939, n14938, n14937, 
        n14936, n14935, n14934, n14933, n14932, n14931, n14930, 
        n14929, n14928, n14927, n14926, n14925, n14924, n14923, 
        n14922, n14921, n14920, n14919, n14918, n14839, n14836, 
        n14835, n14834, n14833, n14832, n14917, n14916, n14915, 
        n14914, n14913, n14912, n14911, n14910, n14830, n14829, 
        n14828, n14827, n14826, n14825, n14824, n14823, n14909, 
        n14908, n14907, n14906, n14905, n14904, n14903, n14902, 
        n14901, n14900, n14899, n14898, n14897, n14896, n14895, 
        n14894, n14893, n14892, n14891, n14890, n14889, n14888, 
        n14887, n29637, n29627, n28285, n27156, n7375, n13407, 
        n4_adj_4519, n26029, n29903, n14822, n14821, n29819, n29821, 
        n25777, n14820, n14818, n14817, n30261, n4_adj_4520, n28241, 
        n28236, n24343, n13405, n13399, n29235, n13556, n29233, 
        n3_adj_4521, n10896, n30128, n26399, n29210, n28;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .data_o({quadA_debounced, quadB_debounced}), 
            .GND_net(GND_net), .n28241(n28241), .reg_B({reg_B}), .VCC_net(VCC_net), 
            .n14834(n14834), .ENCODER0_B_c_0(ENCODER0_B_c_0), .n15347(n15347), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(185[15] 190[4])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_26 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF h2_25 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 i11284_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n10896), .I3(GND_net), .O(n15089));   // verilog/coms.v(127[12] 300[6])
    defparam i11284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[14]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4483));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    neopixel nx (.GND_net(GND_net), .clk32MHz(clk32MHz), .n26858(n26858), 
            .n28(n28), .\state[0] (state[0]), .\state[1] (state[1]), .\one_wire_N_399[11] (one_wire_N_399[11]), 
            .n1554(n1554), .timer({timer}), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .VCC_net(VCC_net), .n20822(n20822), .n29233(n29233), .n14869(n14869), 
            .n14868(n14868), .n4(n4_adj_4519), .neopxl_color({neopxl_color}), 
            .n14867(n14867), .n14866(n14866), .n29210(n29210), .n14865(n14865), 
            .n14864(n14864), .n14863(n14863), .n14862(n14862), .n14861(n14861), 
            .n14860(n14860), .n14859(n14859), .n14858(n14858), .n14857(n14857), 
            .n14856(n14856), .n14855(n14855), .n14854(n14854), .n14853(n14853), 
            .n14852(n14852), .n14851(n14851), .n14850(n14850), .n14849(n14849), 
            .n14848(n14848), .n14847(n14847), .n14846(n14846), .n14845(n14845), 
            .n14844(n14844), .n14843(n14843), .n14842(n14842), .n14841(n14841), 
            .n14840(n14840), .n14839(n14839), .n12(n12_adj_4465), .n25063(n25063), 
            .LED_c(LED_c), .n14817(n14817), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(44[10] 50[2])
    SB_LUT4 i11064_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n1554), .I3(GND_net), .O(n14869));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[15]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11285_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n10896), .I3(GND_net), .O(n15090));   // verilog/coms.v(127[12] 300[6])
    defparam i11285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11286_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n10896), .I3(GND_net), .O(n15091));   // verilog/coms.v(127[12] 300[6])
    defparam i11286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11287_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n10896), .I3(GND_net), .O(n15092));   // verilog/coms.v(127[12] 300[6])
    defparam i11287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11288_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n10896), .I3(GND_net), .O(n15093));   // verilog/coms.v(127[12] 300[6])
    defparam i11288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[16]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11289_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n10896), .I3(GND_net), .O(n15094));   // verilog/coms.v(127[12] 300[6])
    defparam i11289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11290_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n10896), .I3(GND_net), .O(n15095));   // verilog/coms.v(127[12] 300[6])
    defparam i11290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11291_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n10896), .I3(GND_net), .O(n15096));   // verilog/coms.v(127[12] 300[6])
    defparam i11291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11292_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n10896), .I3(GND_net), .O(n15097));   // verilog/coms.v(127[12] 300[6])
    defparam i11292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11293_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n10896), .I3(GND_net), .O(n15098));   // verilog/coms.v(127[12] 300[6])
    defparam i11293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[17]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11294_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n10896), .I3(GND_net), .O(n15099));   // verilog/coms.v(127[12] 300[6])
    defparam i11294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11295_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n10896), .I3(GND_net), .O(n15100));   // verilog/coms.v(127[12] 300[6])
    defparam i11295_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dir_30 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 i11296_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n10896), .I3(GND_net), .O(n15101));   // verilog/coms.v(127[12] 300[6])
    defparam i11296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11297_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n10896), .I3(GND_net), .O(n15102));   // verilog/coms.v(127[12] 300[6])
    defparam i11297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11298_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n10896), .I3(GND_net), .O(n15103));   // verilog/coms.v(127[12] 300[6])
    defparam i11298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[18]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11299_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n10896), .I3(GND_net), .O(n15104));   // verilog/coms.v(127[12] 300[6])
    defparam i11299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4482));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11300_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n10896), .I3(GND_net), .O(n15105));   // verilog/coms.v(127[12] 300[6])
    defparam i11300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[19]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11301_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n10896), .I3(GND_net), .O(n15106));   // verilog/coms.v(127[12] 300[6])
    defparam i11301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11302_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n10896), .I3(GND_net), .O(n15107));   // verilog/coms.v(127[12] 300[6])
    defparam i11302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11303_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n10896), .I3(GND_net), .O(n15108));   // verilog/coms.v(127[12] 300[6])
    defparam i11303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11305_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n4141), .I3(GND_net), .O(n15110));   // verilog/coms.v(127[12] 300[6])
    defparam i11305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11306_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n4141), .I3(GND_net), .O(n15111));   // verilog/coms.v(127[12] 300[6])
    defparam i11306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11307_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n4141), .I3(GND_net), .O(n15112));   // verilog/coms.v(127[12] 300[6])
    defparam i11307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11308_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n4141), .I3(GND_net), .O(n15113));   // verilog/coms.v(127[12] 300[6])
    defparam i11308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11309_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n4141), .I3(GND_net), .O(n15114));   // verilog/coms.v(127[12] 300[6])
    defparam i11309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11310_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n4141), .I3(GND_net), .O(n15115));   // verilog/coms.v(127[12] 300[6])
    defparam i11310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11311_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n4141), .I3(GND_net), .O(n15116));   // verilog/coms.v(127[12] 300[6])
    defparam i11311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11312_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n4141), .I3(GND_net), .O(n15117));   // verilog/coms.v(127[12] 300[6])
    defparam i11312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11313_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n4141), .I3(GND_net), .O(n15118));   // verilog/coms.v(127[12] 300[6])
    defparam i11313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11314_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n4141), .I3(GND_net), .O(n15119));   // verilog/coms.v(127[12] 300[6])
    defparam i11314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11315_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n4141), .I3(GND_net), .O(n15120));   // verilog/coms.v(127[12] 300[6])
    defparam i11315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11061_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n1554), .I3(GND_net), .O(n14866));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11316_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n4141), .I3(GND_net), .O(n15121));   // verilog/coms.v(127[12] 300[6])
    defparam i11316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11317_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n4141), .I3(GND_net), .O(n15122));   // verilog/coms.v(127[12] 300[6])
    defparam i11317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[20]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[21]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11318_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n4141), .I3(GND_net), .O(n15123));   // verilog/coms.v(127[12] 300[6])
    defparam i11318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11319_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n4141), .I3(GND_net), .O(n15124));   // verilog/coms.v(127[12] 300[6])
    defparam i11319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11320_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n4141), .I3(GND_net), .O(n15125));   // verilog/coms.v(127[12] 300[6])
    defparam i11320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11321_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n4141), .I3(GND_net), .O(n15126));   // verilog/coms.v(127[12] 300[6])
    defparam i11321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11322_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n4141), .I3(GND_net), .O(n15127));   // verilog/coms.v(127[12] 300[6])
    defparam i11322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[22]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11323_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n4141), .I3(GND_net), .O(n15128));   // verilog/coms.v(127[12] 300[6])
    defparam i11323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4470));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11324_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n4141), .I3(GND_net), .O(n15129));   // verilog/coms.v(127[12] 300[6])
    defparam i11324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11325_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n4141), .I3(GND_net), .O(n15130));   // verilog/coms.v(127[12] 300[6])
    defparam i11325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11326_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n4141), .I3(GND_net), .O(n15131));   // verilog/coms.v(127[12] 300[6])
    defparam i11326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(control_mode[3]), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(control_mode[7]), .O(n10_adj_4464));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11327_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n4141), .I3(GND_net), .O(n15132));   // verilog/coms.v(127[12] 300[6])
    defparam i11327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4464), .I2(control_mode[2]), 
            .I3(GND_net), .O(n13497));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(n13399), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4478));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n13497), 
            .I3(GND_net), .O(n15_adj_4463));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_38_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[23]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11062_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n1554), .I3(GND_net), .O(n14867));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4489));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4471));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4472));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4488));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[7]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[8]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4487));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4462));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[9]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11067_3_lut (.I0(n26880), .I1(r_Bit_Index_adj_4569[0]), .I2(n26856), 
            .I3(GND_net), .O(n14872));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11067_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i11068_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n4137), .I3(GND_net), .O(n14873));   // verilog/coms.v(127[12] 300[6])
    defparam i11068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4486));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4485));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11063_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n1554), .I3(GND_net), .O(n14868));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[10]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4484));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[11]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11069_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n4137), .I3(GND_net), .O(n14874));   // verilog/coms.v(127[12] 300[6])
    defparam i11069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(143[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[12]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[13]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11070_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n4137), .I3(GND_net), .O(n14875));   // verilog/coms.v(127[12] 300[6])
    defparam i11070_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF h1_24 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCL_pad (.PACKAGE_PIN(SCL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCL_pad.PIN_TYPE = 6'b011001;
    defparam SCL_pad.PULLUP = 1'b0;
    defparam SCL_pad.NEG_TRIGGER = 1'b0;
    defparam SCL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_483_24_lut (.I0(duty[22]), .I1(n30261), .I2(n3), .I3(n22050), 
            .O(pwm_setpoint_22__N_3[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_483_23_lut (.I0(duty[21]), .I1(n30261), .I2(n4_adj_4462), 
            .I3(n22049), .O(pwm_setpoint_22__N_3[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_23_lut.LUT_INIT = 16'h8BB8;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[0]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_CARRY add_483_23 (.CI(n22049), .I0(n30261), .I1(n4_adj_4462), .CO(n22050));
    SB_LUT4 add_483_22_lut (.I0(duty[20]), .I1(n30261), .I2(n5), .I3(n22048), 
            .O(pwm_setpoint_22__N_3[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_22 (.CI(n22048), .I0(n30261), .I1(n5), .CO(n22049));
    SB_LUT4 add_483_21_lut (.I0(duty[19]), .I1(n30261), .I2(n6), .I3(n22047), 
            .O(pwm_setpoint_22__N_3[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_21 (.CI(n22047), .I0(n30261), .I1(n6), .CO(n22048));
    SB_LUT4 add_483_20_lut (.I0(duty[18]), .I1(n30261), .I2(n7), .I3(n22046), 
            .O(pwm_setpoint_22__N_3[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_20 (.CI(n22046), .I0(n30261), .I1(n7), .CO(n22047));
    SB_LUT4 add_483_19_lut (.I0(duty[17]), .I1(n30261), .I2(n8), .I3(n22045), 
            .O(pwm_setpoint_22__N_3[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_19 (.CI(n22045), .I0(n30261), .I1(n8), .CO(n22046));
    SB_LUT4 i11078_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n4137), .I3(GND_net), .O(n14883));   // verilog/coms.v(127[12] 300[6])
    defparam i11078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11071_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n4137), .I3(GND_net), .O(n14876));   // verilog/coms.v(127[12] 300[6])
    defparam i11071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11072_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n4137), .I3(GND_net), .O(n14877));   // verilog/coms.v(127[12] 300[6])
    defparam i11072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11073_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n4137), .I3(GND_net), .O(n14878));   // verilog/coms.v(127[12] 300[6])
    defparam i11073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_483_18_lut (.I0(duty[16]), .I1(n30261), .I2(n9), .I3(n22044), 
            .O(pwm_setpoint_22__N_3[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_18 (.CI(n22044), .I0(n30261), .I1(n9), .CO(n22045));
    SB_LUT4 i11079_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n4137), .I3(GND_net), .O(n14884));   // verilog/coms.v(127[12] 300[6])
    defparam i11079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_483_17_lut (.I0(duty[15]), .I1(n30261), .I2(n10), .I3(n22043), 
            .O(pwm_setpoint_22__N_3[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_17 (.CI(n22043), .I0(n30261), .I1(n10), .CO(n22044));
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n2), .I3(n22113), .O(displacement_23__N_26[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_483_16_lut (.I0(duty[14]), .I1(n30261), .I2(n11), .I3(n22042), 
            .O(pwm_setpoint_22__N_3[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4472), .I3(n22112), .O(displacement_23__N_26[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11074_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n4137), .I3(GND_net), .O(n14879));   // verilog/coms.v(127[12] 300[6])
    defparam i11074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11075_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n4137), .I3(GND_net), .O(n14880));   // verilog/coms.v(127[12] 300[6])
    defparam i11075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11076_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n4137), .I3(GND_net), .O(n14881));   // verilog/coms.v(127[12] 300[6])
    defparam i11076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11077_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n4137), .I3(GND_net), .O(n14882));   // verilog/coms.v(127[12] 300[6])
    defparam i11077_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n22112), .I0(encoder1_position[22]), 
            .I1(n3_adj_4472), .CO(n22113));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_26[23]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n4_adj_4471), .I3(n22111), .O(displacement_23__N_26[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11503_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4137), .I3(GND_net), .O(n15308));   // verilog/coms.v(127[12] 300[6])
    defparam i11503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11504_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4137), .I3(GND_net), .O(n15309));   // verilog/coms.v(127[12] 300[6])
    defparam i11504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11505_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4137), .I3(GND_net), .O(n15310));   // verilog/coms.v(127[12] 300[6])
    defparam i11505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11506_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4137), .I3(GND_net), .O(n15311));   // verilog/coms.v(127[12] 300[6])
    defparam i11506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11507_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4137), .I3(GND_net), .O(n15312));   // verilog/coms.v(127[12] 300[6])
    defparam i11507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11508_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4137), .I3(GND_net), .O(n15313));   // verilog/coms.v(127[12] 300[6])
    defparam i11508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11509_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4137), .I3(GND_net), .O(n15314));   // verilog/coms.v(127[12] 300[6])
    defparam i11509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11510_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n4137), .I3(GND_net), .O(n15315));   // verilog/coms.v(127[12] 300[6])
    defparam i11510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11511_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n4137), .I3(GND_net), .O(n15316));   // verilog/coms.v(127[12] 300[6])
    defparam i11511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11512_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n4137), .I3(GND_net), .O(n15317));   // verilog/coms.v(127[12] 300[6])
    defparam i11512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11513_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n4137), .I3(GND_net), .O(n15318));   // verilog/coms.v(127[12] 300[6])
    defparam i11513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11514_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n4137), .I3(GND_net), .O(n15319));   // verilog/coms.v(127[12] 300[6])
    defparam i11514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11515_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n4137), .I3(GND_net), .O(n15320));   // verilog/coms.v(127[12] 300[6])
    defparam i11515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11516_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n4137), .I3(GND_net), .O(n15321));   // verilog/coms.v(127[12] 300[6])
    defparam i11516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11517_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n4137), .I3(GND_net), .O(n15322));   // verilog/coms.v(127[12] 300[6])
    defparam i11517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11518_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n4137), .I3(GND_net), .O(n15323));   // verilog/coms.v(127[12] 300[6])
    defparam i11518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11519_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n4137), .I3(GND_net), .O(n15324));   // verilog/coms.v(127[12] 300[6])
    defparam i11519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11520_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n4137), .I3(GND_net), .O(n15325));   // verilog/coms.v(127[12] 300[6])
    defparam i11520_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_26[22]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_26[21]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_26[20]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_26[19]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_26[18]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_26[17]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_26[16]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_26[15]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_26[14]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_26[13]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_26[12]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_26[11]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_26[10]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_26[9]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_26[8]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_26[7]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_26[6]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_26[5]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_26[4]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_26[3]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_26[2]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_26[1]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[22]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[21]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[20]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[19]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[18]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[17]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[16]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[15]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[14]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[13]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[12]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[11]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[10]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[9]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[8]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[7]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[6]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[5]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[4]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[3]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[2]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[1]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 i11521_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n4137), .I3(GND_net), .O(n15326));   // verilog/coms.v(127[12] 300[6])
    defparam i11521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11522_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n4137), .I3(GND_net), .O(n15327));   // verilog/coms.v(127[12] 300[6])
    defparam i11522_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_483_16 (.CI(n22042), .I0(n30261), .I1(n11), .CO(n22043));
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n22111), .I0(encoder1_position[21]), 
            .I1(n4_adj_4471), .CO(n22112));
    SB_LUT4 i11523_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n4137), .I3(GND_net), .O(n15328));   // verilog/coms.v(127[12] 300[6])
    defparam i11523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11524_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n4137), .I3(GND_net), .O(n15329));   // verilog/coms.v(127[12] 300[6])
    defparam i11524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11525_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n4137), .I3(GND_net), .O(n15330));   // verilog/coms.v(127[12] 300[6])
    defparam i11525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11526_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n4137), .I3(GND_net), .O(n15331));   // verilog/coms.v(127[12] 300[6])
    defparam i11526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11527_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n4137), .I3(GND_net), .O(n15332));   // verilog/coms.v(127[12] 300[6])
    defparam i11527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4470), .I3(n22110), .O(displacement_23__N_26[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11528_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n4137), .I3(GND_net), .O(n15333));   // verilog/coms.v(127[12] 300[6])
    defparam i11528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11529_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n4137), .I3(GND_net), .O(n15334));   // verilog/coms.v(127[12] 300[6])
    defparam i11529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11530_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n4137), .I3(GND_net), .O(n15335));   // verilog/coms.v(127[12] 300[6])
    defparam i11530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11531_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n4137), .I3(GND_net), .O(n15336));   // verilog/coms.v(127[12] 300[6])
    defparam i11531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11532_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n4137), .I3(GND_net), .O(n15337));   // verilog/coms.v(127[12] 300[6])
    defparam i11532_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n22110), .I0(encoder1_position[20]), 
            .I1(n5_adj_4470), .CO(n22111));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4482), .I3(n22109), .O(displacement_23__N_26[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(n63), .I1(n7_adj_4466), .I2(n4_adj_4467), .I3(n1), 
            .O(n30820));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i21779_4_lut (.I0(\FRAME_MATCHER.state_31__N_2380 [2]), .I1(n26748), 
            .I2(n2252), .I3(n3_adj_4521), .O(n26836));
    defparam i21779_4_lut.LUT_INIT = 16'haaa8;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n22109), .I0(encoder1_position[19]), 
            .I1(n6_adj_4482), .CO(n22110));
    SB_LUT4 i25166_4_lut (.I0(n63), .I1(n7_adj_4518), .I2(n26836), .I3(n5_adj_4517), 
            .O(n28285));   // verilog/coms.v(127[12] 300[6])
    defparam i25166_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4483), .I3(n22108), .O(displacement_23__N_26[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n22108), .I0(encoder1_position[18]), 
            .I1(n7_adj_4483), .CO(n22109));
    SB_LUT4 add_483_15_lut (.I0(duty[13]), .I1(n30261), .I2(n12), .I3(n22041), 
            .O(pwm_setpoint_22__N_3[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_15 (.CI(n22041), .I0(n30261), .I1(n12), .CO(n22042));
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4484), .I3(n22107), .O(displacement_23__N_26[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11541_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4473), 
            .I3(n13551), .O(n15346));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11541_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11542_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n28241), 
            .I3(GND_net), .O(n15347));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11542_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11543_3_lut (.I0(quadA_debounced_adj_4468), .I1(reg_B_adj_4578[1]), 
            .I2(n28236), .I3(GND_net), .O(n15348));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11543_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11537_3_lut (.I0(n14766), .I1(r_Bit_Index[0]), .I2(n14672), 
            .I3(GND_net), .O(n15342));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11537_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i24360_4_lut (.I0(n28), .I1(one_wire_N_399[11]), .I2(n26858), 
            .I3(state[0]), .O(n29235));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24360_4_lut.LUT_INIT = 16'hfcee;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i18_4_lut (.I0(n29235), .I1(n29233), .I2(state[1]), .I3(n4_adj_4519), 
            .O(n25063));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4501));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_483_14_lut (.I0(duty[12]), .I1(n30261), .I2(n13), .I3(n22040), 
            .O(pwm_setpoint_22__N_3[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n22107), .I0(encoder1_position[17]), 
            .I1(n8_adj_4484), .CO(n22108));
    SB_CARRY add_483_14 (.CI(n22040), .I0(n30261), .I1(n13), .CO(n22041));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4485), .I3(n22106), .O(displacement_23__N_26[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n22106), .I0(encoder1_position[16]), 
            .I1(n9_adj_4485), .CO(n22107));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4486), .I3(n22105), .O(displacement_23__N_26[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_483_13_lut (.I0(duty[11]), .I1(n30261), .I2(n14), .I3(n22039), 
            .O(pwm_setpoint_22__N_3[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11027_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4137), .I3(GND_net), .O(n14832));   // verilog/coms.v(127[12] 300[6])
    defparam i11027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11028_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n4137), .I3(GND_net), .O(n14833));   // verilog/coms.v(127[12] 300[6])
    defparam i11028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11029_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n28241), 
            .I3(GND_net), .O(n14834));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11029_3_lut.LUT_INIT = 16'hacac;
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i11030_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_4567[1]), .I2(n7375), 
            .I3(n4_adj_4520), .O(n14835));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11030_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i11031_3_lut (.I0(quadB_debounced_adj_4469), .I1(reg_B_adj_4578[0]), 
            .I2(n28236), .I3(GND_net), .O(n14836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26_4_lut (.I0(n29210), .I1(state[1]), .I2(n20822), .I3(GND_net), 
            .O(n12_adj_4465));   // verilog/neopixel.v(35[12] 117[6])
    defparam i26_4_lut.LUT_INIT = 16'h7474;
    SB_LUT4 i11034_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n1554), .I3(GND_net), .O(n14839));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11035_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n1554), .I3(GND_net), .O(n14840));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11036_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n1554), .I3(GND_net), .O(n14841));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11037_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n1554), .I3(GND_net), .O(n14842));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11038_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n1554), .I3(GND_net), .O(n14843));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11039_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n1554), .I3(GND_net), .O(n14844));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11040_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n1554), .I3(GND_net), .O(n14845));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11041_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n1554), .I3(GND_net), .O(n14846));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11042_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n1554), .I3(GND_net), .O(n14847));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11043_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n1554), .I3(GND_net), .O(n14848));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11044_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n1554), .I3(GND_net), .O(n14849));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11045_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n1554), .I3(GND_net), .O(n14850));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11046_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n1554), .I3(GND_net), .O(n14851));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11047_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n1554), .I3(GND_net), .O(n14852));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11048_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n1554), .I3(GND_net), .O(n14853));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11049_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n1554), .I3(GND_net), .O(n14854));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11050_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n1554), .I3(GND_net), .O(n14855));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11051_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n1554), .I3(GND_net), .O(n14856));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11052_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n1554), .I3(GND_net), .O(n14857));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11053_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n1554), .I3(GND_net), .O(n14858));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11054_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n1554), .I3(GND_net), .O(n14859));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11055_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n1554), .I3(GND_net), .O(n14860));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11056_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n1554), .I3(GND_net), .O(n14861));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11057_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n1554), .I3(GND_net), .O(n14862));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4500));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4499));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4498));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4497));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_483_13 (.CI(n22039), .I0(n30261), .I1(n14), .CO(n22040));
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n22105), .I0(encoder1_position[15]), 
            .I1(n10_adj_4486), .CO(n22106));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4487), .I3(n22104), .O(displacement_23__N_26[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_483_12_lut (.I0(duty[10]), .I1(n30261), .I2(n15), .I3(n22038), 
            .O(pwm_setpoint_22__N_3[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11058_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n1554), .I3(GND_net), .O(n14863));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11080_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n4137), .I3(GND_net), .O(n14885));   // verilog/coms.v(127[12] 300[6])
    defparam i11080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11059_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n1554), .I3(GND_net), .O(n14864));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11059_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_483_12 (.CI(n22038), .I0(n30261), .I1(n15), .CO(n22039));
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n22104), .I0(encoder1_position[14]), 
            .I1(n11_adj_4487), .CO(n22105));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4488), .I3(n22103), .O(displacement_23__N_26[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n22103), .I0(encoder1_position[13]), 
            .I1(n12_adj_4488), .CO(n22104));
    SB_LUT4 add_483_11_lut (.I0(duty[9]), .I1(n30261), .I2(n16), .I3(n22037), 
            .O(pwm_setpoint_22__N_3[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_11 (.CI(n22037), .I0(n30261), .I1(n16), .CO(n22038));
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4489), .I3(n22102), .O(displacement_23__N_26[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_483_10_lut (.I0(duty[8]), .I1(n30261), .I2(n17), .I3(n22036), 
            .O(pwm_setpoint_22__N_3[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4496));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3262[2]), 
            .I3(r_SM_Main[0]), .O(n14621));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n14621), 
            .I3(rx_data_ready), .O(n25777));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4495));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[0]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[1]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i25176_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n26029));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i25176_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4494));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n22102), .I0(encoder1_position[12]), 
            .I1(n13_adj_4489), .CO(n22103));
    SB_LUT4 mux_38_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[2]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4493));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11060_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n1554), .I3(GND_net), .O(n14865));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4490), .I3(n22101), .O(displacement_23__N_26[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_483_10 (.CI(n22036), .I0(n30261), .I1(n17), .CO(n22037));
    SB_LUT4 add_483_9_lut (.I0(duty[7]), .I1(n30261), .I2(n18), .I3(n22035), 
            .O(pwm_setpoint_22__N_3[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_38_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[3]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4492));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4491));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[4]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_37_i1_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[0]), 
            .I3(encoder0_position[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i2_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[1]), 
            .I3(encoder0_position[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i3_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[2]), 
            .I3(encoder0_position[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n22101), .I0(encoder1_position[11]), 
            .I1(n14_adj_4490), .CO(n22102));
    SB_CARRY add_483_9 (.CI(n22035), .I0(n30261), .I1(n18), .CO(n22036));
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_4567[1]), .I1(r_SM_Main_adj_4567[0]), 
            .I2(r_SM_Main_adj_4567[2]), .I3(r_SM_Main_2__N_3333[1]), .O(n30875));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 add_483_8_lut (.I0(duty[6]), .I1(n30261), .I2(n19), .I3(n22034), 
            .O(pwm_setpoint_22__N_3[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_483_8 (.CI(n22034), .I0(n30261), .I1(n19), .CO(n22035));
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4491), .I3(n22100), .O(displacement_23__N_26[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_483_7_lut (.I0(duty[5]), .I1(n30261), .I2(n20), .I3(n22033), 
            .O(pwm_setpoint_22__N_3[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n22100), .I0(encoder1_position[10]), 
            .I1(n15_adj_4491), .CO(n22101));
    SB_LUT4 LessThan_555_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4506));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4508));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4512));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4492), .I3(n22099), .O(displacement_23__N_26[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_555_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4511));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4510));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4504));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_483_7 (.CI(n22033), .I0(n30261), .I1(n20), .CO(n22034));
    SB_LUT4 LessThan_555_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4503));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_555_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4507));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24278_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n29341));
    defparam i24278_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_555_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4509));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_555_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4505));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_555_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4514));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4515));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24293_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n29356));
    defparam i24293_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_555_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4513));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_483_6_lut (.I0(duty[4]), .I1(n30261), .I2(n21), .I3(n22032), 
            .O(pwm_setpoint_22__N_3[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n22099), .I0(encoder1_position[9]), 
            .I1(n16_adj_4492), .CO(n22100));
    SB_LUT4 LessThan_555_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4516));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11081_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n4137), .I3(GND_net), .O(n14886));   // verilog/coms.v(127[12] 300[6])
    defparam i11081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11082_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n4137), .I3(GND_net), .O(n14887));   // verilog/coms.v(127[12] 300[6])
    defparam i11082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11083_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n4137), .I3(GND_net), .O(n14888));   // verilog/coms.v(127[12] 300[6])
    defparam i11083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11084_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n4137), .I3(GND_net), .O(n14889));   // verilog/coms.v(127[12] 300[6])
    defparam i11084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11085_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n4137), .I3(GND_net), .O(n14890));   // verilog/coms.v(127[12] 300[6])
    defparam i11085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11086_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n4137), .I3(GND_net), .O(n14891));   // verilog/coms.v(127[12] 300[6])
    defparam i11086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11087_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n4137), .I3(GND_net), .O(n14892));   // verilog/coms.v(127[12] 300[6])
    defparam i11087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11088_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n4137), .I3(GND_net), .O(n14893));   // verilog/coms.v(127[12] 300[6])
    defparam i11088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11089_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n4137), .I3(GND_net), .O(n14894));   // verilog/coms.v(127[12] 300[6])
    defparam i11089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11090_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n4137), .I3(GND_net), .O(n14895));   // verilog/coms.v(127[12] 300[6])
    defparam i11090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11091_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14896));   // verilog/coms.v(127[12] 300[6])
    defparam i11091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11092_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14897));   // verilog/coms.v(127[12] 300[6])
    defparam i11092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11093_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14898));   // verilog/coms.v(127[12] 300[6])
    defparam i11093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11094_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14899));   // verilog/coms.v(127[12] 300[6])
    defparam i11094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11095_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14900));   // verilog/coms.v(127[12] 300[6])
    defparam i11095_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_483_6 (.CI(n22032), .I0(n30261), .I1(n21), .CO(n22033));
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4493), .I3(n22098), .O(displacement_23__N_26[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n22098), .I0(encoder1_position[8]), 
            .I1(n17_adj_4493), .CO(n22099));
    SB_LUT4 i11096_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14901));   // verilog/coms.v(127[12] 300[6])
    defparam i11096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11097_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14902));   // verilog/coms.v(127[12] 300[6])
    defparam i11097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_483_5_lut (.I0(duty[3]), .I1(n30261), .I2(n22), .I3(n22031), 
            .O(pwm_setpoint_22__N_3[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11098_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14903));   // verilog/coms.v(127[12] 300[6])
    defparam i11098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4494), .I3(n22097), .O(displacement_23__N_26[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11099_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14904));   // verilog/coms.v(127[12] 300[6])
    defparam i11099_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n22097), .I0(encoder1_position[7]), 
            .I1(n18_adj_4494), .CO(n22098));
    SB_CARRY add_483_5 (.CI(n22031), .I0(n30261), .I1(n22), .CO(n22032));
    SB_LUT4 i11100_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14905));   // verilog/coms.v(127[12] 300[6])
    defparam i11100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11101_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14906));   // verilog/coms.v(127[12] 300[6])
    defparam i11101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11102_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14907));   // verilog/coms.v(127[12] 300[6])
    defparam i11102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11103_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14908));   // verilog/coms.v(127[12] 300[6])
    defparam i11103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4495), .I3(n22096), .O(displacement_23__N_26[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_483_4_lut (.I0(duty[2]), .I1(n30261), .I2(n23), .I3(n22030), 
            .O(pwm_setpoint_22__N_3[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11104_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14909));   // verilog/coms.v(127[12] 300[6])
    defparam i11104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11105_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14910));   // verilog/coms.v(127[12] 300[6])
    defparam i11105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11106_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14911));   // verilog/coms.v(127[12] 300[6])
    defparam i11106_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n22096), .I0(encoder1_position[6]), 
            .I1(n19_adj_4495), .CO(n22097));
    SB_LUT4 i11107_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14912));   // verilog/coms.v(127[12] 300[6])
    defparam i11107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4496), .I3(n22095), .O(displacement_23__N_26[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11108_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14913));   // verilog/coms.v(127[12] 300[6])
    defparam i11108_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n22095), .I0(encoder1_position[5]), 
            .I1(n20_adj_4496), .CO(n22096));
    SB_CARRY add_483_4 (.CI(n22030), .I0(n30261), .I1(n23), .CO(n22031));
    SB_LUT4 i11109_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14914));   // verilog/coms.v(127[12] 300[6])
    defparam i11109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_483_3_lut (.I0(duty[1]), .I1(n30261), .I2(n24), .I3(n22029), 
            .O(pwm_setpoint_22__N_3[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11110_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14915));   // verilog/coms.v(127[12] 300[6])
    defparam i11110_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_483_3 (.CI(n22029), .I0(n30261), .I1(n24), .CO(n22030));
    SB_LUT4 i11111_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14916));   // verilog/coms.v(127[12] 300[6])
    defparam i11111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11112_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14917));   // verilog/coms.v(127[12] 300[6])
    defparam i11112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11113_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14918));   // verilog/coms.v(127[12] 300[6])
    defparam i11113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11114_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14919));   // verilog/coms.v(127[12] 300[6])
    defparam i11114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11115_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14920));   // verilog/coms.v(127[12] 300[6])
    defparam i11115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11116_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14921));   // verilog/coms.v(127[12] 300[6])
    defparam i11116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4497), .I3(n22094), .O(displacement_23__N_26[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11117_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14922));   // verilog/coms.v(127[12] 300[6])
    defparam i11117_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n22094), .I0(encoder1_position[4]), 
            .I1(n21_adj_4497), .CO(n22095));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4498), .I3(n22093), .O(displacement_23__N_26[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11118_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14923));   // verilog/coms.v(127[12] 300[6])
    defparam i11118_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n22093), .I0(encoder1_position[3]), 
            .I1(n22_adj_4498), .CO(n22094));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4499), .I3(n22092), .O(displacement_23__N_26[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n22092), .I0(encoder1_position[2]), 
            .I1(n23_adj_4499), .CO(n22093));
    SB_LUT4 i11119_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14924));   // verilog/coms.v(127[12] 300[6])
    defparam i11119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11120_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14925));   // verilog/coms.v(127[12] 300[6])
    defparam i11120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[5]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11121_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14926));   // verilog/coms.v(127[12] 300[6])
    defparam i11121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11122_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n27156), 
            .I3(GND_net), .O(n14927));   // verilog/coms.v(127[12] 300[6])
    defparam i11122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11123_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n27156), 
            .I3(GND_net), .O(n14928));   // verilog/coms.v(127[12] 300[6])
    defparam i11123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_483_2_lut (.I0(duty[0]), .I1(n30261), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_3[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_483_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4500), .I3(n22091), .O(displacement_23__N_26[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_483_2 (.CI(VCC_net), .I0(n30261), .I1(n25), .CO(n22029));
    SB_LUT4 mux_37_i4_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[3]), 
            .I3(encoder0_position[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11124_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n27156), 
            .I3(GND_net), .O(n14929));   // verilog/coms.v(127[12] 300[6])
    defparam i11124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11125_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n27156), 
            .I3(GND_net), .O(n14930));   // verilog/coms.v(127[12] 300[6])
    defparam i11125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11126_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n27156), 
            .I3(GND_net), .O(n14931));   // verilog/coms.v(127[12] 300[6])
    defparam i11126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4490));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11127_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n27156), 
            .I3(GND_net), .O(n14932));   // verilog/coms.v(127[12] 300[6])
    defparam i11127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11128_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n27156), 
            .I3(GND_net), .O(n14933));   // verilog/coms.v(127[12] 300[6])
    defparam i11128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11129_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n27156), 
            .I3(GND_net), .O(n14934));   // verilog/coms.v(127[12] 300[6])
    defparam i11129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11130_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n27156), 
            .I3(GND_net), .O(n14935));   // verilog/coms.v(127[12] 300[6])
    defparam i11130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11131_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n27156), 
            .I3(GND_net), .O(n14936));   // verilog/coms.v(127[12] 300[6])
    defparam i11131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11132_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n27156), 
            .I3(GND_net), .O(n14937));   // verilog/coms.v(127[12] 300[6])
    defparam i11132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11133_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n27156), 
            .I3(GND_net), .O(n14938));   // verilog/coms.v(127[12] 300[6])
    defparam i11133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11134_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n27156), 
            .I3(GND_net), .O(n14939));   // verilog/coms.v(127[12] 300[6])
    defparam i11134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11135_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n27156), 
            .I3(GND_net), .O(n14940));   // verilog/coms.v(127[12] 300[6])
    defparam i11135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_37_i5_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[4]), 
            .I3(encoder0_position[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11136_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n27156), 
            .I3(GND_net), .O(n14941));   // verilog/coms.v(127[12] 300[6])
    defparam i11136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11137_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n27156), 
            .I3(GND_net), .O(n14942));   // verilog/coms.v(127[12] 300[6])
    defparam i11137_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n22091), .I0(encoder1_position[1]), 
            .I1(n24_adj_4500), .CO(n22092));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4501), .I3(VCC_net), .O(displacement_23__N_26[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11138_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n27156), 
            .I3(GND_net), .O(n14943));   // verilog/coms.v(127[12] 300[6])
    defparam i11138_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11139_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n27156), 
            .I3(GND_net), .O(n14944));   // verilog/coms.v(127[12] 300[6])
    defparam i11139_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4501), .CO(n22091));
    SB_LUT4 i11140_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n27156), 
            .I3(GND_net), .O(n14945));   // verilog/coms.v(127[12] 300[6])
    defparam i11140_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11141_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n27156), 
            .I3(GND_net), .O(n14946));   // verilog/coms.v(127[12] 300[6])
    defparam i11141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11142_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n27156), 
            .I3(GND_net), .O(n14947));   // verilog/coms.v(127[12] 300[6])
    defparam i11142_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11143_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n27156), 
            .I3(GND_net), .O(n14948));   // verilog/coms.v(127[12] 300[6])
    defparam i11143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11144_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n27156), 
            .I3(GND_net), .O(n14949));   // verilog/coms.v(127[12] 300[6])
    defparam i11144_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_37_i6_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[5]), 
            .I3(encoder0_position[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_adj_1586 (.I0(n13405), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n13407));
    defparam i1_2_lut_adj_1586.LUT_INIT = 16'heeee;
    SB_LUT4 i24284_4_lut (.I0(n27), .I1(n15_adj_4511), .I2(n13_adj_4510), 
            .I3(n11_adj_4508), .O(n29347));
    defparam i24284_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24571_4_lut (.I0(n9_adj_4506), .I1(n7_adj_4504), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n29637));
    defparam i24571_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i24755_4_lut (.I0(n15_adj_4511), .I1(n13_adj_4510), .I2(n11_adj_4508), 
            .I3(n29637), .O(n29821));
    defparam i24755_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24753_4_lut (.I0(n21_adj_4514), .I1(n19_adj_4513), .I2(n17_adj_4512), 
            .I3(n29821), .O(n29819));
    defparam i24753_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24287_4_lut (.I0(n27), .I1(n25_adj_4516), .I2(n23_adj_4515), 
            .I3(n29819), .O(n29350));
    defparam i24287_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_555_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4502));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i24904_3_lut (.I0(n4_adj_4502), .I1(pwm_setpoint[13]), .I2(n27), 
            .I3(GND_net), .O(n29970));   // verilog/pwm.v(21[8:24])
    defparam i24904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_555_i30_3_lut (.I0(n12_adj_4509), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam LessThan_555_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24905_3_lut (.I0(n29970), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n29971));   // verilog/pwm.v(21[8:24])
    defparam i24905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24280_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n29347), 
            .O(n29343));
    defparam i24280_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25008_4_lut (.I0(n30), .I1(n10_adj_4507), .I2(n35), .I3(n29341), 
            .O(n30074));   // verilog/pwm.v(21[8:24])
    defparam i25008_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24882_3_lut (.I0(n29971), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n29948));   // verilog/pwm.v(21[8:24])
    defparam i24882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24906_3_lut (.I0(n6_adj_4503), .I1(pwm_setpoint[10]), .I2(n21_adj_4514), 
            .I3(GND_net), .O(n29972));   // verilog/pwm.v(21[8:24])
    defparam i24906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24907_3_lut (.I0(n29972), .I1(pwm_setpoint[11]), .I2(n23_adj_4515), 
            .I3(GND_net), .O(n29973));   // verilog/pwm.v(21[8:24])
    defparam i24907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24561_4_lut (.I0(n23_adj_4515), .I1(n21_adj_4514), .I2(n19_adj_4513), 
            .I3(n29356), .O(n29627));
    defparam i24561_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24807_3_lut (.I0(n8_adj_4505), .I1(pwm_setpoint[9]), .I2(n19_adj_4513), 
            .I3(GND_net), .O(n29873));   // verilog/pwm.v(21[8:24])
    defparam i24807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24880_3_lut (.I0(n29973), .I1(pwm_setpoint[12]), .I2(n25_adj_4516), 
            .I3(GND_net), .O(n29946));   // verilog/pwm.v(21[8:24])
    defparam i24880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24837_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n29350), 
            .O(n29903));
    defparam i24837_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25057_4_lut (.I0(n29948), .I1(n30074), .I2(n35), .I3(n29343), 
            .O(n30123));   // verilog/pwm.v(21[8:24])
    defparam i25057_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24900_4_lut (.I0(n29946), .I1(n29873), .I2(n25_adj_4516), 
            .I3(n29627), .O(n29966));   // verilog/pwm.v(21[8:24])
    defparam i24900_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i25061_4_lut (.I0(n29966), .I1(n30123), .I2(n35), .I3(n29903), 
            .O(n30127));   // verilog/pwm.v(21[8:24])
    defparam i25061_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25062_3_lut (.I0(n30127), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n30128));   // verilog/pwm.v(21[8:24])
    defparam i25062_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25060_3_lut (.I0(n30128), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n30126));   // verilog/pwm.v(21[8:24])
    defparam i25060_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24988_3_lut (.I0(n30126), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n30054));   // verilog/pwm.v(21[8:24])
    defparam i24988_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24989_3_lut (.I0(n30054), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n30055));   // verilog/pwm.v(21[8:24])
    defparam i24989_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11145_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n27156), 
            .I3(GND_net), .O(n14950));   // verilog/coms.v(127[12] 300[6])
    defparam i11145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11146_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n27156), 
            .I3(GND_net), .O(n14951));   // verilog/coms.v(127[12] 300[6])
    defparam i11146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11147_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n27156), 
            .I3(GND_net), .O(n14952));   // verilog/coms.v(127[12] 300[6])
    defparam i11147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11148_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n27156), 
            .I3(GND_net), .O(n14953));   // verilog/coms.v(127[12] 300[6])
    defparam i11148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11149_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n27156), 
            .I3(GND_net), .O(n14954));   // verilog/coms.v(127[12] 300[6])
    defparam i11149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11150_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n27156), 
            .I3(GND_net), .O(n14955));   // verilog/coms.v(127[12] 300[6])
    defparam i11150_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11151_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n27156), 
            .I3(GND_net), .O(n14956));   // verilog/coms.v(127[12] 300[6])
    defparam i11151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11152_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n10896), .I3(GND_net), .O(n14957));   // verilog/coms.v(127[12] 300[6])
    defparam i11152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11153_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n10896), .I3(GND_net), .O(n14958));   // verilog/coms.v(127[12] 300[6])
    defparam i11153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11154_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n10896), .I3(GND_net), .O(n14959));   // verilog/coms.v(127[12] 300[6])
    defparam i11154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11155_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n10896), .I3(GND_net), .O(n14960));   // verilog/coms.v(127[12] 300[6])
    defparam i11155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i7_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[6]), 
            .I3(encoder0_position[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i8_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[7]), 
            .I3(encoder0_position[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11156_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n10896), .I3(GND_net), .O(n14961));   // verilog/coms.v(127[12] 300[6])
    defparam i11156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11157_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n10896), .I3(GND_net), .O(n14962));   // verilog/coms.v(127[12] 300[6])
    defparam i11157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i9_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[8]), 
            .I3(encoder0_position[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i10_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[9]), 
            .I3(encoder0_position[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11158_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n10896), .I3(GND_net), .O(n14963));   // verilog/coms.v(127[12] 300[6])
    defparam i11158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11159_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n10896), .I3(GND_net), .O(n14964));   // verilog/coms.v(127[12] 300[6])
    defparam i11159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11160_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n10896), .I3(GND_net), .O(n14965));   // verilog/coms.v(127[12] 300[6])
    defparam i11160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11161_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n10896), .I3(GND_net), .O(n14966));   // verilog/coms.v(127[12] 300[6])
    defparam i11161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11162_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n10896), .I3(GND_net), .O(n14967));   // verilog/coms.v(127[12] 300[6])
    defparam i11162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11163_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n10896), .I3(GND_net), .O(n14968));   // verilog/coms.v(127[12] 300[6])
    defparam i11163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11164_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n10896), .I3(GND_net), .O(n14969));   // verilog/coms.v(127[12] 300[6])
    defparam i11164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11165_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n10896), .I3(GND_net), .O(n14970));   // verilog/coms.v(127[12] 300[6])
    defparam i11165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11166_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n10896), .I3(GND_net), .O(n14971));   // verilog/coms.v(127[12] 300[6])
    defparam i11166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11167_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n10896), .I3(GND_net), .O(n14972));   // verilog/coms.v(127[12] 300[6])
    defparam i11167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11168_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n10896), .I3(GND_net), .O(n14973));   // verilog/coms.v(127[12] 300[6])
    defparam i11168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11169_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n10896), .I3(GND_net), .O(n14974));   // verilog/coms.v(127[12] 300[6])
    defparam i11169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24888_3_lut (.I0(n30055), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n29954));   // verilog/pwm.v(21[8:24])
    defparam i24888_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11170_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n10896), .I3(GND_net), .O(n14975));   // verilog/coms.v(127[12] 300[6])
    defparam i11170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11171_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n10896), .I3(GND_net), .O(n14976));   // verilog/coms.v(127[12] 300[6])
    defparam i11171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11172_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n10896), .I3(GND_net), .O(n14977));   // verilog/coms.v(127[12] 300[6])
    defparam i11172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11173_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n10896), .I3(GND_net), .O(n14978));   // verilog/coms.v(127[12] 300[6])
    defparam i11173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11174_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n10896), .I3(GND_net), .O(n14979));   // verilog/coms.v(127[12] 300[6])
    defparam i11174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11175_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n10896), .I3(GND_net), .O(n14980));   // verilog/coms.v(127[12] 300[6])
    defparam i11175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11176_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n10896), .I3(GND_net), .O(n14981));   // verilog/coms.v(127[12] 300[6])
    defparam i11176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11012_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n1554), .I3(GND_net), .O(n14817));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11013_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n4137), .I3(GND_net), .O(n14818));   // verilog/coms.v(127[12] 300[6])
    defparam i11013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11015_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n18789), 
            .I3(n13556), .O(n14820));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11015_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i11016_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n18789), 
            .I3(n13551), .O(n14821));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11016_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_37_i11_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[10]), 
            .I3(encoder0_position[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11017_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n13556), 
            .O(n14822));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11017_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11018_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n13551), 
            .O(n14823));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11018_4_lut.LUT_INIT = 16'hccca;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_26[0]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_LUT4 i11177_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n10896), .I3(GND_net), .O(n14982));   // verilog/coms.v(127[12] 300[6])
    defparam i11177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11178_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n10896), .I3(GND_net), .O(n14983));   // verilog/coms.v(127[12] 300[6])
    defparam i11178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11179_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n10896), .I3(GND_net), .O(n14984));   // verilog/coms.v(127[12] 300[6])
    defparam i11179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11180_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n10896), .I3(GND_net), .O(n14985));   // verilog/coms.v(127[12] 300[6])
    defparam i11180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11181_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n10896), .I3(GND_net), .O(n14986));   // verilog/coms.v(127[12] 300[6])
    defparam i11181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11182_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n10896), .I3(GND_net), .O(n14987));   // verilog/coms.v(127[12] 300[6])
    defparam i11182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11183_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n10896), .I3(GND_net), .O(n14988));   // verilog/coms.v(127[12] 300[6])
    defparam i11183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11019_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4481), 
            .I3(n13556), .O(n14824));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11019_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11020_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4481), 
            .I3(n13551), .O(n14825));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11020_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11021_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4473), 
            .I3(n13556), .O(n14826));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11021_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11022_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14827));   // verilog/coms.v(127[12] 300[6])
    defparam i11022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11023_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n27156), 
            .I3(GND_net), .O(n14828));   // verilog/coms.v(127[12] 300[6])
    defparam i11023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11024_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n27156), 
            .I3(GND_net), .O(n14829));   // verilog/coms.v(127[12] 300[6])
    defparam i11024_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11025_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n4141), .I3(GND_net), .O(n14830));   // verilog/coms.v(127[12] 300[6])
    defparam i11025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11184_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n10896), .I3(GND_net), .O(n14989));   // verilog/coms.v(127[12] 300[6])
    defparam i11184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11185_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n10896), .I3(GND_net), .O(n14990));   // verilog/coms.v(127[12] 300[6])
    defparam i11185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11186_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n10896), .I3(GND_net), .O(n14991));   // verilog/coms.v(127[12] 300[6])
    defparam i11186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4463), .I3(n15_adj_4478), .O(motor_state_23__N_50[6]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11187_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n10896), .I3(GND_net), .O(n14992));   // verilog/coms.v(127[12] 300[6])
    defparam i11187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11188_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n10896), .I3(GND_net), .O(n14993));   // verilog/coms.v(127[12] 300[6])
    defparam i11188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11189_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n10896), .I3(GND_net), .O(n14994));   // verilog/coms.v(127[12] 300[6])
    defparam i11189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i12_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[11]), 
            .I3(encoder0_position[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11190_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n10896), .I3(GND_net), .O(n14995));   // verilog/coms.v(127[12] 300[6])
    defparam i11190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11191_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n10896), .I3(GND_net), .O(n14996));   // verilog/coms.v(127[12] 300[6])
    defparam i11191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11192_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n10896), .I3(GND_net), .O(n14997));   // verilog/coms.v(127[12] 300[6])
    defparam i11192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11193_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n10896), .I3(GND_net), .O(n14998));   // verilog/coms.v(127[12] 300[6])
    defparam i11193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11194_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n10896), .I3(GND_net), .O(n14999));   // verilog/coms.v(127[12] 300[6])
    defparam i11194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11195_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n10896), .I3(GND_net), .O(n15000));   // verilog/coms.v(127[12] 300[6])
    defparam i11195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i13_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[12]), 
            .I3(encoder0_position[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11196_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n10896), .I3(GND_net), .O(n15001));   // verilog/coms.v(127[12] 300[6])
    defparam i11196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11197_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n10896), .I3(GND_net), .O(n15002));   // verilog/coms.v(127[12] 300[6])
    defparam i11197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11198_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n10896), .I3(GND_net), .O(n15003));   // verilog/coms.v(127[12] 300[6])
    defparam i11198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11199_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n10896), .I3(GND_net), .O(n15004));   // verilog/coms.v(127[12] 300[6])
    defparam i11199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11200_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n10896), .I3(GND_net), .O(n15005));   // verilog/coms.v(127[12] 300[6])
    defparam i11200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i14_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[13]), 
            .I3(encoder0_position[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11201_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n10896), .I3(GND_net), .O(n15006));   // verilog/coms.v(127[12] 300[6])
    defparam i11201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11202_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n10896), .I3(GND_net), .O(n15007));   // verilog/coms.v(127[12] 300[6])
    defparam i11202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11203_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n10896), .I3(GND_net), .O(n15008));   // verilog/coms.v(127[12] 300[6])
    defparam i11203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11204_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n10896), .I3(GND_net), .O(n15009));   // verilog/coms.v(127[12] 300[6])
    defparam i11204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11205_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n10896), .I3(GND_net), .O(n15010));   // verilog/coms.v(127[12] 300[6])
    defparam i11205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11206_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n10896), .I3(GND_net), .O(n15011));   // verilog/coms.v(127[12] 300[6])
    defparam i11206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i15_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[14]), 
            .I3(encoder0_position[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11207_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n10896), .I3(GND_net), .O(n15012));   // verilog/coms.v(127[12] 300[6])
    defparam i11207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11208_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n10896), .I3(GND_net), .O(n15013));   // verilog/coms.v(127[12] 300[6])
    defparam i11208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11209_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n10896), .I3(GND_net), .O(n15014));   // verilog/coms.v(127[12] 300[6])
    defparam i11209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11210_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n10896), .I3(GND_net), .O(n15015));   // verilog/coms.v(127[12] 300[6])
    defparam i11210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11211_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n10896), .I3(GND_net), .O(n15016));   // verilog/coms.v(127[12] 300[6])
    defparam i11211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11212_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n10896), .I3(GND_net), .O(n15017));   // verilog/coms.v(127[12] 300[6])
    defparam i11212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11213_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n10896), .I3(GND_net), .O(n15018));   // verilog/coms.v(127[12] 300[6])
    defparam i11213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11214_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n10896), .I3(GND_net), .O(n15019));   // verilog/coms.v(127[12] 300[6])
    defparam i11214_3_lut.LUT_INIT = 16'hcaca;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4468, 
            quadB_debounced_adj_4469}), .n28236(n28236), .reg_B({reg_B_adj_4578}), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .VCC_net(VCC_net), .n14836(n14836), 
            .ENCODER1_B_c_0(ENCODER1_B_c_0), .n15348(n15348)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(193[15] 198[4])
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 mux_37_i16_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[15]), 
            .I3(encoder0_position[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i17_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[16]), 
            .I3(encoder0_position[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i18_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[17]), 
            .I3(encoder0_position[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11215_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n10896), .I3(GND_net), .O(n15020));   // verilog/coms.v(127[12] 300[6])
    defparam i11215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11216_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n10896), .I3(GND_net), .O(n15021));   // verilog/coms.v(127[12] 300[6])
    defparam i11216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11217_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n10896), .I3(GND_net), .O(n15022));   // verilog/coms.v(127[12] 300[6])
    defparam i11217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11218_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n10896), .I3(GND_net), .O(n15023));   // verilog/coms.v(127[12] 300[6])
    defparam i11218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11219_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n10896), .I3(GND_net), .O(n15024));   // verilog/coms.v(127[12] 300[6])
    defparam i11219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i19_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[18]), 
            .I3(encoder0_position[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11220_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n10896), .I3(GND_net), .O(n15025));   // verilog/coms.v(127[12] 300[6])
    defparam i11220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11221_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n10896), .I3(GND_net), .O(n15026));   // verilog/coms.v(127[12] 300[6])
    defparam i11221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11222_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n10896), .I3(GND_net), .O(n15027));   // verilog/coms.v(127[12] 300[6])
    defparam i11222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11223_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n10896), .I3(GND_net), .O(n15028));   // verilog/coms.v(127[12] 300[6])
    defparam i11223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11224_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n10896), .I3(GND_net), .O(n15029));   // verilog/coms.v(127[12] 300[6])
    defparam i11224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11225_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n10896), .I3(GND_net), .O(n15030));   // verilog/coms.v(127[12] 300[6])
    defparam i11225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11226_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n10896), .I3(GND_net), .O(n15031));   // verilog/coms.v(127[12] 300[6])
    defparam i11226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11227_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n10896), .I3(GND_net), .O(n15032));   // verilog/coms.v(127[12] 300[6])
    defparam i11227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11228_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n10896), .I3(GND_net), .O(n15033));   // verilog/coms.v(127[12] 300[6])
    defparam i11228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11229_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n10896), .I3(GND_net), .O(n15034));   // verilog/coms.v(127[12] 300[6])
    defparam i11229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11230_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n10896), .I3(GND_net), .O(n15035));   // verilog/coms.v(127[12] 300[6])
    defparam i11230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11231_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n10896), .I3(GND_net), .O(n15036));   // verilog/coms.v(127[12] 300[6])
    defparam i11231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11232_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n10896), 
            .I3(GND_net), .O(n15037));   // verilog/coms.v(127[12] 300[6])
    defparam i11232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11233_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n10896), 
            .I3(GND_net), .O(n15038));   // verilog/coms.v(127[12] 300[6])
    defparam i11233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11234_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n10896), 
            .I3(GND_net), .O(n15039));   // verilog/coms.v(127[12] 300[6])
    defparam i11234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11235_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n10896), 
            .I3(GND_net), .O(n15040));   // verilog/coms.v(127[12] 300[6])
    defparam i11235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11236_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n10896), 
            .I3(GND_net), .O(n15041));   // verilog/coms.v(127[12] 300[6])
    defparam i11236_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i11237_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n10896), 
            .I3(GND_net), .O(n15042));   // verilog/coms.v(127[12] 300[6])
    defparam i11237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11238_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n10896), 
            .I3(GND_net), .O(n15043));   // verilog/coms.v(127[12] 300[6])
    defparam i11238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11239_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n10896), 
            .I3(GND_net), .O(n15044));   // verilog/coms.v(127[12] 300[6])
    defparam i11239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11240_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n10896), 
            .I3(GND_net), .O(n15045));   // verilog/coms.v(127[12] 300[6])
    defparam i11240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11241_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n10896), 
            .I3(GND_net), .O(n15046));   // verilog/coms.v(127[12] 300[6])
    defparam i11241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i20_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[19]), 
            .I3(encoder0_position[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11242_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n10896), 
            .I3(GND_net), .O(n15047));   // verilog/coms.v(127[12] 300[6])
    defparam i11242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11243_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n10896), 
            .I3(GND_net), .O(n15048));   // verilog/coms.v(127[12] 300[6])
    defparam i11243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_4464), .I3(control_mode[2]), .O(n13399));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11304_3_lut_4_lut (.I0(\data_out_frame[27] [0]), .I1(n24343), 
            .I2(n26399), .I3(n14641), .O(n15109));   // verilog/coms.v(127[12] 300[6])
    defparam i11304_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i11244_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n10896), 
            .I3(GND_net), .O(n15049));   // verilog/coms.v(127[12] 300[6])
    defparam i11244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11245_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n10896), 
            .I3(GND_net), .O(n15050));   // verilog/coms.v(127[12] 300[6])
    defparam i11245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11246_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n10896), 
            .I3(GND_net), .O(n15051));   // verilog/coms.v(127[12] 300[6])
    defparam i11246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11247_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n10896), 
            .I3(GND_net), .O(n15052));   // verilog/coms.v(127[12] 300[6])
    defparam i11247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11248_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n10896), 
            .I3(GND_net), .O(n15053));   // verilog/coms.v(127[12] 300[6])
    defparam i11248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11249_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n10896), 
            .I3(GND_net), .O(n15054));   // verilog/coms.v(127[12] 300[6])
    defparam i11249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11250_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n10896), 
            .I3(GND_net), .O(n15055));   // verilog/coms.v(127[12] 300[6])
    defparam i11250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11251_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n10896), 
            .I3(GND_net), .O(n15056));   // verilog/coms.v(127[12] 300[6])
    defparam i11251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11252_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n10896), 
            .I3(GND_net), .O(n15057));   // verilog/coms.v(127[12] 300[6])
    defparam i11252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11253_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n10896), 
            .I3(GND_net), .O(n15058));   // verilog/coms.v(127[12] 300[6])
    defparam i11253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11254_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n10896), 
            .I3(GND_net), .O(n15059));   // verilog/coms.v(127[12] 300[6])
    defparam i11254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11255_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n10896), 
            .I3(GND_net), .O(n15060));   // verilog/coms.v(127[12] 300[6])
    defparam i11255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11256_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n10896), .I3(GND_net), .O(n15061));   // verilog/coms.v(127[12] 300[6])
    defparam i11256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11257_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n10896), .I3(GND_net), .O(n15062));   // verilog/coms.v(127[12] 300[6])
    defparam i11257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11258_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n10896), .I3(GND_net), .O(n15063));   // verilog/coms.v(127[12] 300[6])
    defparam i11258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11259_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n10896), .I3(GND_net), .O(n15064));   // verilog/coms.v(127[12] 300[6])
    defparam i11259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11260_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n10896), .I3(GND_net), .O(n15065));   // verilog/coms.v(127[12] 300[6])
    defparam i11260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i21_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[20]), 
            .I3(encoder0_position[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11261_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n10896), .I3(GND_net), .O(n15066));   // verilog/coms.v(127[12] 300[6])
    defparam i11261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11262_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n10896), .I3(GND_net), .O(n15067));   // verilog/coms.v(127[12] 300[6])
    defparam i11262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11263_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n10896), .I3(GND_net), .O(n15068));   // verilog/coms.v(127[12] 300[6])
    defparam i11263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11264_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n10896), .I3(GND_net), .O(n15069));   // verilog/coms.v(127[12] 300[6])
    defparam i11264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11265_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n10896), .I3(GND_net), .O(n15070));   // verilog/coms.v(127[12] 300[6])
    defparam i11265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11266_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n10896), .I3(GND_net), .O(n15071));   // verilog/coms.v(127[12] 300[6])
    defparam i11266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11267_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n10896), .I3(GND_net), .O(n15072));   // verilog/coms.v(127[12] 300[6])
    defparam i11267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11268_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n10896), .I3(GND_net), .O(n15073));   // verilog/coms.v(127[12] 300[6])
    defparam i11268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11269_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n10896), .I3(GND_net), .O(n15074));   // verilog/coms.v(127[12] 300[6])
    defparam i11269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11270_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n10896), .I3(GND_net), .O(n15075));   // verilog/coms.v(127[12] 300[6])
    defparam i11270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i22_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[21]), 
            .I3(encoder0_position[21]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i23_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[22]), 
            .I3(encoder0_position[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11271_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n10896), .I3(GND_net), .O(n15076));   // verilog/coms.v(127[12] 300[6])
    defparam i11271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11272_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n10896), .I3(GND_net), .O(n15077));   // verilog/coms.v(127[12] 300[6])
    defparam i11272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11274_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n10896), .I3(GND_net), .O(n15079));   // verilog/coms.v(127[12] 300[6])
    defparam i11274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11275_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n10896), .I3(GND_net), .O(n15080));   // verilog/coms.v(127[12] 300[6])
    defparam i11275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11276_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n10896), .I3(GND_net), .O(n15081));   // verilog/coms.v(127[12] 300[6])
    defparam i11276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11277_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n10896), .I3(GND_net), .O(n15082));   // verilog/coms.v(127[12] 300[6])
    defparam i11277_3_lut.LUT_INIT = 16'hcaca;
    motorControl control (.GND_net(GND_net), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), 
            .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .IntegralLimit({IntegralLimit}), 
            .PWMLimit({PWMLimit}), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), 
            .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
            .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
            .\Ki[15] (Ki[15]), .duty({duty}), .n30261(n30261), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz), .setpoint({setpoint}), .motor_state({motor_state})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(170[16] 182[4])
    SB_LUT4 i11278_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n10896), .I3(GND_net), .O(n15083));   // verilog/coms.v(127[12] 300[6])
    defparam i11278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11279_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n10896), .I3(GND_net), .O(n15084));   // verilog/coms.v(127[12] 300[6])
    defparam i11279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i24_3_lut_4_lut (.I0(n13399), .I1(control_mode[1]), .I2(motor_state_23__N_50[23]), 
            .I3(encoder0_position[23]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11280_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n10896), .I3(GND_net), .O(n15085));   // verilog/coms.v(127[12] 300[6])
    defparam i11280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11281_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n10896), .I3(GND_net), .O(n15086));   // verilog/coms.v(127[12] 300[6])
    defparam i11281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11282_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n10896), .I3(GND_net), .O(n15087));   // verilog/coms.v(127[12] 300[6])
    defparam i11282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11283_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n10896), .I3(GND_net), .O(n15088));   // verilog/coms.v(127[12] 300[6])
    defparam i11283_3_lut.LUT_INIT = 16'hcaca;
    pwm PWM (.n29954(n29954), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n13407(n13407), .GND_net(GND_net), .n13405(n13405), .\pwm_counter[6] (pwm_counter[6]), 
        .\pwm_counter[8] (pwm_counter[8]), .\pwm_counter[7] (pwm_counter[7]), 
        .\pwm_counter[13] (pwm_counter[13]), .\pwm_counter[10] (pwm_counter[10]), 
        .\pwm_counter[9] (pwm_counter[9]), .\pwm_counter[17] (pwm_counter[17]), 
        .\pwm_counter[22] (pwm_counter[22]), .\pwm_counter[14] (pwm_counter[14]), 
        .\pwm_counter[18] (pwm_counter[18]), .\pwm_counter[21] (pwm_counter[21]), 
        .\pwm_counter[16] (pwm_counter[16]), .\pwm_counter[12] (pwm_counter[12]), 
        .\pwm_counter[15] (pwm_counter[15]), .\pwm_counter[19] (pwm_counter[19]), 
        .\pwm_counter[11] (pwm_counter[11]), .\pwm_counter[20] (pwm_counter[20]), 
        .\pwm_counter[31] (pwm_counter[31]), .\pwm_counter[0] (pwm_counter[0]), 
        .\pwm_counter[5] (pwm_counter[5]), .\pwm_counter[4] (pwm_counter[4]), 
        .\pwm_counter[3] (pwm_counter[3]), .\pwm_counter[2] (pwm_counter[2]), 
        .\pwm_counter[1] (pwm_counter[1])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(90[6] 95[3])
    coms neopxl_color_23__I_0 (.GND_net(GND_net), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .rx_data({rx_data}), .setpoint({setpoint}), .clk32MHz(clk32MHz), 
         .n14885(n14885), .IntegralLimit({IntegralLimit}), .n14884(n14884), 
         .n14883(n14883), .n10896(n10896), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .n4141(n4141), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[20] ({\data_out_frame[20] [7:2], 
         Open_0, \data_out_frame[20] [0]}), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .n14882(n14882), .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n14881(n14881), .n14880(n14880), .n14879(n14879), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n14878(n14878), .\data_in_frame[4] ({\data_in_frame[4] }), .n14877(n14877), 
         .n14876(n14876), .rx_data_ready(rx_data_ready), .n14875(n14875), 
         .n14874(n14874), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n14873(n14873), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n2252(n2252), .\data_in[1] ({\data_in[1] }), .\data_in[0] ({\data_in[0] }), 
         .\data_in[2] ({\data_in[2] }), .\data_in[3] ({\data_in[3] }), .n63(n63), 
         .n3(n3_adj_4521), .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\FRAME_MATCHER.state_31__N_2380[2] (\FRAME_MATCHER.state_31__N_2380 [2]), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .n4137(n4137), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[27][0] (\data_out_frame[27] [0]), .n4(n4_adj_4467), 
         .tx_active(tx_active), .n14641(n14641), .n24343(n24343), .n1(n1), 
         .DE_c(DE_c), .n26748(n26748), .n7(n7_adj_4466), .n7_adj_3(n7_adj_4518), 
         .LED_c(LED_c), .n5(n5_adj_4517), .n26399(n26399), .n14833(n14833), 
         .PWMLimit({PWMLimit}), .n14832(n14832), .control_mode({control_mode}), 
         .n28285(n28285), .n30820(n30820), .n15337(n15337), .n15336(n15336), 
         .n15335(n15335), .n15334(n15334), .n15333(n15333), .n15332(n15332), 
         .n15331(n15331), .n15330(n15330), .n15329(n15329), .n15328(n15328), 
         .n15327(n15327), .n15326(n15326), .n15325(n15325), .n15324(n15324), 
         .n15323(n15323), .n15322(n15322), .n15321(n15321), .n15320(n15320), 
         .n15319(n15319), .n15318(n15318), .n15317(n15317), .n15316(n15316), 
         .n15315(n15315), .n15314(n15314), .n15313(n15313), .n15312(n15312), 
         .n15311(n15311), .n15310(n15310), .n15309(n15309), .n15308(n15308), 
         .n15132(n15132), .neopxl_color({neopxl_color}), .n15131(n15131), 
         .n15130(n15130), .n15129(n15129), .n15128(n15128), .n15127(n15127), 
         .n15126(n15126), .n15125(n15125), .n15124(n15124), .n15123(n15123), 
         .n15122(n15122), .n15121(n15121), .n15120(n15120), .n15119(n15119), 
         .n15118(n15118), .n15117(n15117), .n15116(n15116), .n15115(n15115), 
         .n15114(n15114), .n15113(n15113), .n15112(n15112), .n15111(n15111), 
         .n15110(n15110), .n15109(n15109), .n15108(n15108), .n15107(n15107), 
         .n15106(n15106), .n15105(n15105), .n15104(n15104), .n15103(n15103), 
         .n15102(n15102), .n15101(n15101), .n15100(n15100), .n15099(n15099), 
         .n15098(n15098), .n15097(n15097), .n15096(n15096), .n15095(n15095), 
         .n15094(n15094), .n15093(n15093), .n15092(n15092), .n15091(n15091), 
         .n15090(n15090), .n15089(n15089), .n15088(n15088), .n15087(n15087), 
         .n15086(n15086), .n15085(n15085), .n15084(n15084), .n15083(n15083), 
         .n15082(n15082), .n15081(n15081), .n15080(n15080), .n15079(n15079), 
         .n15077(n15077), .n15076(n15076), .n15075(n15075), .n15074(n15074), 
         .n15073(n15073), .n15072(n15072), .n15071(n15071), .n15070(n15070), 
         .n15069(n15069), .n15068(n15068), .n15067(n15067), .n15066(n15066), 
         .n15065(n15065), .n15064(n15064), .n15063(n15063), .n15062(n15062), 
         .n15061(n15061), .n15060(n15060), .n15059(n15059), .n15058(n15058), 
         .n15057(n15057), .n15056(n15056), .n15055(n15055), .n15054(n15054), 
         .n15053(n15053), .n15052(n15052), .n15051(n15051), .n15050(n15050), 
         .n15049(n15049), .n15048(n15048), .n15047(n15047), .n15046(n15046), 
         .n15045(n15045), .n15044(n15044), .n15043(n15043), .n15042(n15042), 
         .n15041(n15041), .n15040(n15040), .n15039(n15039), .n15038(n15038), 
         .n15037(n15037), .n15036(n15036), .n15035(n15035), .n15034(n15034), 
         .n15033(n15033), .n15032(n15032), .n15031(n15031), .n15030(n15030), 
         .n15029(n15029), .n15028(n15028), .n15027(n15027), .n15026(n15026), 
         .n15025(n15025), .n15024(n15024), .n15023(n15023), .n15022(n15022), 
         .n15021(n15021), .n15020(n15020), .n27156(n27156), .n15019(n15019), 
         .n15018(n15018), .n15017(n15017), .n15016(n15016), .n15015(n15015), 
         .n15014(n15014), .n15013(n15013), .n15012(n15012), .n15011(n15011), 
         .n15010(n15010), .n15009(n15009), .n15008(n15008), .n15007(n15007), 
         .n15006(n15006), .n15005(n15005), .n15004(n15004), .n15003(n15003), 
         .n15002(n15002), .n15001(n15001), .n15000(n15000), .n14999(n14999), 
         .n14998(n14998), .n14997(n14997), .n14996(n14996), .n14995(n14995), 
         .n14994(n14994), .n14993(n14993), .n14992(n14992), .n14991(n14991), 
         .n14990(n14990), .n14989(n14989), .n14830(n14830), .n14829(n14829), 
         .\Ki[0] (Ki[0]), .n14828(n14828), .\Kp[0] (Kp[0]), .n14827(n14827), 
         .n14988(n14988), .n14987(n14987), .n14986(n14986), .n14985(n14985), 
         .n14984(n14984), .n14983(n14983), .n14982(n14982), .n14818(n14818), 
         .n14981(n14981), .n14980(n14980), .n14979(n14979), .n14978(n14978), 
         .n14977(n14977), .n14976(n14976), .n14975(n14975), .n14974(n14974), 
         .n14973(n14973), .n14972(n14972), .n14971(n14971), .n14970(n14970), 
         .n14969(n14969), .n14968(n14968), .n14967(n14967), .n14966(n14966), 
         .n14965(n14965), .n14964(n14964), .n14963(n14963), .n14962(n14962), 
         .n14961(n14961), .n14960(n14960), .n14959(n14959), .n14958(n14958), 
         .n14957(n14957), .n14956(n14956), .\Ki[15] (Ki[15]), .n14955(n14955), 
         .\Ki[14] (Ki[14]), .n14954(n14954), .\Ki[13] (Ki[13]), .n14953(n14953), 
         .\Ki[12] (Ki[12]), .n14952(n14952), .\Ki[11] (Ki[11]), .n14951(n14951), 
         .\Ki[10] (Ki[10]), .n14950(n14950), .\Ki[9] (Ki[9]), .n14949(n14949), 
         .\Ki[8] (Ki[8]), .n14948(n14948), .\Ki[7] (Ki[7]), .n14947(n14947), 
         .\Ki[6] (Ki[6]), .n14946(n14946), .\Ki[5] (Ki[5]), .n14945(n14945), 
         .\Ki[4] (Ki[4]), .n14944(n14944), .\Ki[3] (Ki[3]), .n14943(n14943), 
         .\Ki[2] (Ki[2]), .n14942(n14942), .\Ki[1] (Ki[1]), .n14941(n14941), 
         .\Kp[15] (Kp[15]), .n14940(n14940), .\Kp[14] (Kp[14]), .n14939(n14939), 
         .\Kp[13] (Kp[13]), .n14938(n14938), .\Kp[12] (Kp[12]), .n14937(n14937), 
         .\Kp[11] (Kp[11]), .n14936(n14936), .\Kp[10] (Kp[10]), .n14935(n14935), 
         .\Kp[9] (Kp[9]), .n14934(n14934), .\Kp[8] (Kp[8]), .n14933(n14933), 
         .\Kp[7] (Kp[7]), .n14932(n14932), .\Kp[6] (Kp[6]), .n14931(n14931), 
         .\Kp[5] (Kp[5]), .n14930(n14930), .\Kp[4] (Kp[4]), .n14929(n14929), 
         .\Kp[3] (Kp[3]), .n14928(n14928), .\Kp[2] (Kp[2]), .n14927(n14927), 
         .\Kp[1] (Kp[1]), .n14926(n14926), .n14925(n14925), .n14924(n14924), 
         .n14923(n14923), .n14922(n14922), .n14921(n14921), .n14920(n14920), 
         .n14919(n14919), .n14918(n14918), .n14917(n14917), .n14916(n14916), 
         .n14915(n14915), .n14914(n14914), .n14913(n14913), .n14912(n14912), 
         .n14911(n14911), .n14910(n14910), .n14909(n14909), .n14908(n14908), 
         .n14907(n14907), .n14906(n14906), .n14905(n14905), .n14904(n14904), 
         .n14903(n14903), .n14902(n14902), .n14901(n14901), .\displacement[1] (displacement[1]), 
         .n14900(n14900), .n14899(n14899), .n14898(n14898), .n14897(n14897), 
         .n14896(n14896), .n14895(n14895), .n14894(n14894), .n14893(n14893), 
         .n14892(n14892), .n14891(n14891), .n14890(n14890), .n14889(n14889), 
         .n14888(n14888), .n14887(n14887), .n14886(n14886), .n26856(n26856), 
         .n26880(n26880), .r_SM_Main({r_SM_Main_adj_4567}), .\r_SM_Main_2__N_3333[1] (r_SM_Main_2__N_3333[1]), 
         .tx_o(tx_o), .n14872(n14872), .VCC_net(VCC_net), .\r_Bit_Index[0] (r_Bit_Index_adj_4569[0]), 
         .n7375(n7375), .n14835(n14835), .n4_adj_4(n4_adj_4520), .n30875(n30875), 
         .tx_enable(tx_enable), .n14672(n14672), .n14766(n14766), .\r_SM_Main_2__N_3262[2] (r_SM_Main_2__N_3262[2]), 
         .r_SM_Main_adj_12({r_SM_Main}), .n26029(n26029), .r_Rx_Data(r_Rx_Data), 
         .RX_N_2(RX_N_2), .\r_Bit_Index[0]_adj_8 (r_Bit_Index[0]), .n13551(n13551), 
         .n4_adj_9(n4_adj_4473), .n15342(n15342), .n25777(n25777), .n15346(n15346), 
         .n18789(n18789), .n4_adj_10(n4), .n4_adj_11(n4_adj_4481), .n13556(n13556), 
         .n14826(n14826), .n14825(n14825), .n14824(n14824), .n14823(n14823), 
         .n14822(n14822), .n14821(n14821), .n14820(n14820)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(137[8] 160[4])
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, clk32MHz, data_o, 
            GND_net, n28241, reg_B, VCC_net, n14834, ENCODER0_B_c_0, 
            n15347, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input clk32MHz;
    output [1:0]data_o;
    input GND_net;
    output n28241;
    output [1:0]reg_B;
    input VCC_net;
    input n14834;
    input ENCODER0_B_c_0;
    input n15347;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2472;
    
    wire count_enable, B_delayed, A_delayed, count_direction, n2468, 
        n22090, n22089, n22088, n22087, n22086, n22085, n22084, 
        n22083, n22082, n22081, n22080, n22079, n22078, n22077, 
        n22076, n22075, n22074, n22073, n22072, n22071, n22070, 
        n22069, n22068, n22067;
    
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2472[23]));   // quad.v(35[10] 41[6])
    SB_LUT4 i843_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2468));   // quad.v(37[5] 40[8])
    defparam i843_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_552_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2468), 
            .I3(n22090), .O(n2472[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_552_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2468), 
            .I3(n22089), .O(n2472[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_24 (.CI(n22089), .I0(encoder0_position[22]), .I1(n2468), 
            .CO(n22090));
    SB_LUT4 add_552_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2468), 
            .I3(n22088), .O(n2472[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_23 (.CI(n22088), .I0(encoder0_position[21]), .I1(n2468), 
            .CO(n22089));
    SB_LUT4 add_552_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2468), 
            .I3(n22087), .O(n2472[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_22 (.CI(n22087), .I0(encoder0_position[20]), .I1(n2468), 
            .CO(n22088));
    SB_LUT4 add_552_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2468), 
            .I3(n22086), .O(n2472[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_21 (.CI(n22086), .I0(encoder0_position[19]), .I1(n2468), 
            .CO(n22087));
    SB_LUT4 add_552_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2468), 
            .I3(n22085), .O(n2472[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_20 (.CI(n22085), .I0(encoder0_position[18]), .I1(n2468), 
            .CO(n22086));
    SB_LUT4 add_552_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2468), 
            .I3(n22084), .O(n2472[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_19 (.CI(n22084), .I0(encoder0_position[17]), .I1(n2468), 
            .CO(n22085));
    SB_LUT4 add_552_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2468), 
            .I3(n22083), .O(n2472[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_18 (.CI(n22083), .I0(encoder0_position[16]), .I1(n2468), 
            .CO(n22084));
    SB_LUT4 add_552_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2468), 
            .I3(n22082), .O(n2472[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_17 (.CI(n22082), .I0(encoder0_position[15]), .I1(n2468), 
            .CO(n22083));
    SB_LUT4 add_552_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2468), 
            .I3(n22081), .O(n2472[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_16 (.CI(n22081), .I0(encoder0_position[14]), .I1(n2468), 
            .CO(n22082));
    SB_LUT4 add_552_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2468), 
            .I3(n22080), .O(n2472[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_15 (.CI(n22080), .I0(encoder0_position[13]), .I1(n2468), 
            .CO(n22081));
    SB_LUT4 add_552_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2468), 
            .I3(n22079), .O(n2472[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_14 (.CI(n22079), .I0(encoder0_position[12]), .I1(n2468), 
            .CO(n22080));
    SB_LUT4 add_552_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2468), 
            .I3(n22078), .O(n2472[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_13 (.CI(n22078), .I0(encoder0_position[11]), .I1(n2468), 
            .CO(n22079));
    SB_LUT4 add_552_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2468), 
            .I3(n22077), .O(n2472[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_12 (.CI(n22077), .I0(encoder0_position[10]), .I1(n2468), 
            .CO(n22078));
    SB_LUT4 add_552_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2468), 
            .I3(n22076), .O(n2472[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_11 (.CI(n22076), .I0(encoder0_position[9]), .I1(n2468), 
            .CO(n22077));
    SB_LUT4 add_552_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2468), 
            .I3(n22075), .O(n2472[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_10 (.CI(n22075), .I0(encoder0_position[8]), .I1(n2468), 
            .CO(n22076));
    SB_LUT4 add_552_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2468), 
            .I3(n22074), .O(n2472[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_9 (.CI(n22074), .I0(encoder0_position[7]), .I1(n2468), 
            .CO(n22075));
    SB_LUT4 add_552_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2468), 
            .I3(n22073), .O(n2472[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_8 (.CI(n22073), .I0(encoder0_position[6]), .I1(n2468), 
            .CO(n22074));
    SB_LUT4 add_552_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2468), 
            .I3(n22072), .O(n2472[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_7 (.CI(n22072), .I0(encoder0_position[5]), .I1(n2468), 
            .CO(n22073));
    SB_LUT4 add_552_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2468), 
            .I3(n22071), .O(n2472[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_6 (.CI(n22071), .I0(encoder0_position[4]), .I1(n2468), 
            .CO(n22072));
    SB_LUT4 add_552_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2468), 
            .I3(n22070), .O(n2472[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_5 (.CI(n22070), .I0(encoder0_position[3]), .I1(n2468), 
            .CO(n22071));
    SB_LUT4 add_552_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2468), 
            .I3(n22069), .O(n2472[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_4 (.CI(n22069), .I0(encoder0_position[2]), .I1(n2468), 
            .CO(n22070));
    SB_LUT4 add_552_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2468), 
            .I3(n22068), .O(n2472[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_3 (.CI(n22068), .I0(encoder0_position[1]), .I1(n2468), 
            .CO(n22069));
    SB_LUT4 add_552_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n22067), .O(n2472[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_552_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_552_2 (.CI(n22067), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n22068));
    SB_CARRY add_552_1 (.CI(GND_net), .I0(n2468), .I1(n2468), .CO(n22067));
    \grp_debouncer(2,100)_U0  debounce (.n28241(n28241), .reg_B({reg_B}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .n14834(n14834), .data_o({data_o}), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .n15347(n15347), .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (n28241, reg_B, GND_net, clk32MHz, 
            VCC_net, n14834, data_o, ENCODER0_B_c_0, n15347, ENCODER0_A_c_1);
    output n28241;
    output [1:0]reg_B;
    input GND_net;
    input clk32MHz;
    input VCC_net;
    input n14834;
    output [1:0]data_o;
    input ENCODER0_B_c_0;
    input n15347;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3576;
    wire [6:0]n33;
    
    wire n22430, n22429, n22428, n22427, n22426, n22425;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n28241));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n28241), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1128__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1128_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n22430), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1128_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n22429), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1128_add_4_7 (.CI(n22429), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n22430));
    SB_LUT4 cnt_reg_1128_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n22428), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1128_add_4_6 (.CI(n22428), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n22429));
    SB_LUT4 cnt_reg_1128_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n22427), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1128_add_4_5 (.CI(n22427), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n22428));
    SB_LUT4 cnt_reg_1128_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n22426), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1128_add_4_4 (.CI(n22426), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n22427));
    SB_LUT4 cnt_reg_1128_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n22425), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1128_add_4_3 (.CI(n22425), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n22426));
    SB_LUT4 cnt_reg_1128_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1128_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1128_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n22425));
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n14834));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n15347));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1128__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1128__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1128__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1128__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1128__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1128__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (GND_net, clk32MHz, n26858, n28, \state[0] , \state[1] , 
            \one_wire_N_399[11] , n1554, timer, \neo_pixel_transmitter.t0 , 
            VCC_net, n20822, n29233, n14869, n14868, n4, neopxl_color, 
            n14867, n14866, n29210, n14865, n14864, n14863, n14862, 
            n14861, n14860, n14859, n14858, n14857, n14856, n14855, 
            n14854, n14853, n14852, n14851, n14850, n14849, n14848, 
            n14847, n14846, n14845, n14844, n14843, n14842, n14841, 
            n14840, n14839, n12, n25063, LED_c, n14817, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk32MHz;
    output n26858;
    output n28;
    output \state[0] ;
    output \state[1] ;
    output \one_wire_N_399[11] ;
    output n1554;
    output [31:0]timer;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input VCC_net;
    output n20822;
    output n29233;
    input n14869;
    input n14868;
    output n4;
    input [23:0]neopxl_color;
    input n14867;
    input n14866;
    output n29210;
    input n14865;
    input n14864;
    input n14863;
    input n14862;
    input n14861;
    input n14860;
    input n14859;
    input n14858;
    input n14857;
    input n14856;
    input n14855;
    input n14854;
    input n14853;
    input n14852;
    input n14851;
    input n14850;
    input n14849;
    input n14848;
    input n14847;
    input n14846;
    input n14845;
    input n14844;
    input n14843;
    input n14842;
    input n14841;
    input n14840;
    input n14839;
    input n12;
    input n25063;
    input LED_c;
    input n14817;
    output NEOPXL_c;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n22065, n1995, n2027, n22066, n2126, n30260, \neo_pixel_transmitter.done_N_456 , 
        n27007, \neo_pixel_transmitter.done , n64, start, n2095, n1996, 
        n22064, n22139;
    wire [31:0]n1;
    
    wire n22140;
    wire [31:0]one_wire_N_399;
    
    wire n22138, n2693, n2704, n28_adj_4305, n2699, n2706, n2694, 
        n2691, n38;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n2709, n19275, n2701, n2696, n2697, n36, n2700, n2705, 
        n42, n2702, n2690, n2689, n2708, n40, n2687, n2703, 
        n2695, n41, n2688, n2698, n2692, n2707, n39, n2720, 
        n2819, n30265;
    wire [31:0]n255;
    
    wire n14635, n14745, n2491, n2504, n24, n2496, n2505, n2500, 
        n2499, n34, n2497, n2509, n22, n2490, n2494, n38_adj_4306, 
        n2501, n2502, n2506, n2492, n36_adj_4307, n2495, n2498, 
        n2493, n37, n2507, n2508, n2503, n2489, n35, n2522, 
        n2621, n30267, n2798, n2804, n2791, n2795, n40_adj_4308, 
        n2796, n2793, n2788, n2808, n38_adj_4309, n2789, n2800, 
        n2803, n2805, n39_adj_4310, n2792, n2787, n2801, n2799, 
        n37_adj_4311, n2786, n2797, n34_adj_4312, n2096, n1997, 
        n22063, n2794, n2806, n2807, n2790, n42_adj_4313, n46, 
        n2802, n2809, n33_adj_4314, n2918, n30264, n2907, n2909, 
        n33_adj_4315, n2900, n2891, n2897, n2888, n41_adj_4316, 
        n2906, n2887, n2892, n38_adj_4317, n2896, n2885, n2905, 
        n2902, n43, n2899, n2890, n2898, n2908, n40_adj_4318, 
        n2889, n2901, n46_adj_4319, n2886, n2894, n2895, n2903, 
        n39_adj_4320, n2904, n2893, n47, n3017, n30263, n3209, 
        n19339, n35_adj_4321, n11, n29, n51, n48, n37_adj_4322, 
        n23, n53, n39_adj_4323, n46_adj_4324, n27, n57, n63, n43_adj_4325, 
        n47_adj_4326, n25, n33_adj_4327, n47_adj_4328, n61, n45, 
        n59, n17, n15, n55, n44, n31_adj_4329, n41_adj_4330, n49, 
        n43_adj_4331, n54, n45_adj_4332, n13, n19, n21, n49_adj_4333, 
        n23391, n23679, n3004, n2989, n2990, n3007, n40_adj_4334, 
        n3006, n2984, n2988, n2986, n44_adj_4335, n3008, n3003, 
        n2994, n3002, n42_adj_4336, n2999, n3000, n2992, n2997, 
        n43_adj_4337, n2996, n2985, n2995, n2987, n41_adj_4338, 
        n3001, n2993, n38_adj_4339, n2998, n2991, n46_adj_4340, 
        n50, n3005, n3009, n37_adj_4341, n3116, n30262, n2192, 
        n2093, n23164, n2193, n2094, n23163, n2194, n23162, n2195, 
        n23161, n2196, n2097, n23160, n2197, n2098, n23159, n2198, 
        n2099, n23158, n2199, n2100, n23157, n2200, n2101, n23156, 
        n2201, n2102, n23155, n2202, n2103, n23154, n2203, n2104, 
        n23153, n2204, n2105, n23152, n2205, n2106, n23151, n2206, 
        n2107, n23150, n2207, n2108, n23149, n2208, n2109, n23148, 
        n2209, n1998, n22062, n26, n21916, n3102, n3090, n3103, 
        n3085, n42_adj_4342, n3089, n3094, n3101, n3098, n46_adj_4343, 
        n3099, n3091, n3106, n3100, n44_adj_4344, n3097, n3088, 
        n3104, n3092, n45_adj_4345, n3105, n3083, n3093, n3096, 
        n43_adj_4346, n3108, n3109, n40_adj_4347, n3107, n3087, 
        n3086, n48_adj_4348, n52, n3095, n3084, n39_adj_4349, n30, 
        n21924, n30259, n2591, n2608, n2601, n2605, n36_adj_4350, 
        n2606, n2609, n25_adj_4351, n2593, n2596, n2600, n2590, 
        n34_adj_4352, n2594, n2589, n40_adj_4353, n2602, n2588, 
        n2604, n2607, n38_adj_4354, n2598, n2603, n39_adj_4355, 
        n2592, n2597, n2595, n2599, n37_adj_4356, n30266, n1999, 
        n22061, n28_adj_4357, n2000, n22060, n29_adj_4358, n27_adj_4359, 
        n2001, n22059, n1205, n1206, n1204, n1207, n14, n1203, 
        n1209, n9, n1202, n1208, n1235, n21917, n2002, n22058, 
        n1136, n30273, n21925, n2003, n22057, n1109, n19291, n1105, 
        n1103, n1108, n12_c, n1107, n1106, n1104, n2004, n22056, 
        n2005, n22055, n110, n2006, n22054, n2007, n22053, n2008, 
        n22052, n1037, n30272, n2;
    wire [31:0]n971;
    
    wire n1007, n1006, n906, n1005, n1009, n12133, n1008, n26828, 
        n14692, n8, n905, n28384, n6, n2009, n22051, n21923, 
        n4_c, n21922, n21944, n22661, n22660, n22659, n22658, 
        n22657, n22656, n22655, n22654, n22653, n21915, n46_adj_4360, 
        n44_adj_4361, n45_adj_4362, n43_adj_4363, n42_adj_4364, n41_adj_4365, 
        n52_adj_4366, n47_adj_4367, n24472, n73, n7, n86, n20817, 
        n83, n29305, n34_adj_4368, n22652, n22651, n22650, n22649, 
        n22648, n22647, n22646, n22645, n22644, n22643, n22642, 
        n22641, n22640, n22639, n22638, n22637, n22636, n22635, 
        n22634, n22633, n22632, n22631, n22630, n22629, n22628, 
        n29304, n21943, n22627, n22626, n22625, n22624, n22623, 
        n22622, n22621, n22620, n22619, n22618, n22617, n22616, 
        n22615, n22614, n22613, n22612, n22611, n22610, n22609, 
        n22608, n22607, n22606, n22605, n22604, n22603, n22602, 
        n22601, n22600, n22599, n22598, n22597, n21921, n22596, 
        n22595, n22594, n22593, n22592, n22591, n21942, n22590, 
        n22589, n22588, n22587, n22586, n22585, n22584, n22583, 
        n22582, n22581, n22580, n22579, n22578, n22577, n22576, 
        n22575, n22574, n22573, n22572;
    wire [31:0]n133;
    
    wire n22571, n22570, n22569, n22568, n21941, n22567, n22566, 
        n21940, n22565, n22564, n22563, n22562, n22561, n22560, 
        n22559, n21939, n22558, n50_adj_4369, n22557, n22556, n22555, 
        n26778, n22554, n22553, n21938, n22552, n22551, n22550, 
        n22549, n22548, n22547, n22546, n22545, n22544, n22543, 
        n22542, n22541, n22540, n22539, n22538, n22537, n838, 
        n807, n60, n23695, n5, n22536, n608, n708, n19068, n739, 
        n12135, n26736, n22535, n25_adj_4372, n27_adj_4373, n29_adj_4374, 
        n26_adj_4375, n16, n21_adj_4376, n28_adj_4377, n30_adj_4378, 
        n23_adj_4379, n17_adj_4380, n22_adj_4381, n24_adj_4382, n44_adj_4383, 
        n30571, n28388, n2225, n30271, n22534, n22533, n22532, 
        n22531, n22530, n22529, n22528, n22527, n30457, n30460, 
        n22526, n22525, n22524, n22523, n22522, n30403, n28514, 
        n30397, n28517, n30385, n30388, n30367, n29897, n22521, 
        n21937, n22520, n22519, n30355, n30358, n22518, n22517, 
        n22516, n22515, n22514, n22513, n22512, n22511, n22510, 
        n22509, n22508, n22507, n22506, n22505, n22504, n26774, 
        n9_adj_4386, n7_adj_4387, n8_adj_4388, n26072, n22503, n22502, 
        n28_adj_4389, n32_adj_4390, n30_adj_4391, n31_adj_4392, n29_adj_4393, 
        n2324, n30270, n26073, n2302, n2292, n22_adj_4395, n2299, 
        n2309, n30_adj_4396, n2294, n2306, n2297, n34_adj_4397, 
        n2301, n2307, n2291, n2305, n32_adj_4398, n22501, n2298, 
        n2295, n2304, n2300, n33_adj_4399, n4_adj_4400, n2308, n2296, 
        n2303, n2293, n31_adj_4401;
    wire [3:0]state_3__N_248;
    
    wire n22500, n22499, n22498, n2423, n30269, n22497, n22496, 
        n21936, n29213, n2403, n2409, n27_adj_4402, n2390, n2391, 
        n2397, n2394, n33_adj_4403, n2392, n2405, n2400, n2398, 
        n32_adj_4404, n2396, n2402, n2408, n2399, n31_adj_4405, 
        n2393, n2406, n2395, n2407, n35_adj_4406, n2404, n2401, 
        n37_adj_4407, n22495, n30268, n22494, n22493, n22492, n22491, 
        n22490, n22489, n22488, n22487, n22486, n22485, n22484, 
        n28318, n22483, n22482, n22481, n22480, n22479, n22478, 
        n22477, n22476, n22475, n22474, n28326, n21935, n26854, 
        n21934, n22473, n22472, n22471, n22470, n22469, n22468, 
        n21933, n22467, n21914, n21920, n22466, n22465, n22464, 
        n22463, n22462, n21932, n22461, n22168, n22460, n22459, 
        n22458, n22457, n22456, n22455, n22454, n22453, n22452, 
        n22167, n22451, n22450, n22449, n22448, n22447, n22446, 
        n22445, n22444, n22443, n18, n22442, n28_adj_4410, n22441, 
        n22440, n22439, n22438, n22437, n22166, n26_adj_4411, n1994, 
        n27_adj_4412, n22165, n1928, n30281, n25_adj_4413, n22416, 
        n22415, n22414, n22413, n22164, n22412, n22373, n22372, 
        n22371, n22370, n22369, n22368, n22367, n22366, n22365, 
        n22364, n22363, n22362, n22361, n22360, n22359, n22358, 
        n22357, n22356, n22355, n22354, n22353, n22352, n22351, 
        n22350, n22349, n22348, n22347, n22346, n22345, n22344, 
        n22343, n22342, n22341, n22340, n1895, n1902, n1899, n1897, 
        n26_adj_4419, n1907, n1909, n19_adj_4420, n1908, n1900, 
        n16_adj_4421, n22339, n22338, n22337, n21931, n22336, n22335, 
        n21930, n22334, n22333, n1904, n1901, n1906, n1898, n24_adj_4422, 
        n22332, n1905, n1903, n28_adj_4423, n22331, n22330, n1896, 
        n1829, n30280, n1301, n22329, n1302, n22328, n1806, n1803, 
        n1798, n1805, n24_adj_4428, n1808, n1804, n1802, n1807, 
        n22_adj_4429, n1800, n1799, n1797, n1801, n23_adj_4430, 
        n1796, n1809, n21_adj_4431, n1730, n30279, n1699, n1709, 
        n17_adj_4434, n1698, n1707, n1703, n1705, n21_adj_4435, 
        n1704, n1701, n1708, n20_adj_4436, n1702, n1697, n24_adj_4437, 
        n1700, n1706, n1631, n30278, n29508, n29331, n26884, n26888, 
        n1303, n22327, \neo_pixel_transmitter.done_N_462 , n1304, n22326, 
        n1305, n22325, n1306, n22324, n1307, n22323, n1308, n30274, 
        n22322, n1309, n1400, n1334, n22321, n1401, n22320, n1402, 
        n22319, n21919, n1403, n22318, n1404, n22317, n1405, n22316, 
        n21929, n1406, n22315, n22163, n1407, n22314, n22162, 
        n22161, n22160, n22159, n22158, n1408, n30275, n22313, 
        n1409, n1499, n1433, n22312, n22157, n7_adj_4445, n14750, 
        n1500, n22311, n1501, n22310, n1502, n22309, n1503, n22308, 
        n1504, n22307, n1505, n22306, n1506, n22305, n1507, n22304, 
        n1508, n30276, n22303, n1509, n22156, n1598, n1532, n22302, 
        n1599, n22301, n1600, n22300, n1601, n22299, n1602, n22298, 
        n1603, n22297, n1604, n22296, n1605, n22295, n1606, n22294, 
        n22155, n1607, n22293, n22154, n1608, n30277, n22292, 
        n1609, n22291, n22290, n22289, n21918, n22288, n22287, 
        n22286, n22285, n22284, n22283, n20_adj_4449, n13_adj_4450, 
        n18_adj_4451, n22_adj_4452, n18_adj_4453, n20_adj_4454, n22282, 
        n15_adj_4455, n22153, n22281, n21928, n22280, n22279, n22278, 
        n22277, n22276, n22275, n22274, n22273, n22152, n22272, 
        n22271, n10_adj_4456, n22151, n22270;
    wire [4:0]color_bit_N_442;
    
    wire n29281, n22269, n22268, n22267, n19303, n22266, n22265, 
        n22264, n16_adj_4457, n22263, n17_adj_4458, n22150, n22149, 
        n22262, n22261, n22260, n22259, n10_adj_4459, n22148, n12_adj_4460, 
        n22258, n16_adj_4461, n22257, n22256, n22147, n22146, n22255, 
        n22254, n21927, n22253, n21926, n22252, n22251, n22250, 
        n22249, n22248, n22247, n22246, n22145, n22144, n22245, 
        n22244, n22143, n22243, n22142, n22242, n22241, n22240, 
        n22239, n22238, n22141;
    
    SB_CARRY mod_5_add_1406_17 (.CI(n22065), .I0(n1995), .I1(n2027), .CO(n22066));
    SB_LUT4 i25196_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30260));
    defparam i25196_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n27007), .D(\neo_pixel_transmitter.done_N_456 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i17055_4_lut (.I0(n26858), .I1(n28), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n64));   // verilog/neopixel.v(27[7:11])
    defparam i17055_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(start), .I2(\one_wire_N_399[11] ), 
            .I3(n64), .O(n1554));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n22064), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_4 (.CI(n22139), .I0(timer[2]), .I1(n1[2]), .CO(n22140));
    SB_LUT4 sub_14_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n22138), .O(one_wire_N_399[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_16 (.CI(n22064), .I0(n1996), .I1(n2027), .CO(n22065));
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4305));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15473_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n19275));
    defparam i15473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n19275), 
            .O(n36));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n2700), .I1(n38), .I2(n28_adj_4305), .I3(n2705), 
            .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n2687), .I1(n36), .I2(n2703), .I3(n2695), 
            .O(n41));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25201_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30265));
    defparam i25201_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n14635), 
            .D(n255[5]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1455 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34));
    defparam i13_4_lut_adj_1455.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), .I3(GND_net), 
            .O(n22));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1456 (.I0(n2490), .I1(n34), .I2(n24), .I3(n2494), 
            .O(n38_adj_4306));
    defparam i17_4_lut_adj_1456.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1457 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4307));
    defparam i15_4_lut_adj_1457.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1458 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22), 
            .O(n37));
    defparam i16_4_lut_adj_1458.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37), .I2(n36_adj_4307), .I3(n38_adj_4306), 
            .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25203_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30267));
    defparam i25203_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1459 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4308));
    defparam i16_4_lut_adj_1459.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_3 (.CI(n22138), .I0(timer[1]), .I1(n1[1]), .CO(n22139));
    SB_LUT4 i14_4_lut_adj_1460 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4309));
    defparam i14_4_lut_adj_1460.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1461 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4310));
    defparam i15_4_lut_adj_1461.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1462 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4311));
    defparam i13_4_lut_adj_1462.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4312));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n22063), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1463 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4313));
    defparam i18_4_lut_adj_1463.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1464 (.I0(n37_adj_4311), .I1(n39_adj_4310), .I2(n38_adj_4309), 
            .I3(n40_adj_4308), .O(n46));
    defparam i22_4_lut_adj_1464.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4314));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4314), .I1(n46), .I2(n42_adj_4313), 
            .I3(n34_adj_4312), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25200_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30264));
    defparam i25200_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4315));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1465 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4316));
    defparam i16_4_lut_adj_1465.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4317));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1466 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43));
    defparam i18_4_lut_adj_1466.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1467 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4318));
    defparam i15_4_lut_adj_1467.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n41_adj_4316), .I1(n33_adj_4315), .I2(n2889), 
            .I3(n2901), .O(n46_adj_4319));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1468 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4320));
    defparam i14_4_lut_adj_1468.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1469 (.I0(n43), .I1(n2904), .I2(n38_adj_4317), 
            .I3(n2893), .O(n47));
    defparam i22_4_lut_adj_1469.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_4320), .I2(n46_adj_4319), 
            .I3(n40_adj_4318), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25199_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30263));
    defparam i25199_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15536_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n19339));
    defparam i15536_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1470 (.I0(n35_adj_4321), .I1(n11), .I2(n29), 
            .I3(n51), .O(n48));
    defparam i20_4_lut_adj_1470.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1471 (.I0(n37_adj_4322), .I1(n23), .I2(n53), 
            .I3(n39_adj_4323), .O(n46_adj_4324));
    defparam i18_4_lut_adj_1471.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1472 (.I0(n27), .I1(n57), .I2(n63), .I3(n43_adj_4325), 
            .O(n47_adj_4326));
    defparam i19_4_lut_adj_1472.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1473 (.I0(n25), .I1(n33_adj_4327), .I2(n47_adj_4328), 
            .I3(n61), .O(n45));
    defparam i17_4_lut_adj_1473.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1474 (.I0(n59), .I1(n17), .I2(n15), .I3(n55), 
            .O(n44));
    defparam i16_4_lut_adj_1474.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1475 (.I0(n31_adj_4329), .I1(n41_adj_4330), .I2(n49), 
            .I3(n19339), .O(n43_adj_4331));
    defparam i15_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_adj_4326), .I2(n46_adj_4324), 
            .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1476 (.I0(n45_adj_4332), .I1(n13), .I2(n19), 
            .I3(n21), .O(n49_adj_4333));
    defparam i21_4_lut_adj_1476.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4333), .I1(n54), .I2(n43_adj_4331), 
            .I3(n44), .O(n23391));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[3]), .I1(n23391), .I2(GND_net), .I3(GND_net), 
            .O(n23679));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_1477 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4334));
    defparam i14_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1478 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4335));
    defparam i18_4_lut_adj_1478.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1479 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4336));
    defparam i16_4_lut_adj_1479.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1480 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4337));
    defparam i17_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1481 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4338));
    defparam i15_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_4339));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4334), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4340));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut_adj_1482 (.I0(n41_adj_4338), .I1(n43_adj_4337), .I2(n42_adj_4336), 
            .I3(n44_adj_4335), .O(n50));
    defparam i24_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4341));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_4341), .I1(n50), .I2(n46_adj_4340), 
            .I3(n38_adj_4339), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25198_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30262));
    defparam i25198_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n23164), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n23163), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n23163), .I0(n2094), .I1(n2126), .CO(n23164));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n23162), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n23162), .I0(n2095), .I1(n2126), .CO(n23163));
    SB_LUT4 sub_14_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(one_wire_N_399[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n23161), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n23161), .I0(n2096), .I1(n2126), .CO(n23162));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n23160), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n23160), .I0(n2097), .I1(n2126), .CO(n23161));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n23159), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n23159), .I0(n2098), .I1(n2126), .CO(n23160));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n23158), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n23158), .I0(n2099), .I1(n2126), .CO(n23159));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n23157), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n23157), .I0(n2100), .I1(n2126), .CO(n23158));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n23156), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n23156), .I0(n2101), .I1(n2126), .CO(n23157));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n23155), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n23155), .I0(n2102), .I1(n2126), .CO(n23156));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n23154), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n23154), .I0(n2103), .I1(n2126), .CO(n23155));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n23153), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n22138));
    SB_CARRY mod_5_add_1473_8 (.CI(n23153), .I0(n2104), .I1(n2126), .CO(n23154));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n23152), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n23152), .I0(n2105), .I1(n2126), .CO(n23153));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n23151), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n23151), .I0(n2106), .I1(n2126), .CO(n23152));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n23150), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n23150), .I0(n2107), .I1(n2126), .CO(n23151));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n23149), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n23149), .I0(n2108), .I1(n2126), .CO(n23150));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n30260), 
            .I3(n23148), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n23148), .I0(n2109), .I1(n30260), .CO(n23149));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n30260), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n30260), 
            .CO(n23148));
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n14635), 
            .D(n255[4]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n14635), 
            .D(n255[3]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n14635), 
            .D(n255[2]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n14635), 
            .D(n255[1]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1406_15 (.CI(n22063), .I0(n1997), .I1(n2027), .CO(n22064));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n22062), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_3_lut_adj_1483 (.I0(n2096), .I1(n2103), .I2(n2097), .I3(GND_net), 
            .O(n26));
    defparam i9_3_lut_adj_1483.LUT_INIT = 16'hfefe;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n21916), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1484 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42_adj_4342));
    defparam i15_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1485 (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46_adj_4343));
    defparam i19_4_lut_adj_1485.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1486 (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44_adj_4344));
    defparam i17_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1487 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45_adj_4345));
    defparam i18_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1488 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43_adj_4346));
    defparam i16_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1489 (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), 
            .I3(GND_net), .O(n40_adj_4347));
    defparam i13_3_lut_adj_1489.LUT_INIT = 16'hecec;
    SB_LUT4 i21_4_lut_adj_1490 (.I0(n3107), .I1(n42_adj_4342), .I2(n3087), 
            .I3(n3086), .O(n48_adj_4348));
    defparam i21_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1491 (.I0(n43_adj_4346), .I1(n45_adj_4345), .I2(n44_adj_4344), 
            .I3(n46_adj_4343), .O(n52));
    defparam i25_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut_adj_1492 (.I0(n3095), .I1(n3084), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4349));
    defparam i12_2_lut_adj_1492.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut_adj_1493 (.I0(n39_adj_4349), .I1(n52), .I2(n48_adj_4348), 
            .I3(n40_adj_4347), .O(n3116));
    defparam i26_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1494 (.I0(bit_ctr[14]), .I1(n26), .I2(n2100), 
            .I3(n2109), .O(n30));
    defparam i13_4_lut_adj_1494.LUT_INIT = 16'hfefc;
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n21924), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25195_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30259));
    defparam i25195_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1495 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4350));
    defparam i14_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n25_adj_4351));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4352));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1496 (.I0(n25_adj_4351), .I1(n36_adj_4350), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4353));
    defparam i18_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1497 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4354));
    defparam i16_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4352), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4355));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1498 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4356));
    defparam i15_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1499 (.I0(n37_adj_4356), .I1(n39_adj_4355), .I2(n38_adj_4354), 
            .I3(n40_adj_4353), .O(n2621));
    defparam i21_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 i25202_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30266));
    defparam i25202_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_14 (.CI(n22062), .I0(n1998), .I1(n2027), .CO(n22063));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n22061), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n22061), .I0(n1999), .I1(n2027), .CO(n22062));
    SB_LUT4 i11_4_lut (.I0(n2102), .I1(n2099), .I2(n2094), .I3(n2105), 
            .O(n28_adj_4357));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n22060), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut_adj_1500 (.I0(n2095), .I1(n2108), .I2(n2098), .I3(n2093), 
            .O(n29_adj_4358));
    defparam i12_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_12 (.CI(n22060), .I0(n2000), .I1(n2027), .CO(n22061));
    SB_LUT4 i10_4_lut (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4359));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1501 (.I0(n27_adj_4359), .I1(n29_adj_4358), .I2(n28_adj_4357), 
            .I3(n30), .O(n2126));
    defparam i16_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n22059), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1502 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9));
    defparam i1_3_lut_adj_1502.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut (.I0(n9), .I1(n14), .I2(n1202), .I3(n1208), .O(n1235));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_5 (.CI(n21916), .I0(bit_ctr[3]), .I1(GND_net), .CO(n21917));
    SB_CARRY mod_5_add_1406_11 (.CI(n22059), .I0(n2001), .I1(n2027), .CO(n22060));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n22058), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25209_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30273));
    defparam i25209_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_10 (.CI(n22058), .I0(n2002), .I1(n2027), .CO(n22059));
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n14635), 
            .D(n255[15]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_13 (.CI(n21924), .I0(bit_ctr[11]), .I1(GND_net), .CO(n21925));
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n14635), 
            .D(n255[14]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n22057), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n22057), .I0(n2003), .I1(n2027), .CO(n22058));
    SB_LUT4 i15489_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n19291));
    defparam i15489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n19291), .I3(n1108), 
            .O(n12_c));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1503 (.I0(n1107), .I1(n12_c), .I2(n1106), .I3(n1104), 
            .O(n1136));
    defparam i6_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n14635), 
            .D(n255[8]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n22056), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n22056), .I0(n2004), .I1(n2027), .CO(n22057));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n22055), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n22055), .I0(n2005), .I1(n2027), .CO(n22056));
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n14635), 
            .D(n255[7]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_4_lut_adj_1504 (.I0(one_wire_N_399[4]), .I1(n110), .I2(one_wire_N_399[3]), 
            .I3(one_wire_N_399[2]), .O(n28));   // verilog/neopixel.v(6[16:24])
    defparam i1_4_lut_adj_1504.LUT_INIT = 16'heccc;
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n22054), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n22054), .I0(n2006), .I1(n2027), .CO(n22055));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n22053), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n22053), .I0(n2007), .I1(n2027), .CO(n22054));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n22052), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n22052), .I0(n2008), .I1(n2027), .CO(n22053));
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n14635), 
            .D(n255[6]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i25208_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30272));
    defparam i25208_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25192_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i25192_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i25190_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i25190_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n12133), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_3_lut_adj_1505 (.I0(n26828), .I1(n906), .I2(n14692), .I3(GND_net), 
            .O(n8));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut_adj_1505.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut (.I0(n905), .I1(n8), .I2(bit_ctr[26]), .I3(n12133), 
            .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h0444;
    SB_LUT4 i23321_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n28384));
    defparam i23321_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n30259), 
            .I3(n22051), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_4_lut (.I0(n2), .I1(n6), .I2(n1005), .I3(n28384), .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n21923), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25073_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_c));   // verilog/neopixel.v(22[26:36])
    defparam i25073_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_1406_3 (.CI(n22051), .I0(n2009), .I1(n30259), .CO(n22052));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n30259), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n30259), 
            .CO(n22051));
    SB_CARRY add_21_12 (.CI(n21923), .I0(bit_ctr[10]), .I1(GND_net), .CO(n21924));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n21922), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n21944), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n22661), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n22660), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n22660), .I0(n3084), .I1(n3116), .CO(n22661));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n22659), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n22659), .I0(n3085), .I1(n3116), .CO(n22660));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n22658), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n22658), .I0(n3086), .I1(n3116), .CO(n22659));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n22657), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n22657), .I0(n3087), .I1(n3116), .CO(n22658));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n22656), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n22656), .I0(n3088), .I1(n3116), .CO(n22657));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n22655), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n22655), .I0(n3089), .I1(n3116), .CO(n22656));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n22654), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n22654), .I0(n3090), .I1(n3116), .CO(n22655));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n22653), .O(n47_adj_4328)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n22653), .I0(n3091), .I1(n3116), .CO(n22654));
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n21915), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut_adj_1506 (.I0(bit_ctr[23]), .I1(bit_ctr[16]), .I2(bit_ctr[20]), 
            .I3(bit_ctr[7]), .O(n46_adj_4360));
    defparam i19_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1507 (.I0(bit_ctr[14]), .I1(bit_ctr[9]), .I2(bit_ctr[25]), 
            .I3(bit_ctr[10]), .O(n44_adj_4361));
    defparam i17_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1508 (.I0(bit_ctr[27]), .I1(bit_ctr[12]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[29]), .O(n45_adj_4362));
    defparam i18_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1509 (.I0(bit_ctr[6]), .I1(bit_ctr[31]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[21]), .O(n43_adj_4363));
    defparam i16_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1510 (.I0(bit_ctr[17]), .I1(bit_ctr[28]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[5]), .O(n42_adj_4364));
    defparam i15_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_3_lut (.I0(bit_ctr[26]), .I1(bit_ctr[13]), .I2(bit_ctr[22]), 
            .I3(GND_net), .O(n41_adj_4365));
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i25_4_lut_adj_1511 (.I0(n43_adj_4363), .I1(n45_adj_4362), .I2(n44_adj_4361), 
            .I3(n46_adj_4360), .O(n52_adj_4366));
    defparam i25_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1512 (.I0(bit_ctr[30]), .I1(bit_ctr[18]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[8]), .O(n47_adj_4367));
    defparam i20_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1513 (.I0(n47_adj_4367), .I1(n52_adj_4366), .I2(n41_adj_4365), 
            .I3(n42_adj_4364), .O(n24472));
    defparam i26_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1514 (.I0(one_wire_N_399[3]), .I1(one_wire_N_399[1]), 
            .I2(one_wire_N_399[0]), .I3(one_wire_N_399[2]), .O(n73));   // verilog/neopixel.v(53[15:25])
    defparam i1_4_lut_adj_1514.LUT_INIT = 16'haaa8;
    SB_LUT4 i3_4_lut_adj_1515 (.I0(one_wire_N_399[10]), .I1(n73), .I2(one_wire_N_399[4]), 
            .I3(n7), .O(n26858));
    defparam i3_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\one_wire_N_399[11] ), .I1(n26858), .I2(GND_net), 
            .I3(GND_net), .O(n86));
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1517 (.I0(\neo_pixel_transmitter.done ), .I1(n20817), 
            .I2(n83), .I3(\state[0] ), .O(n20822));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut_adj_1517.LUT_INIT = 16'h0a88;
    SB_LUT4 i17047_4_lut (.I0(n29305), .I1(n20817), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n34_adj_4368));   // verilog/neopixel.v(16[20:25])
    defparam i17047_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i10940_4_lut (.I0(n14635), .I1(\neo_pixel_transmitter.done ), 
            .I2(n86), .I3(n34_adj_4368), .O(n14745));   // verilog/neopixel.v(35[12] 117[6])
    defparam i10940_4_lut.LUT_INIT = 16'haa2a;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n22652), .O(n45_adj_4332)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n22652), .I0(n3092), .I1(n3116), .CO(n22653));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n22651), .O(n43_adj_4325)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n22651), .I0(n3093), .I1(n3116), .CO(n22652));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n22650), .O(n41_adj_4330)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n22650), .I0(n3094), .I1(n3116), .CO(n22651));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n22649), .O(n39_adj_4323)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n22649), .I0(n3095), .I1(n3116), .CO(n22650));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n22648), .O(n37_adj_4322)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n22648), .I0(n3096), .I1(n3116), .CO(n22649));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n22647), .O(n35_adj_4321)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n22647), .I0(n3097), .I1(n3116), .CO(n22648));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n22646), .O(n33_adj_4327)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n22646), .I0(n3098), .I1(n3116), .CO(n22647));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n22645), .O(n31_adj_4329)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n22645), .I0(n3099), .I1(n3116), .CO(n22646));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n22644), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n22644), .I0(n3100), .I1(n3116), .CO(n22645));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n22643), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n22643), .I0(n3101), .I1(n3116), .CO(n22644));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n22642), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n22642), .I0(n3102), .I1(n3116), .CO(n22643));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n22641), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n22641), .I0(n3103), .I1(n3116), .CO(n22642));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n22640), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n22640), .I0(n3104), .I1(n3116), .CO(n22641));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n22639), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n22639), .I0(n3105), .I1(n3116), .CO(n22640));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n22638), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n22638), .I0(n3106), .I1(n3116), .CO(n22639));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n22637), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n22637), .I0(n3107), .I1(n3116), .CO(n22638));
    SB_CARRY add_21_11 (.CI(n21922), .I0(bit_ctr[9]), .I1(GND_net), .CO(n21923));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n22636), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n22636), .I0(n3108), .I1(n3116), .CO(n22637));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n30262), 
            .I3(n22635), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n14635), 
            .D(n255[0]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2143_3 (.CI(n22635), .I0(n3109), .I1(n30262), .CO(n22636));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n30262), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n30262), 
            .CO(n22635));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n22634), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n22633), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n22633), .I0(n2985), .I1(n3017), .CO(n22634));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n22632), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n22632), .I0(n2986), .I1(n3017), .CO(n22633));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n22631), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n22631), .I0(n2987), .I1(n3017), .CO(n22632));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n22630), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n22630), .I0(n2988), .I1(n3017), .CO(n22631));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n22629), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n22629), .I0(n2989), .I1(n3017), .CO(n22630));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n22628), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17038_4_lut (.I0(n20822), .I1(n29304), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n14635));   // verilog/neopixel.v(16[20:25])
    defparam i17038_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n21943), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_22 (.CI(n22628), .I0(n2990), .I1(n3017), .CO(n22629));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n22627), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n22627), .I0(n2991), .I1(n3017), .CO(n22628));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n22626), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n22626), .I0(n2992), .I1(n3017), .CO(n22627));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n22625), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n22625), .I0(n2993), .I1(n3017), .CO(n22626));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n22624), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n22624), .I0(n2994), .I1(n3017), .CO(n22625));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n22623), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n22623), .I0(n2995), .I1(n3017), .CO(n22624));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n22622), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n22622), .I0(n2996), .I1(n3017), .CO(n22623));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n22621), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n22621), .I0(n2997), .I1(n3017), .CO(n22622));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n22620), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n22620), .I0(n2998), .I1(n3017), .CO(n22621));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n22619), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n22619), .I0(n2999), .I1(n3017), .CO(n22620));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n22618), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n22618), .I0(n3000), .I1(n3017), .CO(n22619));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n22617), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n22617), .I0(n3001), .I1(n3017), .CO(n22618));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n22616), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n22616), .I0(n3002), .I1(n3017), .CO(n22617));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n22615), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n22615), .I0(n3003), .I1(n3017), .CO(n22616));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n22614), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n22614), .I0(n3004), .I1(n3017), .CO(n22615));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n22613), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n22613), .I0(n3005), .I1(n3017), .CO(n22614));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n22612), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n22612), .I0(n3006), .I1(n3017), .CO(n22613));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n22611), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n22611), .I0(n3007), .I1(n3017), .CO(n22612));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n22610), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n22610), .I0(n3008), .I1(n3017), .CO(n22611));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n30263), 
            .I3(n22609), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n22609), .I0(n3009), .I1(n30263), .CO(n22610));
    SB_CARRY add_21_32 (.CI(n21943), .I0(bit_ctr[30]), .I1(GND_net), .CO(n21944));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n30263), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_4 (.CI(n21915), .I0(bit_ctr[2]), .I1(GND_net), .CO(n21916));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n30263), 
            .CO(n22609));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n22608), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n22607), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n22607), .I0(n2886), .I1(n2918), .CO(n22608));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n22606), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n22606), .I0(n2887), .I1(n2918), .CO(n22607));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n22605), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n22605), .I0(n2888), .I1(n2918), .CO(n22606));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n22604), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n22604), .I0(n2889), .I1(n2918), .CO(n22605));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n22603), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n22603), .I0(n2890), .I1(n2918), .CO(n22604));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n22602), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n22602), .I0(n2891), .I1(n2918), .CO(n22603));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n22601), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n22601), .I0(n2892), .I1(n2918), .CO(n22602));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n22600), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n22600), .I0(n2893), .I1(n2918), .CO(n22601));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n22599), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n22599), .I0(n2894), .I1(n2918), .CO(n22600));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n22598), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n22598), .I0(n2895), .I1(n2918), .CO(n22599));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n22597), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n22597), .I0(n2896), .I1(n2918), .CO(n22598));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n21921), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n22596), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n22596), .I0(n2897), .I1(n2918), .CO(n22597));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n22595), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n22595), .I0(n2898), .I1(n2918), .CO(n22596));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n22594), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n22594), .I0(n2899), .I1(n2918), .CO(n22595));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n22593), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n22593), .I0(n2900), .I1(n2918), .CO(n22594));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n22592), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n22592), .I0(n2901), .I1(n2918), .CO(n22593));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n22591), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n22591), .I0(n2902), .I1(n2918), .CO(n22592));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n21942), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n22590), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n22590), .I0(n2903), .I1(n2918), .CO(n22591));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n22589), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n22589), .I0(n2904), .I1(n2918), .CO(n22590));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n22588), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n22588), .I0(n2905), .I1(n2918), .CO(n22589));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n22587), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n22587), .I0(n2906), .I1(n2918), .CO(n22588));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n22586), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n22586), .I0(n2907), .I1(n2918), .CO(n22587));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n22585), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n22585), .I0(n2908), .I1(n2918), .CO(n22586));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n30264), 
            .I3(n22584), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n22584), .I0(n2909), .I1(n30264), .CO(n22585));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n30264), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n30264), 
            .CO(n22584));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n22583), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n22582), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n22582), .I0(n2787), .I1(n2819), .CO(n22583));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n22581), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n22581), .I0(n2788), .I1(n2819), .CO(n22582));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n22580), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n22580), .I0(n2789), .I1(n2819), .CO(n22581));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n22579), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n22579), .I0(n2790), .I1(n2819), .CO(n22580));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n22578), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n22578), .I0(n2791), .I1(n2819), .CO(n22579));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n22577), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n22577), .I0(n2792), .I1(n2819), .CO(n22578));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n22576), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n22576), .I0(n2793), .I1(n2819), .CO(n22577));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n22575), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n22575), .I0(n2794), .I1(n2819), .CO(n22576));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n22574), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n22574), .I0(n2795), .I1(n2819), .CO(n22575));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n22573), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n22573), .I0(n2796), .I1(n2819), .CO(n22574));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n22572), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1122__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1942_15 (.CI(n22572), .I0(n2797), .I1(n2819), .CO(n22573));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n22571), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n22571), .I0(n2798), .I1(n2819), .CO(n22572));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n22570), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n22570), .I0(n2799), .I1(n2819), .CO(n22571));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n22569), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n22569), .I0(n2800), .I1(n2819), .CO(n22570));
    SB_CARRY add_21_31 (.CI(n21942), .I0(bit_ctr[29]), .I1(GND_net), .CO(n21943));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n22568), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n21941), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_11 (.CI(n22568), .I0(n2801), .I1(n2819), .CO(n22569));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n22567), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_30 (.CI(n21941), .I0(bit_ctr[28]), .I1(GND_net), .CO(n21942));
    SB_CARRY mod_5_add_1942_10 (.CI(n22567), .I0(n2802), .I1(n2819), .CO(n22568));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n22566), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n22566), .I0(n2803), .I1(n2819), .CO(n22567));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n21940), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n22565), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n22565), .I0(n2804), .I1(n2819), .CO(n22566));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n22564), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n22564), .I0(n2805), .I1(n2819), .CO(n22565));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n22563), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n22563), .I0(n2806), .I1(n2819), .CO(n22564));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n22562), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n22562), .I0(n2807), .I1(n2819), .CO(n22563));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n22561), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n22561), .I0(n2808), .I1(n2819), .CO(n22562));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n30265), 
            .I3(n22560), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n22560), .I0(n2809), .I1(n30265), .CO(n22561));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n30265), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n30265), 
            .CO(n22560));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n22559), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_29 (.CI(n21940), .I0(bit_ctr[27]), .I1(GND_net), .CO(n21941));
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n21939), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n21939), .I0(bit_ctr[26]), .I1(GND_net), .CO(n21940));
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n22558), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n22558), .I0(n2688), .I1(n2720), .CO(n22559));
    SB_LUT4 i24528_3_lut_4_lut (.I0(n50_adj_4369), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(start), .O(n29233));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24528_3_lut_4_lut.LUT_INIT = 16'hff02;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n22557), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n22557), .I0(n2689), .I1(n2720), .CO(n22558));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n22556), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n22556), .I0(n2690), .I1(n2720), .CO(n22557));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n22555), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n22555), .I0(n2691), .I1(n2720), .CO(n22556));
    SB_LUT4 i21724_2_lut_3_lut (.I0(n50_adj_4369), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(GND_net), .O(n26778));   // verilog/neopixel.v(35[12] 117[6])
    defparam i21724_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n14869));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n22554), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n22554), .I0(n2692), .I1(n2720), .CO(n22555));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n22553), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n21938), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_19 (.CI(n22553), .I0(n2693), .I1(n2720), .CO(n22554));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n22552), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n22552), .I0(n2694), .I1(n2720), .CO(n22553));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n22551), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n22551), .I0(n2695), .I1(n2720), .CO(n22552));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n22550), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n22550), .I0(n2696), .I1(n2720), .CO(n22551));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n22549), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n22549), .I0(n2697), .I1(n2720), .CO(n22550));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n22548), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n22548), .I0(n2698), .I1(n2720), .CO(n22549));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n22547), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n22547), .I0(n2699), .I1(n2720), .CO(n22548));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n22546), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n22546), .I0(n2700), .I1(n2720), .CO(n22547));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n22545), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n22545), .I0(n2701), .I1(n2720), .CO(n22546));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n22544), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n22544), .I0(n2702), .I1(n2720), .CO(n22545));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n22543), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n22543), .I0(n2703), .I1(n2720), .CO(n22544));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n22542), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n22542), .I0(n2704), .I1(n2720), .CO(n22543));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n22541), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n22541), .I0(n2705), .I1(n2720), .CO(n22542));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n22540), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n22540), .I0(n2706), .I1(n2720), .CO(n22541));
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n14868));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n22539), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1518 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_adj_1518.LUT_INIT = 16'h4444;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n14635), 
            .D(n255[31]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1875_5 (.CI(n22539), .I0(n2707), .I1(n2720), .CO(n22540));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n22538), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n22538), .I0(n2708), .I1(n2720), .CO(n22539));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n30266), 
            .I3(n22537), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n12133));
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'h9999;
    SB_CARRY mod_5_add_1875_3 (.CI(n22537), .I0(n2709), .I1(n30266), .CO(n22538));
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n30266), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n30266), 
            .CO(n22537));
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i1_2_lut_adj_1520 (.I0(bit_ctr[28]), .I1(n23695), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_adj_1520.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n22536), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15443_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i15443_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n608), .I2(n5), .I3(n19068), .O(n739));
    defparam i2_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n12135));
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i24611_3_lut (.I0(n23695), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n26736));
    defparam i24611_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n12135), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n26736), .O(n26828));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n5), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n22535), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n22535), .I0(n2589), .I1(n2621), .CO(n22536));
    SB_LUT4 i6_4_lut_adj_1522 (.I0(n25_adj_4372), .I1(n27_adj_4373), .I2(n29_adj_4374), 
            .I3(n26_adj_4375), .O(n16));
    defparam i6_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1523 (.I0(n21_adj_4376), .I1(n28_adj_4377), .I2(n30_adj_4378), 
            .I3(n23_adj_4379), .O(n17_adj_4380));
    defparam i7_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n17_adj_4380), .I1(n22_adj_4381), .I2(n16), 
            .I3(n24_adj_4382), .O(n44_adj_4383));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i132_4_lut (.I0(\one_wire_N_399[11] ), .I1(n44_adj_4383), .I2(one_wire_N_399[10]), 
            .I3(one_wire_N_399[9]), .O(n50_adj_4369));   // verilog/neopixel.v(6[16:24])
    defparam i132_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n30571));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30571_bdd_4_lut (.I0(n30571), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n28388));
    defparam n30571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i25207_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30271));
    defparam i25207_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n22534), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n22534), .I0(n2590), .I1(n2621), .CO(n22535));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n22533), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n22533), .I0(n2591), .I1(n2621), .CO(n22534));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n22532), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n22532), .I0(n2592), .I1(n2621), .CO(n22533));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n22531), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n22531), .I0(n2593), .I1(n2621), .CO(n22532));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n22530), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n22530), .I0(n2594), .I1(n2621), .CO(n22531));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n22529), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n22529), .I0(n2595), .I1(n2621), .CO(n22530));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n22528), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n22528), .I0(n2596), .I1(n2621), .CO(n22529));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n22527), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n22527), .I0(n2597), .I1(n2621), .CO(n22528));
    SB_LUT4 bit_ctr_0__bdd_4_lut_25456 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n30457));
    defparam bit_ctr_0__bdd_4_lut_25456.LUT_INIT = 16'he4aa;
    SB_LUT4 n30457_bdd_4_lut (.I0(n30457), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n30460));
    defparam n30457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n22526), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n22526), .I0(n2598), .I1(n2621), .CO(n22527));
    SB_CARRY add_21_27 (.CI(n21938), .I0(bit_ctr[25]), .I1(GND_net), .CO(n21939));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n22525), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n22525), .I0(n2599), .I1(n2621), .CO(n22526));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n22524), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n22524), .I0(n2600), .I1(n2621), .CO(n22525));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n22523), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n22523), .I0(n2601), .I1(n2621), .CO(n22524));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n22522), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n22522), .I0(n2602), .I1(n2621), .CO(n22523));
    SB_LUT4 bit_ctr_0__bdd_4_lut_25361 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n30403));
    defparam bit_ctr_0__bdd_4_lut_25361.LUT_INIT = 16'he4aa;
    SB_LUT4 n30403_bdd_4_lut (.I0(n30403), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n28514));
    defparam n30403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25316 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n30397));
    defparam bit_ctr_0__bdd_4_lut_25316.LUT_INIT = 16'he4aa;
    SB_LUT4 n30397_bdd_4_lut (.I0(n30397), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n28517));
    defparam n30397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25311 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n30385));
    defparam bit_ctr_0__bdd_4_lut_25311.LUT_INIT = 16'he4aa;
    SB_LUT4 n30385_bdd_4_lut (.I0(n30385), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n30388));
    defparam n30385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25301 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n30367));
    defparam bit_ctr_0__bdd_4_lut_25301.LUT_INIT = 16'he4aa;
    SB_LUT4 n30367_bdd_4_lut (.I0(n30367), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n29897));
    defparam n30367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n22521), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n21937), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_26 (.CI(n21937), .I0(bit_ctr[24]), .I1(GND_net), .CO(n21938));
    SB_CARRY mod_5_add_1808_9 (.CI(n22521), .I0(n2603), .I1(n2621), .CO(n22522));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n22520), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n22520), .I0(n2604), .I1(n2621), .CO(n22521));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n22519), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n22519), .I0(n2605), .I1(n2621), .CO(n22520));
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n28514), .I2(n28517), 
            .I3(n23679), .O(n30355));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30355_bdd_4_lut (.I0(n30355), .I1(n29897), .I2(n28388), .I3(n23679), 
            .O(n30358));
    defparam n30355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n14635), 
            .D(n255[13]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n22518), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n22518), .I0(n2606), .I1(n2621), .CO(n22519));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n22517), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n22517), .I0(n2607), .I1(n2621), .CO(n22518));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n22516), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n22516), .I0(n2608), .I1(n2621), .CO(n22517));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n30267), 
            .I3(n22515), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n22515), .I0(n2609), .I1(n30267), .CO(n22516));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n30267), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n30267), 
            .CO(n22515));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n22514), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n22513), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n22513), .I0(n2490), .I1(n2522), .CO(n22514));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n22512), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n22512), .I0(n2491), .I1(n2522), .CO(n22513));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n22511), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n22511), .I0(n2492), .I1(n2522), .CO(n22512));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n22510), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n22510), .I0(n2493), .I1(n2522), .CO(n22511));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n22509), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n22509), .I0(n2494), .I1(n2522), .CO(n22510));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n22508), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n22508), .I0(n2495), .I1(n2522), .CO(n22509));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n22507), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n22507), .I0(n2496), .I1(n2522), .CO(n22508));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n22506), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n14635), 
            .D(n255[30]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n14867));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n14635), 
            .D(n255[29]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_15 (.CI(n22506), .I0(n2497), .I1(n2522), .CO(n22507));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n22505), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_14 (.CI(n22505), .I0(n2498), .I1(n2522), .CO(n22506));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n22504), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i21720_2_lut (.I0(start), .I1(\one_wire_N_399[11] ), .I2(GND_net), 
            .I3(GND_net), .O(n26774));
    defparam i21720_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut (.I0(n9_adj_4386), .I1(n7_adj_4387), .I2(n8_adj_4388), 
            .I3(GND_net), .O(n7));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1524 (.I0(one_wire_N_399[10]), .I1(n7), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/neopixel.v(53[15:25])
    defparam i1_2_lut_adj_1524.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1741_13 (.CI(n22504), .I0(n2499), .I1(n2522), .CO(n22505));
    SB_LUT4 i25063_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n26072));
    defparam i25063_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n22503), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n22503), .I0(n2500), .I1(n2522), .CO(n22504));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n22502), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n14866));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_11 (.CI(n22502), .I0(n2501), .I1(n2522), .CO(n22503));
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1525 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4389));
    defparam i10_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1526 (.I0(n2203), .I1(n28_adj_4389), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4390));
    defparam i14_4_lut_adj_1526.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1527 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4391));
    defparam i12_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1528 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4392));
    defparam i13_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1529 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4393));
    defparam i11_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1530 (.I0(n29_adj_4393), .I1(n31_adj_4392), .I2(n30_adj_4391), 
            .I3(n32_adj_4390), .O(n2225));
    defparam i17_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i25206_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30270));
    defparam i25206_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1531 (.I0(one_wire_N_399[0]), .I1(n26072), .I2(one_wire_N_399[4]), 
            .I3(one_wire_N_399[1]), .O(n26073));
    defparam i1_4_lut_adj_1531.LUT_INIT = 16'hcccd;
    SB_LUT4 i24487_3_lut_4_lut (.I0(\one_wire_N_399[11] ), .I1(n28), .I2(start), 
            .I3(\state[0] ), .O(n29305));   // verilog/neopixel.v(53[15:25])
    defparam i24487_3_lut_4_lut.LUT_INIT = 16'hf0f1;
    SB_LUT4 i3_2_lut_adj_1532 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4395));
    defparam i3_2_lut_adj_1532.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1533 (.I0(bit_ctr[12]), .I1(n22_adj_4395), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4396));
    defparam i11_4_lut_adj_1533.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1534 (.I0(n2294), .I1(n30_adj_4396), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4397));
    defparam i15_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1535 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4398));
    defparam i13_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n22501), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1536 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4399));
    defparam i14_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1537 (.I0(n26072), .I1(one_wire_N_399[4]), .I2(one_wire_N_399[3]), 
            .I3(GND_net), .O(n4_adj_4400));
    defparam i1_3_lut_adj_1537.LUT_INIT = 16'h2b2b;
    SB_LUT4 i12_4_lut_adj_1538 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4401));
    defparam i12_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1539 (.I0(n31_adj_4401), .I1(n33_adj_4399), .I2(n32_adj_4398), 
            .I3(n34_adj_4397), .O(n2324));
    defparam i18_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(\one_wire_N_399[11] ), .I1(n28), .I2(start), 
            .I3(GND_net), .O(n20817));   // verilog/neopixel.v(53[15:25])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i24245_3_lut_4_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n24472), 
            .I3(\state[0] ), .O(n29210));
    defparam i24245_3_lut_4_lut.LUT_INIT = 16'h0700;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n24472), 
            .I3(GND_net), .O(state_3__N_248[1]));
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'hf8f8;
    SB_CARRY mod_5_add_1741_10 (.CI(n22501), .I0(n2502), .I1(n2522), .CO(n22502));
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n14635), 
            .D(n255[28]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n22500), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n22500), .I0(n2503), .I1(n2522), .CO(n22501));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n22499), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n22499), .I0(n2504), .I1(n2522), .CO(n22500));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n22498), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n22498), .I0(n2505), .I1(n2522), .CO(n22499));
    SB_LUT4 i25205_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30269));
    defparam i25205_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n22497), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n22497), .I0(n2506), .I1(n2522), .CO(n22498));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n22496), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n21936), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24531_2_lut_4_lut (.I0(start), .I1(\one_wire_N_399[11] ), .I2(n26858), 
            .I3(\neo_pixel_transmitter.done ), .O(n29213));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24531_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_CARRY mod_5_add_1741_5 (.CI(n22496), .I0(n2507), .I1(n2522), .CO(n22497));
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), .I3(GND_net), 
            .O(n27_adj_4402));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1541 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4403));
    defparam i13_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1542 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4404));
    defparam i12_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1543 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4405));
    defparam i11_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1544 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4406));
    defparam i15_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1545 (.I0(n33_adj_4403), .I1(n27_adj_4402), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4407));
    defparam i17_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1546 (.I0(n37_adj_4407), .I1(n35_adj_4406), .I2(n31_adj_4405), 
            .I3(n32_adj_4404), .O(n2423));
    defparam i19_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n22495), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n22495), .I0(n2508), .I1(n2522), .CO(n22496));
    SB_LUT4 i25204_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30268));
    defparam i25204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n30268), 
            .I3(n22494), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n22494), .I0(n2509), .I1(n30268), .CO(n22495));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n30268), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n30268), 
            .CO(n22494));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n22493), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n22492), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n22492), .I0(n2391), .I1(n2423), .CO(n22493));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n22491), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n22491), .I0(n2392), .I1(n2423), .CO(n22492));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n22490), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n22490), .I0(n2393), .I1(n2423), .CO(n22491));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n22489), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n22489), .I0(n2394), .I1(n2423), .CO(n22490));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n22488), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n22488), .I0(n2395), .I1(n2423), .CO(n22489));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n22487), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n22487), .I0(n2396), .I1(n2423), .CO(n22488));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n22486), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n22486), .I0(n2397), .I1(n2423), .CO(n22487));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n22485), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n22485), .I0(n2398), .I1(n2423), .CO(n22486));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n22484), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut_4_lut (.I0(n50_adj_4369), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n28318));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_CARRY mod_5_add_1674_13 (.CI(n22484), .I0(n2399), .I1(n2423), .CO(n22485));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n22483), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n22483), .I0(n2400), .I1(n2423), .CO(n22484));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n22482), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n22482), .I0(n2401), .I1(n2423), .CO(n22483));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n22481), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n22481), .I0(n2402), .I1(n2423), .CO(n22482));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n22480), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n22480), .I0(n2403), .I1(n2423), .CO(n22481));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n22479), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n22479), .I0(n2404), .I1(n2423), .CO(n22480));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n22478), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n22478), .I0(n2405), .I1(n2423), .CO(n22479));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n22477), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n22477), .I0(n2406), .I1(n2423), .CO(n22478));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n22476), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n22476), .I0(n2407), .I1(n2423), .CO(n22477));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n22475), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n21936), .I0(bit_ctr[23]), .I1(GND_net), .CO(n21937));
    SB_CARRY mod_5_add_1674_4 (.CI(n22475), .I0(n2408), .I1(n2423), .CO(n22476));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n30269), 
            .I3(n22474), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n14865));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i25154_4_lut (.I0(one_wire_N_399[2]), .I1(n28326), .I2(n4_adj_4400), 
            .I3(n26073), .O(n27007));
    defparam i25154_4_lut.LUT_INIT = 16'hcecf;
    SB_CARRY mod_5_add_1674_3 (.CI(n22474), .I0(n2409), .I1(n30269), .CO(n22475));
    SB_LUT4 i23264_2_lut_4_lut (.I0(\state[1] ), .I1(start), .I2(\one_wire_N_399[11] ), 
            .I3(n110), .O(n28326));
    defparam i23264_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n30269), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n30269), 
            .CO(n22474));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n21935), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21797_2_lut_3_lut (.I0(\state[1] ), .I1(start), .I2(\one_wire_N_399[11] ), 
            .I3(GND_net), .O(n26854));
    defparam i21797_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_21_24 (.CI(n21935), .I0(bit_ctr[22]), .I1(GND_net), .CO(n21936));
    SB_CARRY add_21_10 (.CI(n21921), .I0(bit_ctr[8]), .I1(GND_net), .CO(n21922));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n21934), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n22473), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n22472), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n22472), .I0(n2292), .I1(n2324), .CO(n22473));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n22471), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n22471), .I0(n2293), .I1(n2324), .CO(n22472));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n22470), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n22470), .I0(n2294), .I1(n2324), .CO(n22471));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n22469), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n22469), .I0(n2295), .I1(n2324), .CO(n22470));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n22468), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n22468), .I0(n2296), .I1(n2324), .CO(n22469));
    SB_CARRY add_21_23 (.CI(n21934), .I0(bit_ctr[21]), .I1(GND_net), .CO(n21935));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n21933), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n22467), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut_4_lut_adj_1547 (.I0(n26736), .I1(n12135), .I2(n807), 
            .I3(bit_ctr[27]), .O(n838));
    defparam i3_4_lut_4_lut_adj_1547.LUT_INIT = 16'h0405;
    SB_CARRY mod_5_add_1607_15 (.CI(n22467), .I0(n2297), .I1(n2324), .CO(n22468));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n21914), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n21920), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n22466), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n19068), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n23695));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(n19068), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(bit_ctr[29]), .O(n708));
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hb60c;
    SB_CARRY mod_5_add_1607_14 (.CI(n22466), .I0(n2298), .I1(n2324), .CO(n22467));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n22465), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n22465), .I0(n2299), .I1(n2324), .CO(n22466));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n22464), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n22464), .I0(n2300), .I1(n2324), .CO(n22465));
    SB_CARRY add_21_22 (.CI(n21933), .I0(bit_ctr[20]), .I1(GND_net), .CO(n21934));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n22463), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n22463), .I0(n2301), .I1(n2324), .CO(n22464));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n22462), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n21932), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n22462), .I0(n2302), .I1(n2324), .CO(n22463));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n22461), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_399[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n22168), .O(n22_adj_4381)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1607_9 (.CI(n22461), .I0(n2303), .I1(n2324), .CO(n22462));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n22460), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n22460), .I0(n2304), .I1(n2324), .CO(n22461));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n22459), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n22459), .I0(n2305), .I1(n2324), .CO(n22460));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n22458), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17091_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_456 ));   // verilog/neopixel.v(16[20:25])
    defparam i17091_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY mod_5_add_1607_6 (.CI(n22458), .I0(n2306), .I1(n2324), .CO(n22459));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n22457), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n22457), .I0(n2307), .I1(n2324), .CO(n22458));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n22456), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n22456), .I0(n2308), .I1(n2324), .CO(n22457));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n30270), 
            .I3(n22455), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n22455), .I0(n2309), .I1(n30270), .CO(n22456));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n30270), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n30270), 
            .CO(n22455));
    SB_LUT4 i3034_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n26736), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3034_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n22454), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n22453), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n22453), .I0(n2193), .I1(n2225), .CO(n22454));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n22452), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n22452), .I0(n2194), .I1(n2225), .CO(n22453));
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_399[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n22167), .O(n23_adj_4379)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i15271_2_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n19068));
    defparam i15271_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n22451), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n22451), .I0(n2195), .I1(n2225), .CO(n22452));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n22450), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n22450), .I0(n2196), .I1(n2225), .CO(n22451));
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n14635), 
            .D(n255[12]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n22449), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n14635), 
            .D(n255[11]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n14635), 
            .D(n255[27]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_15 (.CI(n22449), .I0(n2197), .I1(n2225), .CO(n22450));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n22448), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n22448), .I0(n2198), .I1(n2225), .CO(n22449));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n22447), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n22447), .I0(n2199), .I1(n2225), .CO(n22448));
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n14864));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n14635), 
            .D(n255[26]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n14635), 
            .D(n255[25]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n14635), 
            .D(n255[10]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n22446), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n22446), .I0(n2200), .I1(n2225), .CO(n22447));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n22445), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n22445), .I0(n2201), .I1(n2225), .CO(n22446));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n22444), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n22444), .I0(n2202), .I1(n2225), .CO(n22445));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n22443), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n22443), .I0(n2203), .I1(n2225), .CO(n22444));
    SB_LUT4 i2_2_lut (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n22442), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n22442), .I0(n2204), .I1(n2225), .CO(n22443));
    SB_LUT4 i12_4_lut_adj_1548 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4410));
    defparam i12_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n22441), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n14635), 
            .D(n255[9]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n14635), 
            .D(n255[24]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1540_7 (.CI(n22441), .I0(n2205), .I1(n2225), .CO(n22442));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n22440), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n14863));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1540_6 (.CI(n22440), .I0(n2206), .I1(n2225), .CO(n22441));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n22439), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n22439), .I0(n2207), .I1(n2225), .CO(n22440));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n22438), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n22438), .I0(n2208), .I1(n2225), .CO(n22439));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n30271), 
            .I3(n22437), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n22437), .I0(n2209), .I1(n30271), .CO(n22438));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n30271), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n30271), 
            .CO(n22437));
    SB_CARRY sub_14_add_2_32 (.CI(n22167), .I0(timer[30]), .I1(n1[30]), 
            .CO(n22168));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_399[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n22166), .O(n28_adj_4377)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i10_4_lut_adj_1549 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4411));
    defparam i10_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1550 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4412));
    defparam i11_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i24614_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n14692));
    defparam i24614_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_CARRY sub_14_add_2_31 (.CI(n22166), .I0(timer[29]), .I1(n1[29]), 
            .CO(n22167));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_399[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n22165), .O(n26_adj_4375)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i25217_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30281));
    defparam i25217_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_30 (.CI(n22165), .I0(timer[28]), .I1(n1[28]), 
            .CO(n22166));
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i9_4_lut_adj_1551 (.I0(bit_ctr[15]), .I1(n18), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4413));
    defparam i9_4_lut_adj_1551.LUT_INIT = 16'hfefc;
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n14861));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n14860));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n14859));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n14858));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n14857));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n14856));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n14855));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n14854));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n14853));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n14852));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n14851));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n14850));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n14849));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n14848));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n14847));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n14846));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n14845));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n14844));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n14843));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n14842));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n14841));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n14840));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n14839));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n12));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n22416), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n22415), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n22415), .I0(n906), .I1(VCC_net), .CO(n22416));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n26828), .I2(VCC_net), 
            .I3(n22414), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n22414), .I0(n26828), .I1(VCC_net), 
            .CO(n22415));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n14692), .I2(VCC_net), 
            .I3(n22413), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n22413), .I0(n14692), .I1(VCC_net), 
            .CO(n22414));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_399[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n22164), .O(n21_adj_4376)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n12133), .I2(GND_net), 
            .I3(n22412), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n22412), .I0(n12133), .I1(GND_net), 
            .CO(n22413));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n22412));
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n25063));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_29 (.CI(n22164), .I0(timer[27]), .I1(n1[27]), 
            .CO(n22165));
    SB_CARRY add_21_9 (.CI(n21920), .I0(bit_ctr[7]), .I1(GND_net), .CO(n21921));
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut_adj_1552 (.I0(n25_adj_4413), .I1(n27_adj_4412), .I2(n26_adj_4411), 
            .I3(n28_adj_4410), .O(n2027));
    defparam i15_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1122_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n22373), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1122_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n22372), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_32 (.CI(n22372), .I0(GND_net), .I1(timer[30]), 
            .CO(n22373));
    SB_LUT4 timer_1122_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n22371), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_31 (.CI(n22371), .I0(GND_net), .I1(timer[29]), 
            .CO(n22372));
    SB_LUT4 timer_1122_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n22370), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_30 (.CI(n22370), .I0(GND_net), .I1(timer[28]), 
            .CO(n22371));
    SB_LUT4 timer_1122_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n22369), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_29 (.CI(n22369), .I0(GND_net), .I1(timer[27]), 
            .CO(n22370));
    SB_LUT4 timer_1122_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n22368), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1122_add_4_28 (.CI(n22368), .I0(GND_net), .I1(timer[26]), 
            .CO(n22369));
    SB_LUT4 timer_1122_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n22367), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_27 (.CI(n22367), .I0(GND_net), .I1(timer[25]), 
            .CO(n22368));
    SB_LUT4 timer_1122_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n22366), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_26 (.CI(n22366), .I0(GND_net), .I1(timer[24]), 
            .CO(n22367));
    SB_LUT4 timer_1122_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n22365), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_25 (.CI(n22365), .I0(GND_net), .I1(timer[23]), 
            .CO(n22366));
    SB_LUT4 timer_1122_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n22364), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_24 (.CI(n22364), .I0(GND_net), .I1(timer[22]), 
            .CO(n22365));
    SB_LUT4 timer_1122_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n22363), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_23 (.CI(n22363), .I0(GND_net), .I1(timer[21]), 
            .CO(n22364));
    SB_LUT4 timer_1122_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n22362), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_22 (.CI(n22362), .I0(GND_net), .I1(timer[20]), 
            .CO(n22363));
    SB_LUT4 timer_1122_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n22361), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_21 (.CI(n22361), .I0(GND_net), .I1(timer[19]), 
            .CO(n22362));
    SB_LUT4 timer_1122_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n22360), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_20 (.CI(n22360), .I0(GND_net), .I1(timer[18]), 
            .CO(n22361));
    SB_LUT4 timer_1122_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n22359), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_19 (.CI(n22359), .I0(GND_net), .I1(timer[17]), 
            .CO(n22360));
    SB_LUT4 timer_1122_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n22358), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_18 (.CI(n22358), .I0(GND_net), .I1(timer[16]), 
            .CO(n22359));
    SB_LUT4 timer_1122_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n22357), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_17 (.CI(n22357), .I0(GND_net), .I1(timer[15]), 
            .CO(n22358));
    SB_LUT4 timer_1122_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n22356), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_16 (.CI(n22356), .I0(GND_net), .I1(timer[14]), 
            .CO(n22357));
    SB_LUT4 timer_1122_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n22355), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_15 (.CI(n22355), .I0(GND_net), .I1(timer[13]), 
            .CO(n22356));
    SB_LUT4 timer_1122_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n22354), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_14 (.CI(n22354), .I0(GND_net), .I1(timer[12]), 
            .CO(n22355));
    SB_LUT4 timer_1122_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n22353), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_13 (.CI(n22353), .I0(GND_net), .I1(timer[11]), 
            .CO(n22354));
    SB_LUT4 timer_1122_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n22352), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_12 (.CI(n22352), .I0(GND_net), .I1(timer[10]), 
            .CO(n22353));
    SB_LUT4 timer_1122_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n22351), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_11 (.CI(n22351), .I0(GND_net), .I1(timer[9]), 
            .CO(n22352));
    SB_LUT4 timer_1122_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n22350), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_10 (.CI(n22350), .I0(GND_net), .I1(timer[8]), 
            .CO(n22351));
    SB_LUT4 timer_1122_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n22349), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_9 (.CI(n22349), .I0(GND_net), .I1(timer[7]), 
            .CO(n22350));
    SB_LUT4 timer_1122_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n22348), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_8 (.CI(n22348), .I0(GND_net), .I1(timer[6]), 
            .CO(n22349));
    SB_LUT4 timer_1122_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n22347), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n14635), 
            .D(n255[23]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_1122_add_4_7 (.CI(n22347), .I0(GND_net), .I1(timer[5]), 
            .CO(n22348));
    SB_LUT4 timer_1122_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n22346), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_6 (.CI(n22346), .I0(GND_net), .I1(timer[4]), 
            .CO(n22347));
    SB_LUT4 timer_1122_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n22345), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_5 (.CI(n22345), .I0(GND_net), .I1(timer[3]), 
            .CO(n22346));
    SB_LUT4 timer_1122_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n22344), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_4 (.CI(n22344), .I0(GND_net), .I1(timer[2]), 
            .CO(n22345));
    SB_LUT4 timer_1122_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n22343), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_3 (.CI(n22343), .I0(GND_net), .I1(timer[1]), 
            .CO(n22344));
    SB_LUT4 timer_1122_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1122_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1122_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n22343));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_c), .I1(n4_c), .I2(n1037), .I3(n22342), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n22341), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n22341), .I0(n1005), .I1(n1037), .CO(n22342));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n22340), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_21 (.CI(n21932), .I0(bit_ctr[19]), .I1(GND_net), .CO(n21933));
    SB_CARRY mod_5_add_736_6 (.CI(n22340), .I0(n1006), .I1(n1037), .CO(n22341));
    SB_LUT4 i11_4_lut_adj_1553 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4419));
    defparam i11_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19_adj_4420));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1554 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4421));
    defparam i1_2_lut_adj_1554.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n22339), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n22339), .I0(n1007), .I1(n1037), .CO(n22340));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n22338), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n22338), .I0(n1008), .I1(n1037), .CO(n22339));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n30272), 
            .I3(n22337), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n22337), .I0(n1009), .I1(n30272), .CO(n22338));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n30272), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n30272), 
            .CO(n22337));
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n21931), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n21931), .I0(bit_ctr[18]), .I1(GND_net), .CO(n21932));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n22336), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n22335), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n21930), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_8 (.CI(n22335), .I0(n1104), .I1(n1136), .CO(n22336));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n22334), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n22334), .I0(n1105), .I1(n1136), .CO(n22335));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n22333), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n22333), .I0(n1106), .I1(n1136), .CO(n22334));
    SB_LUT4 i9_4_lut_adj_1555 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4422));
    defparam i9_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n22332), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut_adj_1556 (.I0(n19_adj_4420), .I1(n26_adj_4419), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4423));
    defparam i13_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_803_5 (.CI(n22332), .I0(n1107), .I1(n1136), .CO(n22333));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n22331), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n22331), .I0(n1108), .I1(n1136), .CO(n22332));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n30273), 
            .I3(n22330), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i14_4_lut_adj_1557 (.I0(n1896), .I1(n28_adj_4423), .I2(n24_adj_4422), 
            .I3(n16_adj_4421), .O(n1928));
    defparam i14_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_803_3 (.CI(n22330), .I0(n1109), .I1(n30273), .CO(n22331));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n30273), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n30273), 
            .CO(n22330));
    SB_CARRY add_21_19 (.CI(n21930), .I0(bit_ctr[17]), .I1(GND_net), .CO(n21931));
    SB_LUT4 i25216_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30280));
    defparam i25216_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n22329), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n22328), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1558 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4428));
    defparam i10_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_4429));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1559 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_4430));
    defparam i9_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1560 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4431));
    defparam i7_3_lut_adj_1560.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1561 (.I0(n21_adj_4431), .I1(n23_adj_4430), .I2(n22_adj_4429), 
            .I3(n24_adj_4428), .O(n1829));
    defparam i13_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i25215_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30279));
    defparam i25215_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1562 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_4434));
    defparam i4_3_lut_adj_1562.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1563 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4435));
    defparam i8_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1564 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4436));
    defparam i7_3_lut_adj_1564.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1565 (.I0(n21_adj_4435), .I1(n17_adj_4434), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4437));
    defparam i11_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1566 (.I0(n1700), .I1(n24_adj_4437), .I2(n20_adj_4436), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_DFF timer_1122__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i25214_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30278));
    defparam i25214_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24693_4_lut (.I0(n28), .I1(n26858), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n29508));
    defparam i24693_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i24268_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n29331));
    defparam i24268_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24489_2_lut_4_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n24472), 
            .I3(LED_c), .O(n29304));   // verilog/neopixel.v(16[20:25])
    defparam i24489_2_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1567 (.I0(start), .I1(\one_wire_N_399[11] ), 
            .I2(n26858), .I3(GND_net), .O(n83));
    defparam i1_2_lut_3_lut_adj_1567.LUT_INIT = 16'habab;
    SB_LUT4 i55_4_lut (.I0(n26774), .I1(n50_adj_4369), .I2(\state[1] ), 
            .I3(n26858), .O(n26884));
    defparam i55_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i58_4_lut (.I0(n26884), .I1(n26854), .I2(n29331), .I3(n29508), 
            .O(n26888));
    defparam i58_4_lut.LUT_INIT = 16'h0535;
    SB_CARRY mod_5_add_870_9 (.CI(n22328), .I0(n1203), .I1(n1235), .CO(n22329));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n22327), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n22327), .I0(n1204), .I1(n1235), .CO(n22328));
    SB_LUT4 i46_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_462 ));
    defparam i46_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n22326), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_870_7 (.CI(n22326), .I0(n1205), .I1(n1235), .CO(n22327));
    SB_CARRY add_21_3 (.CI(n21914), .I0(bit_ctr[1]), .I1(GND_net), .CO(n21915));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n22325), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n22325), .I0(n1206), .I1(n1235), .CO(n22326));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n22324), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n22324), .I0(n1207), .I1(n1235), .CO(n22325));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n22323), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n22323), .I0(n1208), .I1(n1235), .CO(n22324));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n30274), 
            .I3(n22322), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n22322), .I0(n1209), .I1(n30274), .CO(n22323));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n30274), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n30274), 
            .CO(n22322));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n22321), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n22320), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n22320), .I0(n1302), .I1(n1334), .CO(n22321));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n22319), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n22319), .I0(n1303), .I1(n1334), .CO(n22320));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n21919), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n22318), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n22318), .I0(n1304), .I1(n1334), .CO(n22319));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n22317), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n21919), .I0(bit_ctr[6]), .I1(GND_net), .CO(n21920));
    SB_CARRY mod_5_add_937_7 (.CI(n22317), .I0(n1305), .I1(n1334), .CO(n22318));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n22316), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n21929), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_6 (.CI(n22316), .I0(n1306), .I1(n1334), .CO(n22317));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n22315), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n22315), .I0(n1307), .I1(n1334), .CO(n22316));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n22163), .O(one_wire_N_399[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n22314), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n22314), .I0(n1308), .I1(n1334), .CO(n22315));
    SB_CARRY sub_14_add_2_28 (.CI(n22163), .I0(timer[26]), .I1(n1[26]), 
            .CO(n22164));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n22162), .O(one_wire_N_399[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_27 (.CI(n22162), .I0(timer[25]), .I1(n1[25]), 
            .CO(n22163));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n22161), .O(one_wire_N_399[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_26 (.CI(n22161), .I0(timer[24]), .I1(n1[24]), 
            .CO(n22162));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_399[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n22160), .O(n30_adj_4378)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n22160), .I0(timer[23]), .I1(n1[23]), 
            .CO(n22161));
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_399[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n22159), .O(n24_adj_4382)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n22159), .I0(timer[22]), .I1(n1[22]), 
            .CO(n22160));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_399[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n22158), .O(n25_adj_4372)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n30275), 
            .I3(n22313), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n22313), .I0(n1309), .I1(n30275), .CO(n22314));
    SB_CARRY sub_14_add_2_23 (.CI(n22158), .I0(timer[21]), .I1(n1[21]), 
            .CO(n22159));
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n14635), 
            .D(n255[22]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n30275), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n30275), 
            .CO(n22313));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n22312), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_399[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n22157), .O(n29_adj_4374)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n14635), 
            .D(n255[21]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n14635), 
            .D(n255[20]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n14635), 
            .D(n255[19]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n7_adj_4445), 
            .D(state_3__N_248[0]), .S(n14750));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n14635), 
            .D(n255[18]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n22311), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n22311), .I0(n1401), .I1(n1433), .CO(n22312));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n22310), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n22310), .I0(n1402), .I1(n1433), .CO(n22311));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n22309), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n22309), .I0(n1403), .I1(n1433), .CO(n22310));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n22308), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n22308), .I0(n1404), .I1(n1433), .CO(n22309));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n22307), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n22307), .I0(n1405), .I1(n1433), .CO(n22308));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n22306), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n22306), .I0(n1406), .I1(n1433), .CO(n22307));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n22305), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_22 (.CI(n22157), .I0(timer[20]), .I1(n1[20]), 
            .CO(n22158));
    SB_CARRY mod_5_add_1004_5 (.CI(n22305), .I0(n1407), .I1(n1433), .CO(n22306));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n22304), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n22304), .I0(n1408), .I1(n1433), .CO(n22305));
    SB_CARRY add_21_18 (.CI(n21929), .I0(bit_ctr[16]), .I1(GND_net), .CO(n21930));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n30276), 
            .I3(n22303), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n22303), .I0(n1409), .I1(n30276), .CO(n22304));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n30276), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n22156), .O(one_wire_N_399[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n30276), 
            .CO(n22303));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n22302), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n22301), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n22301), .I0(n1500), .I1(n1532), .CO(n22302));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n22300), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n22300), .I0(n1501), .I1(n1532), .CO(n22301));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n22299), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n22299), .I0(n1502), .I1(n1532), .CO(n22300));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n22298), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1122__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1071_9 (.CI(n22298), .I0(n1503), .I1(n1532), .CO(n22299));
    SB_CARRY sub_14_add_2_21 (.CI(n22156), .I0(timer[19]), .I1(n1[19]), 
            .CO(n22157));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n22297), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n22297), .I0(n1504), .I1(n1532), .CO(n22298));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n22296), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n22296), .I0(n1505), .I1(n1532), .CO(n22297));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n22295), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n22295), .I0(n1506), .I1(n1532), .CO(n22296));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n22294), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n22155), .O(one_wire_N_399[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n22155), .I0(timer[18]), .I1(n1[18]), 
            .CO(n22156));
    SB_CARRY mod_5_add_1071_5 (.CI(n22294), .I0(n1507), .I1(n1532), .CO(n22295));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n22293), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n22293), .I0(n1508), .I1(n1532), .CO(n22294));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_399[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n22154), .O(n27_adj_4373)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n30277), 
            .I3(n22292), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n22292), .I0(n1509), .I1(n30277), .CO(n22293));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n30277), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n30277), 
            .CO(n22292));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n22291), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n22290), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n22290), .I0(n1599), .I1(n1631), .CO(n22291));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n22289), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n22289), .I0(n1600), .I1(n1631), .CO(n22290));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n21918), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n22288), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n22288), .I0(n1601), .I1(n1631), .CO(n22289));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n22287), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n22287), .I0(n1602), .I1(n1631), .CO(n22288));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n22286), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n22286), .I0(n1603), .I1(n1631), .CO(n22287));
    SB_CARRY sub_14_add_2_19 (.CI(n22154), .I0(timer[17]), .I1(n1[17]), 
            .CO(n22155));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n22285), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n22285), .I0(n1604), .I1(n1631), .CO(n22286));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n22284), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n22284), .I0(n1605), .I1(n1631), .CO(n22285));
    SB_DFF timer_1122__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1122__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n22283), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_4_lut_adj_1568 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4449));
    defparam i8_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1569 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4450));
    defparam i1_3_lut_adj_1569.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4451));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1570 (.I0(n13_adj_4450), .I1(n20_adj_4449), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4452));
    defparam i10_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1571 (.I0(n1601), .I1(n22_adj_4452), .I2(n18_adj_4451), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n14817));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i25213_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30277));
    defparam i25213_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1572 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4453));
    defparam i7_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_6 (.CI(n22283), .I0(n1606), .I1(n1631), .CO(n22284));
    SB_LUT4 i9_4_lut_adj_1573 (.I0(n1504), .I1(n18_adj_4453), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4454));
    defparam i9_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n22282), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4_3_lut_adj_1574 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4455));
    defparam i4_3_lut_adj_1574.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1138_5 (.CI(n22282), .I0(n1607), .I1(n1631), .CO(n22283));
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n22153), .O(one_wire_N_399[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n22281), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n21928), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_4 (.CI(n22281), .I0(n1608), .I1(n1631), .CO(n22282));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n26888), .D(\neo_pixel_transmitter.done_N_462 ), 
            .R(n28318));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n30278), 
            .I3(n22280), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n22280), .I0(n1609), .I1(n30278), .CO(n22281));
    SB_CARRY sub_14_add_2_18 (.CI(n22153), .I0(timer[16]), .I1(n1[16]), 
            .CO(n22154));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n30278), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n30278), 
            .CO(n22280));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n22279), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n22278), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n22278), .I0(n1698), .I1(n1730), .CO(n22279));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n22277), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n22277), .I0(n1699), .I1(n1730), .CO(n22278));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n22276), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n22276), .I0(n1700), .I1(n1730), .CO(n22277));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n22275), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n22275), .I0(n1701), .I1(n1730), .CO(n22276));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n22274), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n22274), .I0(n1702), .I1(n1730), .CO(n22275));
    SB_LUT4 i10_4_lut_adj_1575 (.I0(n15_adj_4455), .I1(n20_adj_4454), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n22273), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n22273), .I0(n1703), .I1(n1730), .CO(n22274));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n22152), .O(one_wire_N_399[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n22272), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_17 (.CI(n22152), .I0(timer[15]), .I1(n1[15]), 
            .CO(n22153));
    SB_LUT4 i25212_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30276));
    defparam i25212_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_8 (.CI(n22272), .I0(n1704), .I1(n1730), .CO(n22273));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n22271), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24_4_lut_adj_1576 (.I0(n50_adj_4369), .I1(n20817), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n10_adj_4456));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_4_lut_adj_1576.LUT_INIT = 16'h0ac0;
    SB_LUT4 i23_4_lut_adj_1577 (.I0(n10_adj_4456), .I1(n29213), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n14750));   // verilog/neopixel.v(35[12] 117[6])
    defparam i23_4_lut_adj_1577.LUT_INIT = 16'h0aca;
    SB_CARRY mod_5_add_1205_7 (.CI(n22271), .I0(n1705), .I1(n1730), .CO(n22272));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n22151), .O(one_wire_N_399[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n22270), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_3_lut (.I0(n20822), .I1(n26778), .I2(\state[1] ), .I3(GND_net), 
            .O(n7_adj_4445));
    defparam i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2239_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n23391), 
            .I3(GND_net), .O(color_bit_N_442[4]));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2239_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i24532_4_lut (.I0(n30460), .I1(n23679), .I2(n30388), .I3(bit_ctr[2]), 
            .O(n29281));
    defparam i24532_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(state_3__N_248[1]), .I1(n30358), .I2(n29281), 
            .I3(color_bit_N_442[4]), .O(state_3__N_248[0]));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'h5044;
    SB_CARRY sub_14_add_2_16 (.CI(n22151), .I0(timer[14]), .I1(n1[14]), 
            .CO(n22152));
    SB_CARRY mod_5_add_1205_6 (.CI(n22270), .I0(n1706), .I1(n1730), .CO(n22271));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n22269), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n22269), .I0(n1707), .I1(n1730), .CO(n22270));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n22268), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n22268), .I0(n1708), .I1(n1730), .CO(n22269));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n30279), 
            .I3(n22267), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_3 (.CI(n22267), .I0(n1709), .I1(n30279), .CO(n22268));
    SB_LUT4 i15501_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n19303));
    defparam i15501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n30279), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n30279), 
            .CO(n22267));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n22266), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n22265), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n22265), .I0(n1797), .I1(n1829), .CO(n22266));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n22264), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n22264), .I0(n1798), .I1(n1829), .CO(n22265));
    SB_LUT4 i6_4_lut_adj_1579 (.I0(n1405), .I1(n19303), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4457));
    defparam i6_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n22263), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1580 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4458));
    defparam i7_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1581 (.I0(n17_adj_4458), .I1(n1408), .I2(n16_adj_4457), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 i25211_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30275));
    defparam i25211_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n22150), .O(one_wire_N_399[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n22150), .I0(timer[13]), .I1(n1[13]), 
            .CO(n22151));
    SB_CARRY mod_5_add_1272_13 (.CI(n22263), .I0(n1799), .I1(n1829), .CO(n22264));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n22149), .O(one_wire_N_399[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n22262), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n22262), .I0(n1800), .I1(n1829), .CO(n22263));
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n22261), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n22261), .I0(n1801), .I1(n1829), .CO(n22262));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n22260), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n22260), .I0(n1802), .I1(n1829), .CO(n22261));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n22259), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4459));
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1272_9 (.CI(n22259), .I0(n1803), .I1(n1829), .CO(n22260));
    SB_CARRY sub_14_add_2_14 (.CI(n22149), .I0(timer[12]), .I1(n1[12]), 
            .CO(n22150));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n22148), .O(\one_wire_N_399[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_3_lut_adj_1583 (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), 
            .I3(GND_net), .O(n12_adj_4460));
    defparam i3_3_lut_adj_1583.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n22258), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_13 (.CI(n22148), .I0(timer[11]), .I1(n1[11]), 
            .CO(n22149));
    SB_CARRY mod_5_add_1272_8 (.CI(n22258), .I0(n1804), .I1(n1829), .CO(n22259));
    SB_LUT4 i7_4_lut_adj_1584 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4459), 
            .O(n16_adj_4461));
    defparam i7_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1585 (.I0(n1307), .I1(n16_adj_4461), .I2(n12_adj_4460), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i25210_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30274));
    defparam i25210_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_17 (.CI(n21928), .I0(bit_ctr[15]), .I1(GND_net), .CO(n21929));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n22257), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n22257), .I0(n1805), .I1(n1829), .CO(n22258));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n22256), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n22147), .O(one_wire_N_399[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n22147), .I0(timer[10]), .I1(n1[10]), 
            .CO(n22148));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n22146), .O(one_wire_N_399[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n22146), .I0(timer[9]), .I1(n1[9]), 
            .CO(n22147));
    SB_CARRY mod_5_add_1272_6 (.CI(n22256), .I0(n1806), .I1(n1829), .CO(n22257));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n22255), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n22255), .I0(n1807), .I1(n1829), .CO(n22256));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n22254), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n21927), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_4 (.CI(n22254), .I0(n1808), .I1(n1829), .CO(n22255));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n30280), 
            .I3(n22253), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_16 (.CI(n21927), .I0(bit_ctr[14]), .I1(GND_net), .CO(n21928));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n21926), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n21926), .I0(bit_ctr[13]), .I1(GND_net), .CO(n21927));
    SB_CARRY mod_5_add_1272_3 (.CI(n22253), .I0(n1809), .I1(n30280), .CO(n22254));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n30280), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n30280), 
            .CO(n22253));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n22252), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n22251), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n22251), .I0(n1896), .I1(n1928), .CO(n22252));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n22250), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n22250), .I0(n1897), .I1(n1928), .CO(n22251));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n22249), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_7 (.CI(n21918), .I0(bit_ctr[5]), .I1(GND_net), .CO(n21919));
    SB_CARRY mod_5_add_1339_14 (.CI(n22249), .I0(n1898), .I1(n1928), .CO(n22250));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n22248), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n22248), .I0(n1899), .I1(n1928), .CO(n22249));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n22247), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n22247), .I0(n1900), .I1(n1928), .CO(n22248));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n22246), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_399[9]), .I1(timer[8]), 
            .I2(n1[8]), .I3(n22145), .O(n7_adj_4387)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_10 (.CI(n22145), .I0(timer[8]), .I1(n1[8]), 
            .CO(n22146));
    SB_LUT4 sub_14_add_2_9_lut (.I0(one_wire_N_399[5]), .I1(timer[7]), .I2(n1[7]), 
            .I3(n22144), .O(n8_adj_4388)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1339_11 (.CI(n22246), .I0(n1901), .I1(n1928), .CO(n22247));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n22245), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n22245), .I0(n1902), .I1(n1928), .CO(n22246));
    SB_CARRY sub_14_add_2_9 (.CI(n22144), .I0(timer[7]), .I1(n1[7]), .CO(n22145));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n22244), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_8_lut (.I0(n44_adj_4383), .I1(timer[6]), .I2(n1[6]), 
            .I3(n22143), .O(n9_adj_4386)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1339_9 (.CI(n22244), .I0(n1903), .I1(n1928), .CO(n22245));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n22243), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_8 (.CI(n22143), .I0(timer[6]), .I1(n1[6]), .CO(n22144));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n22142), .O(one_wire_N_399[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n22142), .I0(timer[5]), .I1(n1[5]), .CO(n22143));
    SB_CARRY mod_5_add_1339_8 (.CI(n22243), .I0(n1904), .I1(n1928), .CO(n22244));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n22242), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n22242), .I0(n1905), .I1(n1928), .CO(n22243));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n22241), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n22241), .I0(n1906), .I1(n1928), .CO(n22242));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n22240), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n22240), .I0(n1907), .I1(n1928), .CO(n22241));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n22239), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n22239), .I0(n1908), .I1(n1928), .CO(n22240));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n30281), 
            .I3(n22238), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_3 (.CI(n22238), .I0(n1909), .I1(n30281), .CO(n22239));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n30281), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n30281), 
            .CO(n22238));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n21917), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n22141), .O(one_wire_N_399[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n21914));
    SB_CARRY sub_14_add_2_6 (.CI(n22141), .I0(timer[4]), .I1(n1[4]), .CO(n22142));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n22140), .O(one_wire_N_399[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n22140), .I0(timer[3]), .I1(n1[3]), .CO(n22141));
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n14635), 
            .D(n255[17]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n14635), 
            .D(n255[16]), .R(n14745));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_6 (.CI(n21917), .I0(bit_ctr[4]), .I1(GND_net), .CO(n21918));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n22139), .O(one_wire_N_399[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n21925), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n22066), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_14 (.CI(n21925), .I0(bit_ctr[12]), .I1(GND_net), .CO(n21926));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n22065), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, GND_net, clk32MHz, 
            data_o, n28236, reg_B, ENCODER1_A_c_1, VCC_net, n14836, 
            ENCODER1_B_c_0, n15348) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output n28236;
    output [1:0]reg_B;
    input ENCODER1_A_c_1;
    input VCC_net;
    input n14836;
    input ENCODER1_B_c_0;
    input n15348;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2422;
    
    wire n2399, n22137, n22136, n22135, n22134, n22133, count_enable, 
        B_delayed, A_delayed, n22132, n22131, n22130, n22129, n22128, 
        n22127, n22126, n22125, n22124, n22123, n22122, n22121, 
        n22120, n22119, n22118, n22117, n22116, n22115, count_direction, 
        n22114;
    
    SB_LUT4 add_526_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2399), 
            .I3(n22137), .O(n2422[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_526_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2399), 
            .I3(n22136), .O(n2422[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_24 (.CI(n22136), .I0(encoder1_position[22]), .I1(n2399), 
            .CO(n22137));
    SB_LUT4 add_526_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2399), 
            .I3(n22135), .O(n2422[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_23 (.CI(n22135), .I0(encoder1_position[21]), .I1(n2399), 
            .CO(n22136));
    SB_LUT4 add_526_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2399), 
            .I3(n22134), .O(n2422[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_22 (.CI(n22134), .I0(encoder1_position[20]), .I1(n2399), 
            .CO(n22135));
    SB_LUT4 add_526_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2399), 
            .I3(n22133), .O(n2422[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_21 (.CI(n22133), .I0(encoder1_position[19]), .I1(n2399), 
            .CO(n22134));
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_526_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2399), 
            .I3(n22132), .O(n2422[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_20 (.CI(n22132), .I0(encoder1_position[18]), .I1(n2399), 
            .CO(n22133));
    SB_LUT4 add_526_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2399), 
            .I3(n22131), .O(n2422[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_19 (.CI(n22131), .I0(encoder1_position[17]), .I1(n2399), 
            .CO(n22132));
    SB_LUT4 add_526_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2399), 
            .I3(n22130), .O(n2422[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_18 (.CI(n22130), .I0(encoder1_position[16]), .I1(n2399), 
            .CO(n22131));
    SB_LUT4 add_526_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2399), 
            .I3(n22129), .O(n2422[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_17 (.CI(n22129), .I0(encoder1_position[15]), .I1(n2399), 
            .CO(n22130));
    SB_LUT4 add_526_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2399), 
            .I3(n22128), .O(n2422[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_16 (.CI(n22128), .I0(encoder1_position[14]), .I1(n2399), 
            .CO(n22129));
    SB_LUT4 add_526_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2399), 
            .I3(n22127), .O(n2422[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_15 (.CI(n22127), .I0(encoder1_position[13]), .I1(n2399), 
            .CO(n22128));
    SB_LUT4 add_526_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2399), 
            .I3(n22126), .O(n2422[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_14 (.CI(n22126), .I0(encoder1_position[12]), .I1(n2399), 
            .CO(n22127));
    SB_LUT4 add_526_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2399), 
            .I3(n22125), .O(n2422[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_13 (.CI(n22125), .I0(encoder1_position[11]), .I1(n2399), 
            .CO(n22126));
    SB_LUT4 add_526_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2399), 
            .I3(n22124), .O(n2422[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_12 (.CI(n22124), .I0(encoder1_position[10]), .I1(n2399), 
            .CO(n22125));
    SB_LUT4 add_526_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2399), 
            .I3(n22123), .O(n2422[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_11 (.CI(n22123), .I0(encoder1_position[9]), .I1(n2399), 
            .CO(n22124));
    SB_LUT4 add_526_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2399), 
            .I3(n22122), .O(n2422[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_526_10 (.CI(n22122), .I0(encoder1_position[8]), .I1(n2399), 
            .CO(n22123));
    SB_LUT4 add_526_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2399), 
            .I3(n22121), .O(n2422[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_9 (.CI(n22121), .I0(encoder1_position[7]), .I1(n2399), 
            .CO(n22122));
    SB_LUT4 add_526_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2399), 
            .I3(n22120), .O(n2422[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_8 (.CI(n22120), .I0(encoder1_position[6]), .I1(n2399), 
            .CO(n22121));
    SB_LUT4 add_526_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2399), 
            .I3(n22119), .O(n2422[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_7 (.CI(n22119), .I0(encoder1_position[5]), .I1(n2399), 
            .CO(n22120));
    SB_LUT4 add_526_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2399), 
            .I3(n22118), .O(n2422[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_6 (.CI(n22118), .I0(encoder1_position[4]), .I1(n2399), 
            .CO(n22119));
    SB_LUT4 add_526_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2399), 
            .I3(n22117), .O(n2422[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_5 (.CI(n22117), .I0(encoder1_position[3]), .I1(n2399), 
            .CO(n22118));
    SB_LUT4 add_526_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2399), 
            .I3(n22116), .O(n2422[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_4 (.CI(n22116), .I0(encoder1_position[2]), .I1(n2399), 
            .CO(n22117));
    SB_LUT4 add_526_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2399), 
            .I3(n22115), .O(n2422[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_3 (.CI(n22115), .I0(encoder1_position[1]), .I1(n2399), 
            .CO(n22116));
    SB_LUT4 add_526_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n22114), .O(n2422[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_526_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_526_2 (.CI(n22114), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n22115));
    SB_CARRY add_526_1 (.CI(GND_net), .I0(n2399), .I1(n2399), .CO(n22114));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2422[23]));   // quad.v(35[10] 41[6])
    SB_LUT4 i860_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2399));   // quad.v(37[5] 40[8])
    defparam i860_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,100)  debounce (.n28236(n28236), .reg_B({reg_B}), .GND_net(GND_net), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .n14836(n14836), .data_o({data_o}), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n15348(n15348));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (n28236, reg_B, GND_net, ENCODER1_A_c_1, 
            clk32MHz, VCC_net, n14836, data_o, ENCODER1_B_c_0, n15348);
    output n28236;
    output [1:0]reg_B;
    input GND_net;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input VCC_net;
    input n14836;
    output [1:0]data_o;
    input ENCODER1_B_c_0;
    input n15348;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3576;
    wire [6:0]n33;
    
    wire n22436, n22435, n22434, n22433, n22432, n22431;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n28236));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n28236), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1129__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 cnt_reg_1129_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n22436), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1129_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n22435), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1129_add_4_7 (.CI(n22435), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n22436));
    SB_LUT4 cnt_reg_1129_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n22434), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1129_add_4_6 (.CI(n22434), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n22435));
    SB_LUT4 cnt_reg_1129_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n22433), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1129_add_4_5 (.CI(n22433), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n22434));
    SB_LUT4 cnt_reg_1129_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n22432), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1129_add_4_4 (.CI(n22432), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n22433));
    SB_LUT4 cnt_reg_1129_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n22431), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1129_add_4_3 (.CI(n22431), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n22432));
    SB_LUT4 cnt_reg_1129_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1129_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1129_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n22431));
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n14836));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n15348));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1129__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1129__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1129__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1129__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1129__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1129__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] , 
            \Kp[1] , \Kp[0] , \Kp[2] , \Kp[3] , \Kp[4] , \Kp[5] , 
            IntegralLimit, PWMLimit, \Ki[1] , \Ki[0] , \Ki[2] , \Ki[3] , 
            \Ki[4] , \Ki[5] , \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , 
            \Ki[10] , \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , 
            duty, n30261, VCC_net, clk32MHz, setpoint, motor_state) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input [23:0]IntegralLimit;
    input [23:0]PWMLimit;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    output [23:0]duty;
    output n30261;
    input VCC_net;
    input clk32MHz;
    input [23:0]setpoint;
    input [23:0]motor_state;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n22750;
    wire [17:0]n6641;
    
    wire n597, n22751;
    wire [18:0]n6620;
    
    wire n524, n22749;
    wire [23:0]n1;
    
    wire n463, n536, n609, n682, n755, n22013;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n22014, n451, n22748, n828, n901, n21950;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    wire [23:0]n2552;
    
    wire n21951, n378, n22747, n974, n1047, n1120, n101, n305, 
        n22746, n32, n174, n247, n320, n162, n393, n235, n466, 
        n539, n612, n685, n86, n758;
    wire [23:0]n1_adj_4303;
    
    wire n831, n308, n381, n454, n527, n600;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3392 ;
    
    wire n21949, n904, n977, n1050, n104, n35, n177, n250, n323, 
        n396, n469, n542, n615, n688, n761, n834, n907, n980, 
        n107, n38, n180, n253, n326, n399, n472, n545, n618, 
        n691, n764, n837, n910, n110, n41, n183, n256, n329, 
        n402, n475, n548, n621, n694, n767, n840, n113, n44, 
        n186, n259, n332, n673, n405, n478, n551, n624, n697, 
        n770, n116, n47, n189, n262, n335, n408, n481, n554, 
        n746, n819, n892, n627, n700, n119, n50, n192, n265, 
        n338, n411, n484, n557, n630, n232, n22745, n159, n22744, 
        n22219;
    wire [23:0]n1_adj_4304;
    
    wire n22220, n17_adj_3887, n122, n53;
    wire [19:0]n6598;
    
    wire n22743;
    wire [5:0]n7112;
    
    wire n27839, n490, n23147;
    wire [4:0]n7120;
    
    wire n417, n23146, n195_adj_3888, n344, n23145, n271, n23144, 
        n268, n198, n23143, n341, n56, n125;
    wire [6:0]n7103;
    
    wire n560, n23142, n414, n487, n23141, n414_adj_3889, n23140, 
        n341_adj_3891, n23139, n268_adj_3892, n23138, n195_adj_3893, 
        n23137, n53_adj_3894, n122_adj_3895;
    wire [7:0]n7093;
    
    wire n630_adj_3896, n23136, n557_adj_3897, n23135, n487_adj_3898, 
        n484_adj_3899, n23134, n411_adj_3900, n23133, n338_adj_3901, 
        n23132, n560_adj_3902, n265_adj_3903, n23131, n192_adj_3904, 
        n23130, n50_adj_3905, n119_adj_3906, n125_adj_3907;
    wire [8:0]n7082;
    
    wire n700_adj_3908, n23129, n627_adj_3909, n23128, n554_adj_3910, 
        n23127, n481_adj_3911, n23126, n408_adj_3912, n23125, n335_adj_3913, 
        n23124, n262_adj_3914, n23123, n189_adj_3915, n23122, n47_adj_3916, 
        n116_adj_3917, n56_adj_3918;
    wire [9:0]n7070;
    
    wire n770_adj_3919, n23121, n697_adj_3920, n23120, n198_adj_3921, 
        n624_adj_3922, n23119, n551_adj_3923, n23118, n478_adj_3924, 
        n23117, n271_adj_3925, n405_adj_3926, n23116, n332_adj_3927, 
        n23115, n259_adj_3928, n23114, n186_adj_3929, n23113, n44_adj_3930, 
        n113_adj_3931;
    wire [10:0]n7057;
    
    wire n840_adj_3932, n23112, n767_adj_3933, n23111, n694_adj_3934, 
        n23110, n621_adj_3935, n23109, n548_adj_3936, n23108, n475_adj_3937, 
        n23107, n402_adj_3938, n23106, n329_adj_3939, n23105, n344_adj_3940, 
        n256_adj_3941, n23104, n183_adj_3942, n23103, n41_adj_3943, 
        n110_adj_3944;
    wire [11:0]n7043;
    
    wire n910_adj_3945, n23102, n837_adj_3946, n23101, n764_adj_3947, 
        n23100, n691_adj_3948, n23099, n618_adj_3949, n23098, n965, 
        n545_adj_3950, n23097, n472_adj_3951, n23096, n1038, n399_adj_3952, 
        n23095, n326_adj_3953, n23094, n253_adj_3954, n23093, n180_adj_3955, 
        n23092, n38_adj_3956, n107_adj_3957;
    wire [12:0]n7028;
    
    wire n980_adj_3958, n23091, n907_adj_3959, n23090, n417_adj_3960, 
        n6;
    wire [3:0]n6830;
    wire [4:0]n6823;
    
    wire n834_adj_3961, n23089, n761_adj_3962, n23088, n688_adj_3963, 
        n23087, n615_adj_3964, n23086, n542_adj_3965, n23085, n469_adj_3966, 
        n23084, n396_adj_3967, n23083, n323_adj_3968, n23082, n250_adj_3969, 
        n23081, n177_adj_3970, n23080, n35_adj_3971, n104_adj_3972;
    wire [13:0]n7012;
    
    wire n1050_adj_3973, n23079, n977_adj_3974, n23078, n904_adj_3975, 
        n23077, n831_adj_3976, n23076, n758_adj_3977, n23075, n685_adj_3978, 
        n23074, n612_adj_3979, n23073, n539_adj_3980, n23072, n466_adj_3981, 
        n23071, n393_adj_3982, n23070, n320_adj_3983, n23069, n22742, 
        n1111;
    wire [23:0]duty_23__N_3492;
    
    wire n22012, n4;
    wire [2:0]n6836;
    wire [1:0]n6841;
    
    wire n247_adj_3985, n23068, n174_adj_3986, n23067, n32_adj_3987, 
        n101_adj_3988;
    wire [23:0]n257;
    
    wire n22218, n22741, n22740;
    wire [14:0]n6995;
    
    wire n1120_adj_3990, n23066, n22739, n1047_adj_3991, n23065, n1105, 
        n22738, n490_adj_3992, n12_adj_3994, n8_adj_3995, n22217, 
        n11_adj_3997, n6_adj_3998, n21754, n18_adj_3999, n13_adj_4000, 
        n4_adj_4001, n27634, n1032, n22737, n77, n8_adj_4002, n150, 
        n223, n959, n22736, n296, n369, n442, n515, n588, n661, 
        n734, n807, n880, n953, n1026, n1099, n974_adj_4003, n23064, 
        n77_adj_4005, n8_adj_4007, n150_adj_4008, n74, n5_adj_4009, 
        n886, n22735, n147_adj_4010, n220, n293, n366, n223_adj_4012, 
        n439, n512, n585, n658, n731, n296_adj_4013, n901_adj_4014, 
        n23063, n804, n369_adj_4015, n442_adj_4016, n515_adj_4017, 
        \PID_CONTROLLER.integral_23__N_3440 , n813, n22734, n588_adj_4019, 
        n877, n950, n661_adj_4021, n734_adj_4022, n1023, n1096, 
        n807_adj_4023, n880_adj_4024, n953_adj_4025, n1026_adj_4026, 
        n1099_adj_4027, n80, n11_adj_4029, n153, n226, n299, n74_adj_4030, 
        n5_adj_4031, n372, n445, n518, n591, n664, n740, n22733, 
        n667, n22732, n737, n810, n883, n147_adj_4032, n956, n1029, 
        n220_adj_4033, n1102, n293_adj_4034, n366_adj_4036, n439_adj_4037, 
        n512_adj_4038, n83, n14_adj_4040, n156, n229, n92, n585_adj_4042, 
        n302, n658_adj_4043, n23_adj_4045, n731_adj_4046, n804_adj_4047, 
        n375, n448, n521, n594, n667_adj_4048, n740_adj_4049, n877_adj_4051, 
        n813_adj_4053, n22216, n165, n886_adj_4055, n959_adj_4056, 
        n950_adj_4057, n1023_adj_4059, n1096_adj_4060, n1032_adj_4061, 
        n1105_adj_4062, n86_adj_4064, n17_adj_4065, n159_adj_4066, n232_adj_4067, 
        n305_adj_4068, n238, n311, n378_adj_4069, n384, n457, n451_adj_4070, 
        n828_adj_4071, n23062, n524_adj_4072, n530, n597_adj_4073, 
        n670, n743, n816, n889, n962, n1035, n1108, n89, n20_adj_4075, 
        n162_adj_4076, n603, n235_adj_4077, n308_adj_4078, n676, n381_adj_4079, 
        n454_adj_4080, n749, n527_adj_4081, n822, n600_adj_4082, n673_adj_4083, 
        n746_adj_4084, n819_adj_4085, n892_adj_4086, n965_adj_4087, 
        n1038_adj_4088, n1111_adj_4089, n895, n968, n1041, n23_adj_4090, 
        n594_adj_4091, n22731, n165_adj_4092, n1114, n238_adj_4093, 
        n311_adj_4094, n521_adj_4095, n22730, n384_adj_4096, n95, 
        n80_adj_4097, n11_adj_4099, n457_adj_4100, n26_adj_4101, n168, 
        n530_adj_4102, n241, n29535, n153_adj_4103, n603_adj_4104, 
        n755_adj_4105, n23061, n682_adj_4106, n23060, n448_adj_4107, 
        n22729, n609_adj_4108, n23059, n375_adj_4109, n22728, n536_adj_4110, 
        n23058, n463_adj_4111, n23057, n390, n23056, n317, n23055, 
        n314, n302_adj_4112, n22727, n244, n23054, n387, n171, 
        n23053, n29, n98, n229_adj_4113, n22726;
    wire [15:0]n6977;
    
    wire n23052, n156_adj_4114, n22725, n1117, n23051, n14_adj_4115, 
        n83_adj_4116, n1044, n23050, n971, n23049, n460, n22215, 
        n898, n23048, n825, n23047, n752, n23046, n679, n23045, 
        n533, n606, n679_adj_4119;
    wire [20:0]n6575;
    
    wire n22724, n752_adj_4120, n676_adj_4121, n825_adj_4122, n898_adj_4123, 
        n971_adj_4124, n1044_adj_4125, n22723, n22722, n606_adj_4126, 
        n23044, n1117_adj_4127, n98_adj_4128, n22011, n29_adj_4129, 
        n171_adj_4130, n22721, n244_adj_4131, n317_adj_4132, n390_adj_4133, 
        n22720, n226_adj_4134, n749_adj_4135, n299_adj_4136, n822_adj_4137, 
        n372_adj_4138, n6_adj_4139;
    wire [3:0]n7127;
    
    wire n22010, n445_adj_4141, n895_adj_4142, n204, n518_adj_4143, 
        n968_adj_4144, n11_adj_4145, n9_adj_4146, n29532, n591_adj_4147;
    wire [1:0]n7138;
    
    wire n533_adj_4148, n23043, n1041_adj_4149, n21952, n21948, n21695, 
        n1114_adj_4150, n131, n21729, n664_adj_4151, n737_adj_4152, 
        n62, n41_adj_4154, n39, n460_adj_4155, n23042, n45, n37, 
        n22719, n29_adj_4156, n31, n30983, n1102_adj_4157, n22718, 
        n43, n23_adj_4158, n25_adj_4159, n35_adj_4160, n11_adj_4161, 
        n29895, n17_adj_4162, n29778, n1029_adj_4163, n22717, n21953, 
        n13_adj_4164, n387_adj_4165, n23041, n92_adj_4166, n22009, 
        n956_adj_4168, n22716, n314_adj_4169, n23040, n15_adj_4170, 
        n27, n33, n9_adj_4171, n17_adj_4172, n883_adj_4173, n22715, 
        n19_adj_4174, n241_adj_4175, n23039, n168_adj_4176, n23038, 
        n21947, n26_adj_4177, n95_adj_4178;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3443 ;
    
    wire n22214, n810_adj_4179, n22714;
    wire [16:0]n6958;
    
    wire n23037, n21_adj_4180, n23036;
    wire [23:0]duty_23__N_3368;
    
    wire n45_adj_4181, n22213, n22713, n22712, n23035, n23034, n29424, 
        n22711, n29417, n23033, n12_adj_4182, n10_adj_4183, n30, 
        n22710, n23032, n22709, n29435, n29701, n29697, n30006, 
        n22708, n23031, n29847, n22707, n30060, n23030, n22706, 
        n16_adj_4184, n23029, n6_adj_4185, n29992, n23028, n22705, 
        n23027, n21946, n23026, n23025, n23024, n23023, n23022;
    wire [17:0]n6938;
    
    wire n23021, n23020, n23019, n23018, n23017, n23016, n23015, 
        n23014, n23013, n23012, n29993, n8_adj_4186, n24_adj_4187, 
        n29402, n29400, n29869, n29934, n23011, n4_adj_4188, n23010, 
        n29982, n23009, n23008, n23007, n23006, n4_adj_4189, n29983, 
        n29413, n29411, n30070, n29936, n30119, n30120, n30101, 
        n29404, n30024, n4_adj_4190;
    wire [2:0]n7133;
    
    wire n40, n23005, n30026, duty_23__N_3491, n39_adj_4192;
    wire [18:0]n6917;
    
    wire n23004, n22008, n41_adj_4193, n21652, n45_adj_4195, n43_adj_4196, 
        n23003, n43_adj_4197, n22212, n23002;
    wire [0:0]n4998;
    wire [21:0]n6551;
    
    wire n22704, n37_adj_4198, n22007, n23_adj_4199, n23001, n23000, 
        n22999, n25_adj_4200, n22998, n22997, n22996, n22995, n29_adj_4201, 
        n22994, n22993, n22992, n31_adj_4202, n22703, n35_adj_4203, 
        n33_adj_4205, n11_adj_4206, n13_adj_4207, n22991, n22702, 
        n22990, n22701, n15_adj_4208, n12_adj_4209, n27_adj_4211, 
        n22989, n22988, n9_adj_4212, n22987, n17_adj_4213, n22700;
    wire [19:0]n6895;
    
    wire n22986, n19_adj_4214, n22985, n22984, n22699, n41_adj_4215, 
        n22211, n22983, n22698, n22982, n22697, n21_adj_4217, n29388, 
        n29382, n22981, n22006, n22980, n8_adj_4219, n22696, n30965, 
        n12_adj_4220, n29776, n22695, n11_adj_4221, n39_adj_4222, 
        n22210, n29774, n22694, n22979, n22978, n22977, n30959, 
        n10_adj_4223, n37_adj_4224, n22209, n30_adj_4225, n27_adj_4226, 
        n15_adj_4227, n13_adj_4228, n11_adj_4229, n29455, n21_adj_4230, 
        n19_adj_4231, n17_adj_4232, n9_adj_4233, n29464, n16_adj_4234, 
        n22693, n29437, n8_adj_4235, n35_adj_4236, n22208, n22976, 
        n24_adj_4237, n29398, n29667, n29663, n29998, n29831, n6_adj_4238, 
        n30058, n16_adj_4239, n6_adj_4240, n29978, n29979, n8_adj_4241, 
        n24_adj_4242, n29368, n29366, n29871, n29940, n4_adj_4243, 
        n29976, n29977, n29378, n29376, n30072, n29942, n30121, 
        n21886, n30122, n30099, n29370, n30030, n22975, n22974, 
        n40_adj_4244, n22973, n22972, n30032, n7_adj_4245, n5_adj_4246, 
        n29496, n29746, n29742, n25_adj_4247, n23_adj_4248, n30036, 
        n31_adj_4249, n29_adj_4250, n29863, n33_adj_4251, n30062, 
        n22971, n22692, n22691, n22690, n22970, n22689, n22969, 
        n22968, n256_adj_4252;
    wire [20:0]n6872;
    
    wire n22967;
    wire [23:0]duty_23__N_3467;
    
    wire n22207, n18_adj_4253, n22966, n22965, n22688, n22964, n22687, 
        n22686, n22206, n22963, n22962, n22685, n22961, n22684, 
        n22960, n22959, n22683, n22958, n22957, n22956, n13_adj_4254, 
        n22955, n22954, n22953, n22952, n4_adj_4255, n22951, n29780, 
        n30952, n29768, n30947, n12_adj_4256, n29510, n30970, n10_adj_4257, 
        n30_adj_4258, n22950, n29961, n22682, n22681, n29518, n22949, 
        n30950, n22948;
    wire [0:0]n5002;
    wire [21:0]n6848;
    
    wire n22947, n29889, n30976, n30040, n22946, n22945, n22944, 
        n22943, n22205, n21945, n22942, n22680, n22679, n22678, 
        n22677, n22676, n22675, n22674, n22673, n22672, n22941, 
        n22940, n22671, n22939, n22938, n22670, n22669, n22937, 
        n22204, n22936, n22668, n22203, n22667, n22666, n22665, 
        n22935, n22664, n22934, n22933, n22932, n22931, n22930, 
        n22663, n22202, n22929, n22928, n22927, n22926, n22925, 
        n22662, n22924, n22923, n22922, n22921, n22920, n22919, 
        n22918, n22917, n30941, n30094, n30938, n16_adj_4263, n29498, 
        n24_adj_4264, n22916, n6_adj_4265, n29909, n22915, n29910, 
        n29500, n22914, n8_adj_4266, n30936, n29865, n22913, n29722, 
        n22912, n22911, n22910, n22909, n22908, n22907, n22906, 
        n22905;
    wire [5:0]n6815;
    
    wire n22904, n22903, n22902, n22901, n22900;
    wire [6:0]n6806;
    
    wire n22899, n22898, n22201, n22897, n22896, n3_adj_4267, n4_adj_4268, 
        n30008, n30009, n12_adj_4269, n29447, n10_adj_4270, n30_adj_4271, 
        n29449, n30068, n29930, n30117, n30118, n30103, n6_adj_4272, 
        n22895, n22894;
    wire [7:0]n6796;
    
    wire n22893, n22892, n22891, n22890, n22889, n22888, n22887;
    wire [8:0]n6785;
    
    wire n22886, n22885, n22884, n22883, n22882, n22881, n22880, 
        n22879;
    wire [9:0]n6773;
    
    wire n22878, n22877, n22876, n22875, n22874, n22873, n22872, 
        n22871, n22870;
    wire [10:0]n6760;
    
    wire n22869, n22868, n22867, n22866, n22865, n22864, n22863, 
        n22862, n29901, n29902, n29439, n29867, n29732, n29441, 
        n30018, n40_adj_4273, n30020, n4_adj_4274, n29907, n29908, 
        n29512, n22861, n22860;
    wire [11:0]n6746;
    
    wire n22859, n22858, n22857, n22200, n22856, n22855, n22854, 
        n22853, n22852, n22851, n22850, n22849;
    wire [12:0]n6731;
    
    wire n22848, n22847, n22846, n22845, n22844, n30052, n29724, 
        n30104, n30105, n30079, n29502, n30014, n29730, \PID_CONTROLLER.integral_23__N_3442 , 
        n30064, n22843, n22842, n22841, n22840, n22839, n22838, 
        n22199, n22837;
    wire [13:0]n6715;
    
    wire n22836, n22835, n22834, n22198, n22197, n22196, n22195, 
        n22194, n22833, n22193, n22192, n22191, n22832, n22831, 
        n22830, n22190, n22829, n22828, n22189, n22188, n22827, 
        n22826, n22825, n22187, n22186, n22824;
    wire [14:0]n6698;
    
    wire n22823, n22822, n22821, n22820, n22819, n22185, n22818, 
        n22817, n22816, n22815, n22814, n22184, n22183, n22182, 
        n22181, n22180, n22179, n22178, n22813, n22812, n22811, 
        n22810;
    wire [15:0]n6680;
    
    wire n22809, n22808, n22807, n22806, n22805, n22804, n22803, 
        n22802, n22801, n22800, n22799, n22798, n22797, n22796, 
        n22795;
    wire [16:0]n6661;
    
    wire n22794, n22793, n22792, n22791, n22790, n22789, n22788, 
        n22787, n22786, n22785, n22177, n22784, n22783, n22782, 
        n22781, n22780, n22779, n22778, n22777, n22776, n22775, 
        n22774, n22773, n22772, n22771, n22770, n22176, n22769, 
        n22175, n22768, n22767, n22766, n22765, n22764, n22763, 
        n22762, n743_adj_4275, n22174, n20_adj_4276, n89_adj_4277, 
        n22761, n22760, n22759, n22758, n1108_adj_4278, n22757, 
        n1035_adj_4279, n22756, n22173, n962_adj_4280, n22755, n816_adj_4281, 
        n889_adj_4282, n22754, n22753, n22172, n22171, n22170, n22752, 
        n21967, n21966, n21965, n22169, n21964, n21954, n21963, 
        n21962, n21961, n22028, n22027, n22026, n21960, n4_adj_4301, 
        n22025, n21959, n670_adj_4302, n21784, n21958, n22024, n22023, 
        n22022, n21861, n21957, n22021, n21956, n22020, n22019, 
        n22018, n22017, n22016, n22237, n21955, n22236, n22235, 
        n22234, n22233, n22232, n22231, n22230, n22229, n22228, 
        n22227, n22226, n22225, n22224, n22223, n22222, n22221, 
        n22015;
    
    SB_CARRY add_3380_9 (.CI(n22750), .I0(n6641[6]), .I1(n597), .CO(n22751));
    SB_LUT4 add_3380_8_lut (.I0(GND_net), .I1(n6641[5]), .I2(n524), .I3(n22749), 
            .O(n6620[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_8 (.CI(n22749), .I0(n6641[5]), .I1(n524), .CO(n22750));
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_10 (.CI(n22013), .I0(n106[8]), .I1(n155[8]), .CO(n22014));
    SB_LUT4 add_3380_7_lut (.I0(GND_net), .I1(n6641[4]), .I2(n451), .I3(n22748), 
            .O(n6620[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3380_7 (.CI(n22748), .I0(n6641[4]), .I1(n451), .CO(n22749));
    SB_CARRY add_560_8 (.CI(n21950), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n2552[6]), .CO(n21951));
    SB_LUT4 add_3380_6_lut (.I0(GND_net), .I1(n6641[3]), .I2(n378), .I3(n22747), 
            .O(n6620[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3380_6 (.CI(n22747), .I0(n6641[3]), .I1(n378), .CO(n22748));
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3380_5_lut (.I0(GND_net), .I1(n6641[2]), .I2(n305), .I3(n22746), 
            .O(n6620[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3380_5 (.CI(n22746), .I0(n6641[2]), .I1(n305), .CO(n22747));
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_560_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n2552[5]), .I3(n21949), .O(\PID_CONTROLLER.integral_23__N_3392 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3380_4_lut (.I0(GND_net), .I1(n6641[1]), .I2(n232), .I3(n22745), 
            .O(n6620[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_4 (.CI(n22745), .I0(n6641[1]), .I1(n232), .CO(n22746));
    SB_LUT4 add_3380_3_lut (.I0(GND_net), .I1(n6641[0]), .I2(n159), .I3(n22744), 
            .O(n6620[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_3 (.CI(n22744), .I0(n6641[0]), .I1(n159), .CO(n22745));
    SB_CARRY unary_minus_16_add_3_7 (.CI(n22219), .I0(GND_net), .I1(n1_adj_4304[5]), 
            .CO(n22220));
    SB_LUT4 add_3380_2_lut (.I0(GND_net), .I1(n17_adj_3887), .I2(n86), 
            .I3(GND_net), .O(n6620[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3380_2 (.CI(GND_net), .I0(n17_adj_3887), .I1(n86), .CO(n22744));
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_21_lut (.I0(GND_net), .I1(n6620[18]), .I2(GND_net), 
            .I3(n22743), .O(n6598[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3415_7_lut (.I0(GND_net), .I1(n27839), .I2(n490), .I3(n23147), 
            .O(n7112[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3415_6_lut (.I0(GND_net), .I1(n7120[3]), .I2(n417), .I3(n23146), 
            .O(n7112[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_6 (.CI(n23146), .I0(n7120[3]), .I1(n417), .CO(n23147));
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_3888));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3415_5_lut (.I0(GND_net), .I1(n7120[2]), .I2(n344), .I3(n23145), 
            .O(n7112[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_5 (.CI(n23145), .I0(n7120[2]), .I1(n344), .CO(n23146));
    SB_LUT4 add_3415_4_lut (.I0(GND_net), .I1(n7120[1]), .I2(n271), .I3(n23144), 
            .O(n7112[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3415_4 (.CI(n23144), .I0(n7120[1]), .I1(n271), .CO(n23145));
    SB_LUT4 add_3415_3_lut (.I0(GND_net), .I1(n7120[0]), .I2(n198), .I3(n23143), 
            .O(n7112[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3415_3 (.CI(n23143), .I0(n7120[0]), .I1(n198), .CO(n23144));
    SB_LUT4 add_3415_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n7112[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n23143));
    SB_LUT4 add_3414_8_lut (.I0(GND_net), .I1(n7112[5]), .I2(n560), .I3(n23142), 
            .O(n7103[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3414_7_lut (.I0(GND_net), .I1(n7112[4]), .I2(n487), .I3(n23141), 
            .O(n7103[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_7 (.CI(n23141), .I0(n7112[4]), .I1(n487), .CO(n23142));
    SB_LUT4 add_3414_6_lut (.I0(GND_net), .I1(n7112[3]), .I2(n414_adj_3889), 
            .I3(n23140), .O(n7103[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_6 (.CI(n23140), .I0(n7112[3]), .I1(n414_adj_3889), 
            .CO(n23141));
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3414_5_lut (.I0(GND_net), .I1(n7112[2]), .I2(n341_adj_3891), 
            .I3(n23139), .O(n7103[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_5 (.CI(n23139), .I0(n7112[2]), .I1(n341_adj_3891), 
            .CO(n23140));
    SB_LUT4 add_3414_4_lut (.I0(GND_net), .I1(n7112[1]), .I2(n268_adj_3892), 
            .I3(n23138), .O(n7103[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_4 (.CI(n23138), .I0(n7112[1]), .I1(n268_adj_3892), 
            .CO(n23139));
    SB_LUT4 add_3414_3_lut (.I0(GND_net), .I1(n7112[0]), .I2(n195_adj_3893), 
            .I3(n23137), .O(n7103[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_3 (.CI(n23137), .I0(n7112[0]), .I1(n195_adj_3893), 
            .CO(n23138));
    SB_LUT4 add_3414_2_lut (.I0(GND_net), .I1(n53_adj_3894), .I2(n122_adj_3895), 
            .I3(GND_net), .O(n7103[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_2 (.CI(GND_net), .I0(n53_adj_3894), .I1(n122_adj_3895), 
            .CO(n23137));
    SB_LUT4 add_3413_9_lut (.I0(GND_net), .I1(n7103[6]), .I2(n630_adj_3896), 
            .I3(n23136), .O(n7093[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3413_8_lut (.I0(GND_net), .I1(n7103[5]), .I2(n557_adj_3897), 
            .I3(n23135), .O(n7093[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_8 (.CI(n23135), .I0(n7103[5]), .I1(n557_adj_3897), 
            .CO(n23136));
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_3898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3413_7_lut (.I0(GND_net), .I1(n7103[4]), .I2(n484_adj_3899), 
            .I3(n23134), .O(n7093[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_7 (.CI(n23134), .I0(n7103[4]), .I1(n484_adj_3899), 
            .CO(n23135));
    SB_LUT4 add_3413_6_lut (.I0(GND_net), .I1(n7103[3]), .I2(n411_adj_3900), 
            .I3(n23133), .O(n7093[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_6 (.CI(n23133), .I0(n7103[3]), .I1(n411_adj_3900), 
            .CO(n23134));
    SB_LUT4 add_3413_5_lut (.I0(GND_net), .I1(n7103[2]), .I2(n338_adj_3901), 
            .I3(n23132), .O(n7093[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_5 (.CI(n23132), .I0(n7103[2]), .I1(n338_adj_3901), 
            .CO(n23133));
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_3902));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3413_4_lut (.I0(GND_net), .I1(n7103[1]), .I2(n265_adj_3903), 
            .I3(n23131), .O(n7093[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_4 (.CI(n23131), .I0(n7103[1]), .I1(n265_adj_3903), 
            .CO(n23132));
    SB_LUT4 add_3413_3_lut (.I0(GND_net), .I1(n7103[0]), .I2(n192_adj_3904), 
            .I3(n23130), .O(n7093[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_3 (.CI(n23130), .I0(n7103[0]), .I1(n192_adj_3904), 
            .CO(n23131));
    SB_LUT4 add_3413_2_lut (.I0(GND_net), .I1(n50_adj_3905), .I2(n119_adj_3906), 
            .I3(GND_net), .O(n7093[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_2 (.CI(GND_net), .I0(n50_adj_3905), .I1(n119_adj_3906), 
            .CO(n23130));
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_3907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3412_10_lut (.I0(GND_net), .I1(n7093[7]), .I2(n700_adj_3908), 
            .I3(n23129), .O(n7082[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3412_9_lut (.I0(GND_net), .I1(n7093[6]), .I2(n627_adj_3909), 
            .I3(n23128), .O(n7082[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_9 (.CI(n23128), .I0(n7093[6]), .I1(n627_adj_3909), 
            .CO(n23129));
    SB_LUT4 add_3412_8_lut (.I0(GND_net), .I1(n7093[5]), .I2(n554_adj_3910), 
            .I3(n23127), .O(n7082[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_8 (.CI(n23127), .I0(n7093[5]), .I1(n554_adj_3910), 
            .CO(n23128));
    SB_LUT4 add_3412_7_lut (.I0(GND_net), .I1(n7093[4]), .I2(n481_adj_3911), 
            .I3(n23126), .O(n7082[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_7 (.CI(n23126), .I0(n7093[4]), .I1(n481_adj_3911), 
            .CO(n23127));
    SB_LUT4 add_3412_6_lut (.I0(GND_net), .I1(n7093[3]), .I2(n408_adj_3912), 
            .I3(n23125), .O(n7082[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_6 (.CI(n23125), .I0(n7093[3]), .I1(n408_adj_3912), 
            .CO(n23126));
    SB_LUT4 add_3412_5_lut (.I0(GND_net), .I1(n7093[2]), .I2(n335_adj_3913), 
            .I3(n23124), .O(n7082[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_5 (.CI(n23124), .I0(n7093[2]), .I1(n335_adj_3913), 
            .CO(n23125));
    SB_LUT4 add_3412_4_lut (.I0(GND_net), .I1(n7093[1]), .I2(n262_adj_3914), 
            .I3(n23123), .O(n7082[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_4 (.CI(n23123), .I0(n7093[1]), .I1(n262_adj_3914), 
            .CO(n23124));
    SB_LUT4 add_3412_3_lut (.I0(GND_net), .I1(n7093[0]), .I2(n189_adj_3915), 
            .I3(n23122), .O(n7082[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_3 (.CI(n23122), .I0(n7093[0]), .I1(n189_adj_3915), 
            .CO(n23123));
    SB_LUT4 add_3412_2_lut (.I0(GND_net), .I1(n47_adj_3916), .I2(n116_adj_3917), 
            .I3(GND_net), .O(n7082[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_2 (.CI(GND_net), .I0(n47_adj_3916), .I1(n116_adj_3917), 
            .CO(n23122));
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_3918));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3411_11_lut (.I0(GND_net), .I1(n7082[8]), .I2(n770_adj_3919), 
            .I3(n23121), .O(n7070[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3411_10_lut (.I0(GND_net), .I1(n7082[7]), .I2(n697_adj_3920), 
            .I3(n23120), .O(n7070[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_3921));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3411_10 (.CI(n23120), .I0(n7082[7]), .I1(n697_adj_3920), 
            .CO(n23121));
    SB_LUT4 add_3411_9_lut (.I0(GND_net), .I1(n7082[6]), .I2(n624_adj_3922), 
            .I3(n23119), .O(n7070[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_9 (.CI(n23119), .I0(n7082[6]), .I1(n624_adj_3922), 
            .CO(n23120));
    SB_LUT4 add_3411_8_lut (.I0(GND_net), .I1(n7082[5]), .I2(n551_adj_3923), 
            .I3(n23118), .O(n7070[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_8 (.CI(n23118), .I0(n7082[5]), .I1(n551_adj_3923), 
            .CO(n23119));
    SB_LUT4 add_3411_7_lut (.I0(GND_net), .I1(n7082[4]), .I2(n478_adj_3924), 
            .I3(n23117), .O(n7070[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_7 (.CI(n23117), .I0(n7082[4]), .I1(n478_adj_3924), 
            .CO(n23118));
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_3925));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3411_6_lut (.I0(GND_net), .I1(n7082[3]), .I2(n405_adj_3926), 
            .I3(n23116), .O(n7070[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_6 (.CI(n23116), .I0(n7082[3]), .I1(n405_adj_3926), 
            .CO(n23117));
    SB_LUT4 add_3411_5_lut (.I0(GND_net), .I1(n7082[2]), .I2(n332_adj_3927), 
            .I3(n23115), .O(n7070[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_5 (.CI(n23115), .I0(n7082[2]), .I1(n332_adj_3927), 
            .CO(n23116));
    SB_LUT4 add_3411_4_lut (.I0(GND_net), .I1(n7082[1]), .I2(n259_adj_3928), 
            .I3(n23114), .O(n7070[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_4 (.CI(n23114), .I0(n7082[1]), .I1(n259_adj_3928), 
            .CO(n23115));
    SB_LUT4 add_3411_3_lut (.I0(GND_net), .I1(n7082[0]), .I2(n186_adj_3929), 
            .I3(n23113), .O(n7070[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_3 (.CI(n23113), .I0(n7082[0]), .I1(n186_adj_3929), 
            .CO(n23114));
    SB_LUT4 add_3411_2_lut (.I0(GND_net), .I1(n44_adj_3930), .I2(n113_adj_3931), 
            .I3(GND_net), .O(n7070[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_2 (.CI(GND_net), .I0(n44_adj_3930), .I1(n113_adj_3931), 
            .CO(n23113));
    SB_LUT4 add_3410_12_lut (.I0(GND_net), .I1(n7070[9]), .I2(n840_adj_3932), 
            .I3(n23112), .O(n7057[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3410_11_lut (.I0(GND_net), .I1(n7070[8]), .I2(n767_adj_3933), 
            .I3(n23111), .O(n7057[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_11 (.CI(n23111), .I0(n7070[8]), .I1(n767_adj_3933), 
            .CO(n23112));
    SB_LUT4 add_3410_10_lut (.I0(GND_net), .I1(n7070[7]), .I2(n694_adj_3934), 
            .I3(n23110), .O(n7057[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_10 (.CI(n23110), .I0(n7070[7]), .I1(n694_adj_3934), 
            .CO(n23111));
    SB_LUT4 add_3410_9_lut (.I0(GND_net), .I1(n7070[6]), .I2(n621_adj_3935), 
            .I3(n23109), .O(n7057[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_9 (.CI(n23109), .I0(n7070[6]), .I1(n621_adj_3935), 
            .CO(n23110));
    SB_LUT4 add_3410_8_lut (.I0(GND_net), .I1(n7070[5]), .I2(n548_adj_3936), 
            .I3(n23108), .O(n7057[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_8 (.CI(n23108), .I0(n7070[5]), .I1(n548_adj_3936), 
            .CO(n23109));
    SB_LUT4 add_3410_7_lut (.I0(GND_net), .I1(n7070[4]), .I2(n475_adj_3937), 
            .I3(n23107), .O(n7057[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_7 (.CI(n23107), .I0(n7070[4]), .I1(n475_adj_3937), 
            .CO(n23108));
    SB_LUT4 add_3410_6_lut (.I0(GND_net), .I1(n7070[3]), .I2(n402_adj_3938), 
            .I3(n23106), .O(n7057[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_6 (.CI(n23106), .I0(n7070[3]), .I1(n402_adj_3938), 
            .CO(n23107));
    SB_LUT4 add_3410_5_lut (.I0(GND_net), .I1(n7070[2]), .I2(n329_adj_3939), 
            .I3(n23105), .O(n7057[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_5 (.CI(n23105), .I0(n7070[2]), .I1(n329_adj_3939), 
            .CO(n23106));
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_3940));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3410_4_lut (.I0(GND_net), .I1(n7070[1]), .I2(n256_adj_3941), 
            .I3(n23104), .O(n7057[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_4 (.CI(n23104), .I0(n7070[1]), .I1(n256_adj_3941), 
            .CO(n23105));
    SB_LUT4 add_3410_3_lut (.I0(GND_net), .I1(n7070[0]), .I2(n183_adj_3942), 
            .I3(n23103), .O(n7057[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_3 (.CI(n23103), .I0(n7070[0]), .I1(n183_adj_3942), 
            .CO(n23104));
    SB_LUT4 add_3410_2_lut (.I0(GND_net), .I1(n41_adj_3943), .I2(n110_adj_3944), 
            .I3(GND_net), .O(n7057[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_2 (.CI(GND_net), .I0(n41_adj_3943), .I1(n110_adj_3944), 
            .CO(n23103));
    SB_LUT4 add_3409_13_lut (.I0(GND_net), .I1(n7057[10]), .I2(n910_adj_3945), 
            .I3(n23102), .O(n7043[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3409_12_lut (.I0(GND_net), .I1(n7057[9]), .I2(n837_adj_3946), 
            .I3(n23101), .O(n7043[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_12 (.CI(n23101), .I0(n7057[9]), .I1(n837_adj_3946), 
            .CO(n23102));
    SB_LUT4 add_3409_11_lut (.I0(GND_net), .I1(n7057[8]), .I2(n764_adj_3947), 
            .I3(n23100), .O(n7043[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_11 (.CI(n23100), .I0(n7057[8]), .I1(n764_adj_3947), 
            .CO(n23101));
    SB_LUT4 add_3409_10_lut (.I0(GND_net), .I1(n7057[7]), .I2(n691_adj_3948), 
            .I3(n23099), .O(n7043[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_10 (.CI(n23099), .I0(n7057[7]), .I1(n691_adj_3948), 
            .CO(n23100));
    SB_LUT4 add_3409_9_lut (.I0(GND_net), .I1(n7057[6]), .I2(n618_adj_3949), 
            .I3(n23098), .O(n7043[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_9 (.CI(n23098), .I0(n7057[6]), .I1(n618_adj_3949), 
            .CO(n23099));
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3409_8_lut (.I0(GND_net), .I1(n7057[5]), .I2(n545_adj_3950), 
            .I3(n23097), .O(n7043[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_8 (.CI(n23097), .I0(n7057[5]), .I1(n545_adj_3950), 
            .CO(n23098));
    SB_LUT4 add_3409_7_lut (.I0(GND_net), .I1(n7057[4]), .I2(n472_adj_3951), 
            .I3(n23096), .O(n7043[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3409_7 (.CI(n23096), .I0(n7057[4]), .I1(n472_adj_3951), 
            .CO(n23097));
    SB_LUT4 add_3409_6_lut (.I0(GND_net), .I1(n7057[3]), .I2(n399_adj_3952), 
            .I3(n23095), .O(n7043[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_6 (.CI(n23095), .I0(n7057[3]), .I1(n399_adj_3952), 
            .CO(n23096));
    SB_LUT4 add_3409_5_lut (.I0(GND_net), .I1(n7057[2]), .I2(n326_adj_3953), 
            .I3(n23094), .O(n7043[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_5 (.CI(n23094), .I0(n7057[2]), .I1(n326_adj_3953), 
            .CO(n23095));
    SB_LUT4 add_3409_4_lut (.I0(GND_net), .I1(n7057[1]), .I2(n253_adj_3954), 
            .I3(n23093), .O(n7043[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_4 (.CI(n23093), .I0(n7057[1]), .I1(n253_adj_3954), 
            .CO(n23094));
    SB_LUT4 add_3409_3_lut (.I0(GND_net), .I1(n7057[0]), .I2(n180_adj_3955), 
            .I3(n23092), .O(n7043[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_3 (.CI(n23092), .I0(n7057[0]), .I1(n180_adj_3955), 
            .CO(n23093));
    SB_LUT4 add_3409_2_lut (.I0(GND_net), .I1(n38_adj_3956), .I2(n107_adj_3957), 
            .I3(GND_net), .O(n7043[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_2 (.CI(GND_net), .I0(n38_adj_3956), .I1(n107_adj_3957), 
            .CO(n23092));
    SB_LUT4 add_3408_14_lut (.I0(GND_net), .I1(n7043[11]), .I2(n980_adj_3958), 
            .I3(n23091), .O(n7028[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3408_13_lut (.I0(GND_net), .I1(n7043[10]), .I2(n907_adj_3959), 
            .I3(n23090), .O(n7028[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_3960));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3408_13 (.CI(n23090), .I0(n7043[10]), .I1(n907_adj_3959), 
            .CO(n23091));
    SB_LUT4 i2_4_lut (.I0(n6), .I1(\Kp[4] ), .I2(n6830[2]), .I3(n1[18]), 
            .O(n6823[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 add_3408_12_lut (.I0(GND_net), .I1(n7043[9]), .I2(n834_adj_3961), 
            .I3(n23089), .O(n7028[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_12 (.CI(n23089), .I0(n7043[9]), .I1(n834_adj_3961), 
            .CO(n23090));
    SB_LUT4 add_3408_11_lut (.I0(GND_net), .I1(n7043[8]), .I2(n761_adj_3962), 
            .I3(n23088), .O(n7028[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_11 (.CI(n23088), .I0(n7043[8]), .I1(n761_adj_3962), 
            .CO(n23089));
    SB_LUT4 add_3408_10_lut (.I0(GND_net), .I1(n7043[7]), .I2(n688_adj_3963), 
            .I3(n23087), .O(n7028[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_10 (.CI(n23087), .I0(n7043[7]), .I1(n688_adj_3963), 
            .CO(n23088));
    SB_LUT4 add_3408_9_lut (.I0(GND_net), .I1(n7043[6]), .I2(n615_adj_3964), 
            .I3(n23086), .O(n7028[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_9 (.CI(n23086), .I0(n7043[6]), .I1(n615_adj_3964), 
            .CO(n23087));
    SB_LUT4 add_3408_8_lut (.I0(GND_net), .I1(n7043[5]), .I2(n542_adj_3965), 
            .I3(n23085), .O(n7028[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_8 (.CI(n23085), .I0(n7043[5]), .I1(n542_adj_3965), 
            .CO(n23086));
    SB_LUT4 add_3408_7_lut (.I0(GND_net), .I1(n7043[4]), .I2(n469_adj_3966), 
            .I3(n23084), .O(n7028[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_7 (.CI(n23084), .I0(n7043[4]), .I1(n469_adj_3966), 
            .CO(n23085));
    SB_LUT4 add_3408_6_lut (.I0(GND_net), .I1(n7043[3]), .I2(n396_adj_3967), 
            .I3(n23083), .O(n7028[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_6 (.CI(n23083), .I0(n7043[3]), .I1(n396_adj_3967), 
            .CO(n23084));
    SB_LUT4 add_3408_5_lut (.I0(GND_net), .I1(n7043[2]), .I2(n323_adj_3968), 
            .I3(n23082), .O(n7028[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_5 (.CI(n23082), .I0(n7043[2]), .I1(n323_adj_3968), 
            .CO(n23083));
    SB_LUT4 add_3408_4_lut (.I0(GND_net), .I1(n7043[1]), .I2(n250_adj_3969), 
            .I3(n23081), .O(n7028[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_4 (.CI(n23081), .I0(n7043[1]), .I1(n250_adj_3969), 
            .CO(n23082));
    SB_LUT4 add_3408_3_lut (.I0(GND_net), .I1(n7043[0]), .I2(n177_adj_3970), 
            .I3(n23080), .O(n7028[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_3 (.CI(n23080), .I0(n7043[0]), .I1(n177_adj_3970), 
            .CO(n23081));
    SB_LUT4 add_3408_2_lut (.I0(GND_net), .I1(n35_adj_3971), .I2(n104_adj_3972), 
            .I3(GND_net), .O(n7028[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_2 (.CI(GND_net), .I0(n35_adj_3971), .I1(n104_adj_3972), 
            .CO(n23080));
    SB_LUT4 add_3407_15_lut (.I0(GND_net), .I1(n7028[12]), .I2(n1050_adj_3973), 
            .I3(n23079), .O(n7012[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_14_lut (.I0(GND_net), .I1(n7028[11]), .I2(n977_adj_3974), 
            .I3(n23078), .O(n7012[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_14 (.CI(n23078), .I0(n7028[11]), .I1(n977_adj_3974), 
            .CO(n23079));
    SB_LUT4 add_3407_13_lut (.I0(GND_net), .I1(n7028[10]), .I2(n904_adj_3975), 
            .I3(n23077), .O(n7012[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_13 (.CI(n23077), .I0(n7028[10]), .I1(n904_adj_3975), 
            .CO(n23078));
    SB_LUT4 add_3407_12_lut (.I0(GND_net), .I1(n7028[9]), .I2(n831_adj_3976), 
            .I3(n23076), .O(n7012[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_12 (.CI(n23076), .I0(n7028[9]), .I1(n831_adj_3976), 
            .CO(n23077));
    SB_LUT4 add_3407_11_lut (.I0(GND_net), .I1(n7028[8]), .I2(n758_adj_3977), 
            .I3(n23075), .O(n7012[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_11 (.CI(n23075), .I0(n7028[8]), .I1(n758_adj_3977), 
            .CO(n23076));
    SB_LUT4 add_3407_10_lut (.I0(GND_net), .I1(n7028[7]), .I2(n685_adj_3978), 
            .I3(n23074), .O(n7012[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_10 (.CI(n23074), .I0(n7028[7]), .I1(n685_adj_3978), 
            .CO(n23075));
    SB_LUT4 add_3407_9_lut (.I0(GND_net), .I1(n7028[6]), .I2(n612_adj_3979), 
            .I3(n23073), .O(n7012[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_9 (.CI(n23073), .I0(n7028[6]), .I1(n612_adj_3979), 
            .CO(n23074));
    SB_LUT4 add_3407_8_lut (.I0(GND_net), .I1(n7028[5]), .I2(n539_adj_3980), 
            .I3(n23072), .O(n7012[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_8 (.CI(n23072), .I0(n7028[5]), .I1(n539_adj_3980), 
            .CO(n23073));
    SB_LUT4 add_3407_7_lut (.I0(GND_net), .I1(n7028[4]), .I2(n466_adj_3981), 
            .I3(n23071), .O(n7012[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_7 (.CI(n23071), .I0(n7028[4]), .I1(n466_adj_3981), 
            .CO(n23072));
    SB_LUT4 add_3407_6_lut (.I0(GND_net), .I1(n7028[3]), .I2(n393_adj_3982), 
            .I3(n23070), .O(n7012[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_6 (.CI(n23070), .I0(n7028[3]), .I1(n393_adj_3982), 
            .CO(n23071));
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3887));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_5_lut (.I0(GND_net), .I1(n7028[2]), .I2(n320_adj_3983), 
            .I3(n23069), .O(n7012[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3379_20_lut (.I0(GND_net), .I1(n6620[17]), .I2(GND_net), 
            .I3(n22742), .O(n6598[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3407_5 (.CI(n23069), .I0(n7028[2]), .I1(n320_adj_3983), 
            .CO(n23070));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n22012), 
            .O(duty_23__N_3492[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1439 (.I0(n4), .I1(\Kp[3] ), .I2(n6836[1]), .I3(n1[19]), 
            .O(n6830[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1439.LUT_INIT = 16'h965a;
    SB_LUT4 i17965_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n6841[0]));   // verilog/motorControl.v(34[16:22])
    defparam i17965_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_4_lut (.I0(GND_net), .I1(n7028[1]), .I2(n247_adj_3985), 
            .I3(n23068), .O(n7012[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_4 (.CI(n23068), .I0(n7028[1]), .I1(n247_adj_3985), 
            .CO(n23069));
    SB_LUT4 add_3407_3_lut (.I0(GND_net), .I1(n7028[0]), .I2(n174_adj_3986), 
            .I3(n23067), .O(n7012[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_3 (.CI(n23067), .I0(n7028[0]), .I1(n174_adj_3986), 
            .CO(n23068));
    SB_CARRY add_3379_20 (.CI(n22742), .I0(n6620[17]), .I1(GND_net), .CO(n22743));
    SB_LUT4 add_3407_2_lut (.I0(GND_net), .I1(n32_adj_3987), .I2(n101_adj_3988), 
            .I3(GND_net), .O(n7012[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[4]), 
            .I3(n22218), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3379_19_lut (.I0(GND_net), .I1(n6620[16]), .I2(GND_net), 
            .I3(n22741), .O(n6598[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_19 (.CI(n22741), .I0(n6620[16]), .I1(GND_net), .CO(n22742));
    SB_CARRY add_3407_2 (.CI(GND_net), .I0(n32_adj_3987), .I1(n101_adj_3988), 
            .CO(n23067));
    SB_LUT4 add_3379_18_lut (.I0(GND_net), .I1(n6620[15]), .I2(GND_net), 
            .I3(n22740), .O(n6598[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3406_16_lut (.I0(GND_net), .I1(n7012[13]), .I2(n1120_adj_3990), 
            .I3(n23066), .O(n6995[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_18 (.CI(n22740), .I0(n6620[15]), .I1(GND_net), .CO(n22741));
    SB_LUT4 add_3379_17_lut (.I0(GND_net), .I1(n6620[14]), .I2(GND_net), 
            .I3(n22739), .O(n6598[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_7 (.CI(n21949), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n2552[5]), .CO(n21950));
    SB_CARRY add_3379_17 (.CI(n22739), .I0(n6620[14]), .I1(GND_net), .CO(n22740));
    SB_LUT4 add_3406_15_lut (.I0(GND_net), .I1(n7012[12]), .I2(n1047_adj_3991), 
            .I3(n23065), .O(n6995[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3379_16_lut (.I0(GND_net), .I1(n6620[13]), .I2(n1105), 
            .I3(n22738), .O(n6598[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n22218), .I0(GND_net), .I1(n1_adj_4304[4]), 
            .CO(n22219));
    SB_CARRY add_3406_15 (.CI(n23065), .I0(n7012[12]), .I1(n1047_adj_3991), 
            .CO(n23066));
    SB_CARRY add_3379_16 (.CI(n22738), .I0(n6620[13]), .I1(n1105), .CO(n22739));
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_3992));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1440 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_3994));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1440.LUT_INIT = 16'h9c50;
    SB_LUT4 i17901_4_lut (.I0(n6830[2]), .I1(\Kp[4] ), .I2(n6), .I3(n1[18]), 
            .O(n8_adj_3995));   // verilog/motorControl.v(34[16:22])
    defparam i17901_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[3]), 
            .I3(n22217), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n22012), .I0(n106[7]), .I1(n155[7]), .CO(n22013));
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), .I3(n1[21]), 
            .O(n11_adj_3997));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i17932_4_lut (.I0(n6836[1]), .I1(\Kp[3] ), .I2(n4), .I3(n1[19]), 
            .O(n6_adj_3998));   // verilog/motorControl.v(34[16:22])
    defparam i17932_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i17967_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n21754));   // verilog/motorControl.v(34[16:22])
    defparam i17967_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_3998), .I1(n11_adj_3997), .I2(n8_adj_3995), 
            .I3(n12_adj_3994), .O(n18_adj_3999));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), .I3(n1[22]), 
            .O(n13_adj_4000));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4000), .I1(n18_adj_3999), .I2(n21754), 
            .I3(n4_adj_4001), .O(n27634));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3379_15_lut (.I0(GND_net), .I1(n6620[12]), .I2(n1032), 
            .I3(n22737), .O(n6598[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_15 (.CI(n22737), .I0(n6620[12]), .I1(n1032), .CO(n22738));
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4002));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_14_lut (.I0(GND_net), .I1(n6620[11]), .I2(n959), 
            .I3(n22736), .O(n6598[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3379_14 (.CI(n22736), .I0(n6620[11]), .I1(n959), .CO(n22737));
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3406_14_lut (.I0(GND_net), .I1(n7012[11]), .I2(n974_adj_4003), 
            .I3(n23064), .O(n6995[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_14 (.CI(n23064), .I0(n7012[11]), .I1(n974_adj_4003), 
            .CO(n23065));
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4005));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4007));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4008));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4009));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_13_lut (.I0(GND_net), .I1(n6620[10]), .I2(n886), 
            .I3(n22735), .O(n6598[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4010));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n22217), .I0(GND_net), .I1(n1_adj_4304[3]), 
            .CO(n22218));
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4012));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4013));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3406_13_lut (.I0(GND_net), .I1(n7012[10]), .I2(n901_adj_4014), 
            .I3(n23063), .O(n6995[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_13 (.CI(n22735), .I0(n6620[10]), .I1(n886), .CO(n22736));
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4015));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4016));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4017));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14954_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i14954_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3379_12_lut (.I0(GND_net), .I1(n6620[9]), .I2(n813), .I3(n22734), 
            .O(n6598[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4019));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4021));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4022));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3379_12 (.CI(n22734), .I0(n6620[9]), .I1(n813), .CO(n22735));
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4024));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4025));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4027));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15182_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15182_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4030));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_13 (.CI(n23063), .I0(n7012[10]), .I1(n901_adj_4014), 
            .CO(n23064));
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4031));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_11_lut (.I0(GND_net), .I1(n6620[8]), .I2(n740), .I3(n22733), 
            .O(n6598[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_11 (.CI(n22733), .I0(n6620[8]), .I1(n740), .CO(n22734));
    SB_LUT4 add_3379_10_lut (.I0(GND_net), .I1(n6620[7]), .I2(n667), .I3(n22732), 
            .O(n6598[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_10 (.CI(n22732), .I0(n6620[7]), .I1(n667), .CO(n22733));
    SB_LUT4 i25197_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30261));   // verilog/motorControl.v(29[14] 48[8])
    defparam i25197_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4033));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4034));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4036));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4037));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4040));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4042));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4043));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4045));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4046));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4048));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4049));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4051));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4053));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[2]), 
            .I3(n22216), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4055));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4056));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4057));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4059));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4060));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4061));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4062));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4064));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4065));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4066));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4067));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4068));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4069));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4070));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3406_12_lut (.I0(GND_net), .I1(n7012[9]), .I2(n828_adj_4071), 
            .I3(n23062), .O(n6995[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4072));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4073));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15188_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15188_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4075));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4076));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4077));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4078));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4079));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4080));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4081));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4082));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4083));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4084));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4085));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4086));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4087));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4088));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4089));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_3900));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4090));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_9_lut (.I0(GND_net), .I1(n6620[6]), .I2(n594_adj_4091), 
            .I3(n22731), .O(n6598[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_9 (.CI(n22731), .I0(n6620[6]), .I1(n594_adj_4091), 
            .CO(n22732));
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4092));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4093));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4094));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3379_8_lut (.I0(GND_net), .I1(n6620[5]), .I2(n521_adj_4095), 
            .I3(n22730), .O(n6598[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_3899));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4097));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4100));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15183_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4101));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_12 (.CI(n23062), .I0(n7012[9]), .I1(n828_adj_4071), 
            .CO(n23063));
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24471_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n29535));
    defparam i24471_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4103));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3406_11_lut (.I0(GND_net), .I1(n7012[8]), .I2(n755_adj_4105), 
            .I3(n23061), .O(n6995[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_8 (.CI(n22730), .I0(n6620[5]), .I1(n521_adj_4095), 
            .CO(n22731));
    SB_CARRY add_3406_11 (.CI(n23061), .I0(n7012[8]), .I1(n755_adj_4105), 
            .CO(n23062));
    SB_LUT4 add_3406_10_lut (.I0(GND_net), .I1(n7012[7]), .I2(n682_adj_4106), 
            .I3(n23060), .O(n6995[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_10 (.CI(n23060), .I0(n7012[7]), .I1(n682_adj_4106), 
            .CO(n23061));
    SB_LUT4 add_3379_7_lut (.I0(GND_net), .I1(n6620[4]), .I2(n448_adj_4107), 
            .I3(n22729), .O(n6598[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_7 (.CI(n22729), .I0(n6620[4]), .I1(n448_adj_4107), 
            .CO(n22730));
    SB_LUT4 add_3406_9_lut (.I0(GND_net), .I1(n7012[6]), .I2(n609_adj_4108), 
            .I3(n23059), .O(n6995[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_3897));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_9 (.CI(n23059), .I0(n7012[6]), .I1(n609_adj_4108), 
            .CO(n23060));
    SB_LUT4 add_3379_6_lut (.I0(GND_net), .I1(n6620[3]), .I2(n375_adj_4109), 
            .I3(n22728), .O(n6598[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_6 (.CI(n22728), .I0(n6620[3]), .I1(n375_adj_4109), 
            .CO(n22729));
    SB_LUT4 add_3406_8_lut (.I0(GND_net), .I1(n7012[5]), .I2(n536_adj_4110), 
            .I3(n23058), .O(n6995[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_8 (.CI(n23058), .I0(n7012[5]), .I1(n536_adj_4110), 
            .CO(n23059));
    SB_LUT4 add_3406_7_lut (.I0(GND_net), .I1(n7012[4]), .I2(n463_adj_4111), 
            .I3(n23057), .O(n6995[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_7 (.CI(n23057), .I0(n7012[4]), .I1(n463_adj_4111), 
            .CO(n23058));
    SB_LUT4 add_3406_6_lut (.I0(GND_net), .I1(n7012[3]), .I2(n390), .I3(n23056), 
            .O(n6995[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_6 (.CI(n23056), .I0(n7012[3]), .I1(n390), .CO(n23057));
    SB_LUT4 add_3406_5_lut (.I0(GND_net), .I1(n7012[2]), .I2(n317), .I3(n23055), 
            .O(n6995[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_5 (.CI(n23055), .I0(n7012[2]), .I1(n317), .CO(n23056));
    SB_LUT4 add_3379_5_lut (.I0(GND_net), .I1(n6620[2]), .I2(n302_adj_4112), 
            .I3(n22727), .O(n6598[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_5 (.CI(n22727), .I0(n6620[2]), .I1(n302_adj_4112), 
            .CO(n22728));
    SB_LUT4 add_3406_4_lut (.I0(GND_net), .I1(n7012[1]), .I2(n244), .I3(n23054), 
            .O(n6995[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_4 (.CI(n23054), .I0(n7012[1]), .I1(n244), .CO(n23055));
    SB_LUT4 add_3406_3_lut (.I0(GND_net), .I1(n7012[0]), .I2(n171), .I3(n23053), 
            .O(n6995[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_3 (.CI(n23053), .I0(n7012[0]), .I1(n171), .CO(n23054));
    SB_LUT4 add_3406_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n6995[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3379_4_lut (.I0(GND_net), .I1(n6620[1]), .I2(n229_adj_4113), 
            .I3(n22726), .O(n6598[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n22216), .I0(GND_net), .I1(n1_adj_4304[2]), 
            .CO(n22217));
    SB_CARRY add_3406_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n23053));
    SB_LUT4 add_3405_17_lut (.I0(GND_net), .I1(n6995[14]), .I2(GND_net), 
            .I3(n23052), .O(n6977[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_4 (.CI(n22726), .I0(n6620[1]), .I1(n229_adj_4113), 
            .CO(n22727));
    SB_LUT4 add_3379_3_lut (.I0(GND_net), .I1(n6620[0]), .I2(n156_adj_4114), 
            .I3(n22725), .O(n6598[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3405_16_lut (.I0(GND_net), .I1(n6995[13]), .I2(n1117), 
            .I3(n23051), .O(n6977[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_16 (.CI(n23051), .I0(n6995[13]), .I1(n1117), .CO(n23052));
    SB_CARRY add_3379_3 (.CI(n22725), .I0(n6620[0]), .I1(n156_adj_4114), 
            .CO(n22726));
    SB_LUT4 add_3379_2_lut (.I0(GND_net), .I1(n14_adj_4115), .I2(n83_adj_4116), 
            .I3(GND_net), .O(n6598[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3379_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_3896));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3405_15_lut (.I0(GND_net), .I1(n6995[12]), .I2(n1044), 
            .I3(n23050), .O(n6977[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_15 (.CI(n23050), .I0(n6995[12]), .I1(n1044), .CO(n23051));
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3405_14_lut (.I0(GND_net), .I1(n6995[11]), .I2(n971), 
            .I3(n23049), .O(n6977[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3405_14 (.CI(n23049), .I0(n6995[11]), .I1(n971), .CO(n23050));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[1]), 
            .I3(n22215), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n22215), .I0(GND_net), .I1(n1_adj_4304[1]), 
            .CO(n22216));
    SB_LUT4 add_3405_13_lut (.I0(GND_net), .I1(n6995[10]), .I2(n898), 
            .I3(n23048), .O(n6977[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_13 (.CI(n23048), .I0(n6995[10]), .I1(n898), .CO(n23049));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3405_12_lut (.I0(GND_net), .I1(n6995[9]), .I2(n825), .I3(n23047), 
            .O(n6977[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3379_2 (.CI(GND_net), .I0(n14_adj_4115), .I1(n83_adj_4116), 
            .CO(n22725));
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4304[0]), 
            .CO(n22215));
    SB_CARRY add_3405_12 (.CI(n23047), .I0(n6995[9]), .I1(n825), .CO(n23048));
    SB_LUT4 add_3405_11_lut (.I0(GND_net), .I1(n6995[8]), .I2(n752), .I3(n23046), 
            .O(n6977[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_11 (.CI(n23046), .I0(n6995[8]), .I1(n752), .CO(n23047));
    SB_LUT4 add_3405_10_lut (.I0(GND_net), .I1(n6995[7]), .I2(n679), .I3(n23045), 
            .O(n6977[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3894));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3378_22_lut (.I0(GND_net), .I1(n6598[19]), .I2(GND_net), 
            .I3(n22724), .O(n6575[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4120));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3893));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4121));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3405_10 (.CI(n23045), .I0(n6995[7]), .I1(n679), .CO(n23046));
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_3891));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_3889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4123));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4124));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3378_21_lut (.I0(GND_net), .I1(n6598[18]), .I2(GND_net), 
            .I3(n22723), .O(n6575[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3378_21 (.CI(n22723), .I0(n6598[18]), .I1(GND_net), .CO(n22724));
    SB_LUT4 add_3378_20_lut (.I0(GND_net), .I1(n6598[17]), .I2(GND_net), 
            .I3(n22722), .O(n6575[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_20 (.CI(n22722), .I0(n6598[17]), .I1(GND_net), .CO(n22723));
    SB_LUT4 add_3405_9_lut (.I0(GND_net), .I1(n6995[6]), .I2(n606_adj_4126), 
            .I3(n23044), .O(n6977[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4127));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4128));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n22011), 
            .O(duty_23__N_3492[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4129));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4130));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3378_19_lut (.I0(GND_net), .I1(n6598[16]), .I2(GND_net), 
            .I3(n22721), .O(n6575[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4131));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4132));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4133));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_8 (.CI(n22011), .I0(n106[6]), .I1(n155[6]), .CO(n22012));
    SB_CARRY add_3378_19 (.CI(n22721), .I0(n6598[16]), .I1(GND_net), .CO(n22722));
    SB_LUT4 add_3378_18_lut (.I0(GND_net), .I1(n6598[15]), .I2(GND_net), 
            .I3(n22720), .O(n6575[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4134));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3378_18 (.CI(n22720), .I0(n6598[15]), .I1(GND_net), .CO(n22721));
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4135));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4136));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4137));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3405_9 (.CI(n23044), .I0(n6995[6]), .I1(n606_adj_4126), 
            .CO(n23045));
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4138));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1441 (.I0(n6_adj_4139), .I1(\Ki[4] ), .I2(n7127[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [18]), .O(n7120[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1441.LUT_INIT = 16'h965a;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n22010), 
            .O(duty_23__N_3492[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4141));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4142));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4143));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4144));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24468_3_lut (.I0(n11_adj_4145), .I1(n9_adj_4146), .I2(n29535), 
            .I3(GND_net), .O(n29532));
    defparam i24468_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18087_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3392 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [21]), .O(n7138[0]));   // verilog/motorControl.v(34[25:36])
    defparam i18087_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_3405_8_lut (.I0(GND_net), .I1(n6995[5]), .I2(n533_adj_4148), 
            .I3(n23043), .O(n6977[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4149));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3405_8 (.CI(n23043), .I0(n6995[5]), .I1(n533_adj_4148), 
            .CO(n23044));
    SB_LUT4 add_560_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n2552[8]), .I3(n21952), .O(\PID_CONTROLLER.integral_23__N_3392 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n2552[4]), .I3(n21948), .O(\PID_CONTROLLER.integral_23__N_3392 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17924_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n21695), 
            .I3(n6836[0]), .O(n4));   // verilog/motorControl.v(34[16:22])
    defparam i17924_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n6836[0]), 
            .I3(n21695), .O(n6830[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17955_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n21729), 
            .I3(n6841[0]), .O(n4_adj_4001));   // verilog/motorControl.v(34[16:22])
    defparam i17955_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4151));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4152));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1442 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n6841[0]), 
            .I3(n21729), .O(n6836[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1442.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_831_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3492[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4154));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3492[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3405_7_lut (.I0(GND_net), .I1(n6995[4]), .I2(n460_adj_4155), 
            .I3(n23042), .O(n6977[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3492[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17944_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n21729));   // verilog/motorControl.v(34[16:22])
    defparam i17944_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 duty_23__I_831_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3492[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3378_17_lut (.I0(GND_net), .I1(n6598[14]), .I2(GND_net), 
            .I3(n22719), .O(n6575[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n22010), .I0(n106[5]), .I1(n155[5]), .CO(n22011));
    SB_LUT4 duty_23__I_831_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3492[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4156));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17942_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n6836[0]));   // verilog/motorControl.v(34[16:22])
    defparam i17942_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 duty_23__I_831_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3492[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_64_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n30983));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_64_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3378_17 (.CI(n22719), .I0(n6598[14]), .I1(GND_net), .CO(n22720));
    SB_LUT4 add_3378_16_lut (.I0(GND_net), .I1(n6598[13]), .I2(n1102_adj_4157), 
            .I3(n22718), .O(n6575[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3492[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3492[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4158));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3492[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4159));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15196_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15196_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_831_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3492[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4160));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3492[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4161));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24829_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n30983), 
            .I2(IntegralLimit[7]), .I3(n29532), .O(n29895));
    defparam i24829_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_3378_16 (.CI(n22718), .I0(n6598[13]), .I1(n1102_adj_4157), 
            .CO(n22719));
    SB_LUT4 i24712_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4162), 
            .I2(IntegralLimit[9]), .I3(n29895), .O(n29778));
    defparam i24712_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_3405_7 (.CI(n23042), .I0(n6995[4]), .I1(n460_adj_4155), 
            .CO(n23043));
    SB_LUT4 add_3378_15_lut (.I0(GND_net), .I1(n6598[12]), .I2(n1029_adj_4163), 
            .I3(n22717), .O(n6575[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_10 (.CI(n21952), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n2552[8]), .CO(n21953));
    SB_LUT4 duty_23__I_831_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3492[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4164));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3405_6_lut (.I0(GND_net), .I1(n6995[3]), .I2(n387_adj_4165), 
            .I3(n23041), .O(n6977[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4166));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3378_15 (.CI(n22717), .I0(n6598[12]), .I1(n1029_adj_4163), 
            .CO(n22718));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n22009), 
            .O(duty_23__N_3492[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3378_14_lut (.I0(GND_net), .I1(n6598[11]), .I2(n956_adj_4168), 
            .I3(n22716), .O(n6575[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_6 (.CI(n23041), .I0(n6995[3]), .I1(n387_adj_4165), 
            .CO(n23042));
    SB_LUT4 add_3405_5_lut (.I0(GND_net), .I1(n6995[2]), .I2(n314_adj_4169), 
            .I3(n23040), .O(n6977[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_14 (.CI(n22716), .I0(n6598[11]), .I1(n956_adj_4168), 
            .CO(n22717));
    SB_CARRY add_3405_5 (.CI(n23040), .I0(n6995[2]), .I1(n314_adj_4169), 
            .CO(n23041));
    SB_LUT4 duty_23__I_831_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3492[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4170));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3492[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3492[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3492[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4171));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_560_6 (.CI(n21948), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n2552[4]), .CO(n21949));
    SB_LUT4 duty_23__I_831_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3492[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4172));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3378_13_lut (.I0(GND_net), .I1(n6598[10]), .I2(n883_adj_4173), 
            .I3(n22715), .O(n6575[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3492[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4174));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3405_4_lut (.I0(GND_net), .I1(n6995[1]), .I2(n241_adj_4175), 
            .I3(n23039), .O(n6977[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_13 (.CI(n22715), .I0(n6598[10]), .I1(n883_adj_4173), 
            .CO(n22716));
    SB_CARRY add_3405_4 (.CI(n23039), .I0(n6995[1]), .I1(n241_adj_4175), 
            .CO(n23040));
    SB_CARRY add_12_6 (.CI(n22009), .I0(n106[4]), .I1(n155[4]), .CO(n22010));
    SB_LUT4 add_3405_3_lut (.I0(GND_net), .I1(n6995[0]), .I2(n168_adj_4176), 
            .I3(n23038), .O(n6977[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_3 (.CI(n23038), .I0(n6995[0]), .I1(n168_adj_4176), 
            .CO(n23039));
    SB_LUT4 add_560_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n2552[3]), .I3(n21947), .O(\PID_CONTROLLER.integral_23__N_3392 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3405_2_lut (.I0(GND_net), .I1(n26_adj_4177), .I2(n95_adj_4178), 
            .I3(GND_net), .O(n6977[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3405_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4303[23]), 
            .I3(n22214), .O(\PID_CONTROLLER.integral_23__N_3443 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3378_12_lut (.I0(GND_net), .I1(n6598[9]), .I2(n810_adj_4179), 
            .I3(n22714), .O(n6575[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3405_2 (.CI(GND_net), .I0(n26_adj_4177), .I1(n95_adj_4178), 
            .CO(n23038));
    SB_LUT4 add_3404_18_lut (.I0(GND_net), .I1(n6977[15]), .I2(GND_net), 
            .I3(n23037), .O(n6958[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3492[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4180));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3404_17_lut (.I0(GND_net), .I1(n6977[14]), .I2(GND_net), 
            .I3(n23036), .O(n6958[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_12 (.CI(n22714), .I0(n6598[9]), .I1(n810_adj_4179), 
            .CO(n22715));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3368[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4303[22]), .I3(n22213), .O(n45_adj_4181)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_3378_11_lut (.I0(GND_net), .I1(n6598[8]), .I2(n737_adj_4152), 
            .I3(n22713), .O(n6575[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_11 (.CI(n22713), .I0(n6598[8]), .I1(n737_adj_4152), 
            .CO(n22714));
    SB_CARRY add_3404_17 (.CI(n23036), .I0(n6977[14]), .I1(GND_net), .CO(n23037));
    SB_LUT4 add_3378_10_lut (.I0(GND_net), .I1(n6598[7]), .I2(n664_adj_4151), 
            .I3(n22712), .O(n6575[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3404_16_lut (.I0(GND_net), .I1(n6977[13]), .I2(n1114_adj_4150), 
            .I3(n23035), .O(n6958[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_16 (.CI(n23035), .I0(n6977[13]), .I1(n1114_adj_4150), 
            .CO(n23036));
    SB_CARRY add_3378_10 (.CI(n22712), .I0(n6598[7]), .I1(n664_adj_4151), 
            .CO(n22713));
    SB_LUT4 add_3404_15_lut (.I0(GND_net), .I1(n6977[12]), .I2(n1041_adj_4149), 
            .I3(n23034), .O(n6958[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24361_4_lut (.I0(n21_adj_4180), .I1(n19_adj_4174), .I2(n17_adj_4172), 
            .I3(n9_adj_4171), .O(n29424));
    defparam i24361_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3378_9_lut (.I0(GND_net), .I1(n6598[6]), .I2(n591_adj_4147), 
            .I3(n22711), .O(n6575[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24354_4_lut (.I0(n27), .I1(n15_adj_4170), .I2(n13_adj_4164), 
            .I3(n11_adj_4161), .O(n29417));
    defparam i24354_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3404_15 (.CI(n23034), .I0(n6977[12]), .I1(n1041_adj_4149), 
            .CO(n23035));
    SB_LUT4 add_3404_14_lut (.I0(GND_net), .I1(n6977[11]), .I2(n968_adj_4144), 
            .I3(n23033), .O(n6958[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_14 (.CI(n23033), .I0(n6977[11]), .I1(n968_adj_4144), 
            .CO(n23034));
    SB_LUT4 duty_23__I_831_i12_3_lut (.I0(duty_23__N_3492[7]), .I1(duty_23__N_3492[16]), 
            .I2(n33), .I3(GND_net), .O(n12_adj_4182));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i10_3_lut (.I0(duty_23__N_3492[5]), .I1(duty_23__N_3492[6]), 
            .I2(n13_adj_4164), .I3(GND_net), .O(n10_adj_4183));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i30_3_lut (.I0(n12_adj_4182), .I1(duty_23__N_3492[17]), 
            .I2(n35_adj_4160), .I3(GND_net), .O(n30));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3378_9 (.CI(n22711), .I0(n6598[6]), .I1(n591_adj_4147), 
            .CO(n22712));
    SB_LUT4 add_3378_8_lut (.I0(GND_net), .I1(n6598[5]), .I2(n518_adj_4143), 
            .I3(n22710), .O(n6575[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_8 (.CI(n22710), .I0(n6598[5]), .I1(n518_adj_4143), 
            .CO(n22711));
    SB_LUT4 add_3404_13_lut (.I0(GND_net), .I1(n6977[10]), .I2(n895_adj_4142), 
            .I3(n23032), .O(n6958[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3378_7_lut (.I0(GND_net), .I1(n6598[4]), .I2(n445_adj_4141), 
            .I3(n22709), .O(n6575[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_13 (.CI(n23032), .I0(n6977[10]), .I1(n895_adj_4142), 
            .CO(n23033));
    SB_LUT4 i24635_4_lut (.I0(n13_adj_4164), .I1(n11_adj_4161), .I2(n9_adj_4171), 
            .I3(n29435), .O(n29701));
    defparam i24635_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24631_4_lut (.I0(n19_adj_4174), .I1(n17_adj_4172), .I2(n15_adj_4170), 
            .I3(n29701), .O(n29697));
    defparam i24631_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24940_4_lut (.I0(n25_adj_4159), .I1(n23_adj_4158), .I2(n21_adj_4180), 
            .I3(n29697), .O(n30006));
    defparam i24940_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3378_7 (.CI(n22709), .I0(n6598[4]), .I1(n445_adj_4141), 
            .CO(n22710));
    SB_LUT4 add_3378_6_lut (.I0(GND_net), .I1(n6598[3]), .I2(n372_adj_4138), 
            .I3(n22708), .O(n6575[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_6 (.CI(n22708), .I0(n6598[3]), .I1(n372_adj_4138), 
            .CO(n22709));
    SB_LUT4 add_3404_12_lut (.I0(GND_net), .I1(n6977[9]), .I2(n822_adj_4137), 
            .I3(n23031), .O(n6958[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_12 (.CI(n23031), .I0(n6977[9]), .I1(n822_adj_4137), 
            .CO(n23032));
    SB_LUT4 i24781_4_lut (.I0(n31), .I1(n29_adj_4156), .I2(n27), .I3(n30006), 
            .O(n29847));
    defparam i24781_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_3378_5_lut (.I0(GND_net), .I1(n6598[2]), .I2(n299_adj_4136), 
            .I3(n22707), .O(n6575[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24994_4_lut (.I0(n37), .I1(n35_adj_4160), .I2(n33), .I3(n29847), 
            .O(n30060));
    defparam i24994_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3404_11_lut (.I0(GND_net), .I1(n6977[8]), .I2(n749_adj_4135), 
            .I3(n23030), .O(n6958[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_5 (.CI(n22707), .I0(n6598[2]), .I1(n299_adj_4136), 
            .CO(n22708));
    SB_LUT4 add_3378_4_lut (.I0(GND_net), .I1(n6598[1]), .I2(n226_adj_4134), 
            .I3(n22706), .O(n6575[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_11 (.CI(n23030), .I0(n6977[8]), .I1(n749_adj_4135), 
            .CO(n23031));
    SB_LUT4 duty_23__I_831_i16_3_lut (.I0(duty_23__N_3492[9]), .I1(duty_23__N_3492[21]), 
            .I2(n43), .I3(GND_net), .O(n16_adj_4184));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3404_10_lut (.I0(GND_net), .I1(n6977[7]), .I2(n676_adj_4121), 
            .I3(n23029), .O(n6958[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_10 (.CI(n23029), .I0(n6977[7]), .I1(n676_adj_4121), 
            .CO(n23030));
    SB_LUT4 i24926_3_lut (.I0(n6_adj_4185), .I1(duty_23__N_3492[10]), .I2(n21_adj_4180), 
            .I3(GND_net), .O(n29992));   // verilog/motorControl.v(36[10:25])
    defparam i24926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3404_9_lut (.I0(GND_net), .I1(n6977[6]), .I2(n603_adj_4104), 
            .I3(n23028), .O(n6958[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_4 (.CI(n22706), .I0(n6598[1]), .I1(n226_adj_4134), 
            .CO(n22707));
    SB_CARRY add_3404_9 (.CI(n23028), .I0(n6977[6]), .I1(n603_adj_4104), 
            .CO(n23029));
    SB_LUT4 add_3378_3_lut (.I0(GND_net), .I1(n6598[0]), .I2(n153_adj_4103), 
            .I3(n22705), .O(n6575[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3404_8_lut (.I0(GND_net), .I1(n6977[5]), .I2(n530_adj_4102), 
            .I3(n23027), .O(n6958[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_5 (.CI(n21947), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n2552[3]), .CO(n21948));
    SB_CARRY add_3404_8 (.CI(n23027), .I0(n6977[5]), .I1(n530_adj_4102), 
            .CO(n23028));
    SB_CARRY unary_minus_5_add_3_24 (.CI(n22213), .I0(GND_net), .I1(n1_adj_4303[22]), 
            .CO(n22214));
    SB_LUT4 add_560_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n2552[2]), .I3(n21946), .O(\PID_CONTROLLER.integral_23__N_3392 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_3 (.CI(n22705), .I0(n6598[0]), .I1(n153_adj_4103), 
            .CO(n22706));
    SB_LUT4 add_3404_7_lut (.I0(GND_net), .I1(n6977[4]), .I2(n457_adj_4100), 
            .I3(n23026), .O(n6958[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3378_2_lut (.I0(GND_net), .I1(n11_adj_4099), .I2(n80_adj_4097), 
            .I3(GND_net), .O(n6575[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3378_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_7 (.CI(n23026), .I0(n6977[4]), .I1(n457_adj_4100), 
            .CO(n23027));
    SB_LUT4 add_3404_6_lut (.I0(GND_net), .I1(n6977[3]), .I2(n384_adj_4096), 
            .I3(n23025), .O(n6958[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_6 (.CI(n23025), .I0(n6977[3]), .I1(n384_adj_4096), 
            .CO(n23026));
    SB_LUT4 add_3404_5_lut (.I0(GND_net), .I1(n6977[2]), .I2(n311_adj_4094), 
            .I3(n23024), .O(n6958[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_5 (.CI(n23024), .I0(n6977[2]), .I1(n311_adj_4094), 
            .CO(n23025));
    SB_LUT4 add_3404_4_lut (.I0(GND_net), .I1(n6977[1]), .I2(n238_adj_4093), 
            .I3(n23023), .O(n6958[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_4 (.CI(n23023), .I0(n6977[1]), .I1(n238_adj_4093), 
            .CO(n23024));
    SB_LUT4 add_3404_3_lut (.I0(GND_net), .I1(n6977[0]), .I2(n165_adj_4092), 
            .I3(n23022), .O(n6958[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_3 (.CI(n23022), .I0(n6977[0]), .I1(n165_adj_4092), 
            .CO(n23023));
    SB_LUT4 add_3404_2_lut (.I0(GND_net), .I1(n23_adj_4090), .I2(n92_adj_4166), 
            .I3(GND_net), .O(n6958[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3404_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3404_2 (.CI(GND_net), .I0(n23_adj_4090), .I1(n92_adj_4166), 
            .CO(n23022));
    SB_LUT4 add_3403_19_lut (.I0(GND_net), .I1(n6958[16]), .I2(GND_net), 
            .I3(n23021), .O(n6938[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3403_18_lut (.I0(GND_net), .I1(n6958[15]), .I2(GND_net), 
            .I3(n23020), .O(n6938[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_18 (.CI(n23020), .I0(n6958[15]), .I1(GND_net), .CO(n23021));
    SB_LUT4 add_3403_17_lut (.I0(GND_net), .I1(n6958[14]), .I2(GND_net), 
            .I3(n23019), .O(n6938[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_17 (.CI(n23019), .I0(n6958[14]), .I1(GND_net), .CO(n23020));
    SB_LUT4 add_3403_16_lut (.I0(GND_net), .I1(n6958[13]), .I2(n1111_adj_4089), 
            .I3(n23018), .O(n6938[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_16 (.CI(n23018), .I0(n6958[13]), .I1(n1111_adj_4089), 
            .CO(n23019));
    SB_LUT4 add_3403_15_lut (.I0(GND_net), .I1(n6958[12]), .I2(n1038_adj_4088), 
            .I3(n23017), .O(n6938[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_15 (.CI(n23017), .I0(n6958[12]), .I1(n1038_adj_4088), 
            .CO(n23018));
    SB_LUT4 add_3403_14_lut (.I0(GND_net), .I1(n6958[11]), .I2(n965_adj_4087), 
            .I3(n23016), .O(n6938[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_14 (.CI(n23016), .I0(n6958[11]), .I1(n965_adj_4087), 
            .CO(n23017));
    SB_LUT4 add_3403_13_lut (.I0(GND_net), .I1(n6958[10]), .I2(n892_adj_4086), 
            .I3(n23015), .O(n6938[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_13 (.CI(n23015), .I0(n6958[10]), .I1(n892_adj_4086), 
            .CO(n23016));
    SB_LUT4 add_3403_12_lut (.I0(GND_net), .I1(n6958[9]), .I2(n819_adj_4085), 
            .I3(n23014), .O(n6938[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_12 (.CI(n23014), .I0(n6958[9]), .I1(n819_adj_4085), 
            .CO(n23015));
    SB_LUT4 add_3403_11_lut (.I0(GND_net), .I1(n6958[8]), .I2(n746_adj_4084), 
            .I3(n23013), .O(n6938[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3378_2 (.CI(GND_net), .I0(n11_adj_4099), .I1(n80_adj_4097), 
            .CO(n22705));
    SB_CARRY add_3403_11 (.CI(n23013), .I0(n6958[8]), .I1(n746_adj_4084), 
            .CO(n23014));
    SB_LUT4 add_3403_10_lut (.I0(GND_net), .I1(n6958[7]), .I2(n673_adj_4083), 
            .I3(n23012), .O(n6938[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24927_3_lut (.I0(n29992), .I1(duty_23__N_3492[11]), .I2(n23_adj_4158), 
            .I3(GND_net), .O(n29993));   // verilog/motorControl.v(36[10:25])
    defparam i24927_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3403_10 (.CI(n23012), .I0(n6958[7]), .I1(n673_adj_4083), 
            .CO(n23013));
    SB_LUT4 duty_23__I_831_i8_3_lut (.I0(duty_23__N_3492[4]), .I1(duty_23__N_3492[8]), 
            .I2(n17_adj_4172), .I3(GND_net), .O(n8_adj_4186));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i24_3_lut (.I0(n16_adj_4184), .I1(duty_23__N_3492[22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_4187));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24339_4_lut (.I0(n43), .I1(n25_adj_4159), .I2(n23_adj_4158), 
            .I3(n29424), .O(n29402));
    defparam i24339_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24803_4_lut (.I0(n24_adj_4187), .I1(n8_adj_4186), .I2(n45), 
            .I3(n29400), .O(n29869));   // verilog/motorControl.v(36[10:25])
    defparam i24803_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24868_3_lut (.I0(n29993), .I1(duty_23__N_3492[12]), .I2(n25_adj_4159), 
            .I3(GND_net), .O(n29934));   // verilog/motorControl.v(36[10:25])
    defparam i24868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3403_9_lut (.I0(GND_net), .I1(n6958[6]), .I2(n600_adj_4082), 
            .I3(n23011), .O(n6938[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i4_4_lut (.I0(duty_23__N_3492[0]), .I1(duty_23__N_3492[1]), 
            .I2(PWMLimit[1]), .I3(n1_adj_4304[0]), .O(n4_adj_4188));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i4_4_lut.LUT_INIT = 16'h8e0c;
    SB_CARRY add_3403_9 (.CI(n23011), .I0(n6958[6]), .I1(n600_adj_4082), 
            .CO(n23012));
    SB_LUT4 add_3403_8_lut (.I0(GND_net), .I1(n6958[5]), .I2(n527_adj_4081), 
            .I3(n23010), .O(n6938[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_8 (.CI(n23010), .I0(n6958[5]), .I1(n527_adj_4081), 
            .CO(n23011));
    SB_LUT4 i24916_3_lut (.I0(n4_adj_4188), .I1(duty_23__N_3492[13]), .I2(n27), 
            .I3(GND_net), .O(n29982));   // verilog/motorControl.v(36[10:25])
    defparam i24916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3403_7_lut (.I0(GND_net), .I1(n6958[4]), .I2(n454_adj_4080), 
            .I3(n23009), .O(n6938[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_7 (.CI(n23009), .I0(n6958[4]), .I1(n454_adj_4080), 
            .CO(n23010));
    SB_LUT4 add_3403_6_lut (.I0(GND_net), .I1(n6958[3]), .I2(n381_adj_4079), 
            .I3(n23008), .O(n6938[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_6 (.CI(n23008), .I0(n6958[3]), .I1(n381_adj_4079), 
            .CO(n23009));
    SB_LUT4 add_3403_5_lut (.I0(GND_net), .I1(n6958[2]), .I2(n308_adj_4078), 
            .I3(n23007), .O(n6938[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_5 (.CI(n23007), .I0(n6958[2]), .I1(n308_adj_4078), 
            .CO(n23008));
    SB_LUT4 add_3403_4_lut (.I0(GND_net), .I1(n6958[1]), .I2(n235_adj_4077), 
            .I3(n23006), .O(n6938[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17893_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4189), 
            .I3(n6830[1]), .O(n6));   // verilog/motorControl.v(34[16:22])
    defparam i17893_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i24917_3_lut (.I0(n29982), .I1(duty_23__N_3492[14]), .I2(n29_adj_4156), 
            .I3(GND_net), .O(n29983));   // verilog/motorControl.v(36[10:25])
    defparam i24917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24350_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4156), .I3(n29417), 
            .O(n29413));
    defparam i24350_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25004_4_lut (.I0(n30), .I1(n10_adj_4183), .I2(n35_adj_4160), 
            .I3(n29411), .O(n30070));   // verilog/motorControl.v(36[10:25])
    defparam i25004_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i2_3_lut_4_lut_adj_1443 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n6830[1]), 
            .I3(n4_adj_4189), .O(n6823[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1443.LUT_INIT = 16'h8778;
    SB_LUT4 i24870_3_lut (.I0(n29983), .I1(duty_23__N_3492[15]), .I2(n31), 
            .I3(GND_net), .O(n29936));   // verilog/motorControl.v(36[10:25])
    defparam i24870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25053_4_lut (.I0(n29936), .I1(n30070), .I2(n35_adj_4160), 
            .I3(n29413), .O(n30119));   // verilog/motorControl.v(36[10:25])
    defparam i25053_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25054_3_lut (.I0(n30119), .I1(duty_23__N_3492[18]), .I2(n37), 
            .I3(GND_net), .O(n30120));   // verilog/motorControl.v(36[10:25])
    defparam i25054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25035_3_lut (.I0(n30120), .I1(duty_23__N_3492[19]), .I2(n39), 
            .I3(GND_net), .O(n30101));   // verilog/motorControl.v(36[10:25])
    defparam i25035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24341_4_lut (.I0(n43), .I1(n41_adj_4154), .I2(n39), .I3(n30060), 
            .O(n29404));
    defparam i24341_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24958_4_lut (.I0(n29934), .I1(n29869), .I2(n45), .I3(n29402), 
            .O(n30024));   // verilog/motorControl.v(36[10:25])
    defparam i24958_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_4_lut_adj_1444 (.I0(n4_adj_4190), .I1(\Ki[3] ), .I2(n7133[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [19]), .O(n7127[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1444.LUT_INIT = 16'h965a;
    SB_CARRY add_3403_4 (.CI(n23006), .I0(n6958[1]), .I1(n235_adj_4077), 
            .CO(n23007));
    SB_LUT4 i25023_3_lut (.I0(n30101), .I1(duty_23__N_3492[20]), .I2(n41_adj_4154), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(36[10:25])
    defparam i25023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3403_3_lut (.I0(GND_net), .I1(n6958[0]), .I2(n162_adj_4076), 
            .I3(n23005), .O(n6938[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3403_3 (.CI(n23005), .I0(n6958[0]), .I1(n162_adj_4076), 
            .CO(n23006));
    SB_LUT4 add_3403_2_lut (.I0(GND_net), .I1(n20_adj_4075), .I2(n89), 
            .I3(GND_net), .O(n6938[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3403_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24960_4_lut (.I0(n40), .I1(n30024), .I2(n45), .I3(n29404), 
            .O(n30026));   // verilog/motorControl.v(36[10:25])
    defparam i24960_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24961_3_lut (.I0(n30026), .I1(PWMLimit[23]), .I2(duty_23__N_3492[23]), 
            .I3(GND_net), .O(duty_23__N_3491));   // verilog/motorControl.v(36[10:25])
    defparam i24961_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_560_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n2552[7]), .I3(n21951), .O(\PID_CONTROLLER.integral_23__N_3392 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3492[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4192));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3403_2 (.CI(GND_net), .I0(n20_adj_4075), .I1(n89), .CO(n23005));
    SB_LUT4 add_3402_20_lut (.I0(GND_net), .I1(n6938[17]), .I2(GND_net), 
            .I3(n23004), .O(n6917[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n22008), 
            .O(duty_23__N_3492[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3492[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4193));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1445 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n6830[0]), 
            .I3(n21652), .O(n6823[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1445.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3492[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4195));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3492[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4196));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3402_19_lut (.I0(GND_net), .I1(n6938[16]), .I2(GND_net), 
            .I3(n23003), .O(n6917[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4303[21]), .I3(n22212), .O(n43_adj_4197)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3402_19 (.CI(n23003), .I0(n6938[16]), .I1(GND_net), .CO(n23004));
    SB_LUT4 add_3402_18_lut (.I0(GND_net), .I1(n6938[15]), .I2(GND_net), 
            .I3(n23002), .O(n6917[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_18 (.CI(n23002), .I0(n6938[15]), .I1(GND_net), .CO(n23003));
    SB_LUT4 i17885_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n21652), 
            .I3(n6830[0]), .O(n4_adj_4189));   // verilog/motorControl.v(34[16:22])
    defparam i17885_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n6551[21]), .I2(GND_net), 
            .I3(n22704), .O(n4998[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_12_5 (.CI(n22008), .I0(n106[3]), .I1(n155[3]), .CO(n22009));
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3492[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4198));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n22007), 
            .O(duty_23__N_3492[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3492[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4199));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3402_17_lut (.I0(GND_net), .I1(n6938[14]), .I2(GND_net), 
            .I3(n23001), .O(n6917[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_17 (.CI(n23001), .I0(n6938[14]), .I1(GND_net), .CO(n23002));
    SB_LUT4 add_3402_16_lut (.I0(GND_net), .I1(n6938[13]), .I2(n1108), 
            .I3(n23000), .O(n6917[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_16 (.CI(n23000), .I0(n6938[13]), .I1(n1108), .CO(n23001));
    SB_LUT4 add_3402_15_lut (.I0(GND_net), .I1(n6938[12]), .I2(n1035), 
            .I3(n22999), .O(n6917[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3492[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4200));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3402_15 (.CI(n22999), .I0(n6938[12]), .I1(n1035), .CO(n23000));
    SB_LUT4 add_3402_14_lut (.I0(GND_net), .I1(n6938[11]), .I2(n962), 
            .I3(n22998), .O(n6917[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_14 (.CI(n22998), .I0(n6938[11]), .I1(n962), .CO(n22999));
    SB_LUT4 add_3402_13_lut (.I0(GND_net), .I1(n6938[10]), .I2(n889), 
            .I3(n22997), .O(n6917[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_13 (.CI(n22997), .I0(n6938[10]), .I1(n889), .CO(n22998));
    SB_LUT4 add_3402_12_lut (.I0(GND_net), .I1(n6938[9]), .I2(n816), .I3(n22996), 
            .O(n6917[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_12 (.CI(n22996), .I0(n6938[9]), .I1(n816), .CO(n22997));
    SB_LUT4 add_3402_11_lut (.I0(GND_net), .I1(n6938[8]), .I2(n743), .I3(n22995), 
            .O(n6917[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3492[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4201));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3402_11 (.CI(n22995), .I0(n6938[8]), .I1(n743), .CO(n22996));
    SB_LUT4 add_3402_10_lut (.I0(GND_net), .I1(n6938[7]), .I2(n670), .I3(n22994), 
            .O(n6917[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_10 (.CI(n22994), .I0(n6938[7]), .I1(n670), .CO(n22995));
    SB_LUT4 add_3402_9_lut (.I0(GND_net), .I1(n6938[6]), .I2(n597_adj_4073), 
            .I3(n22993), .O(n6917[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_9 (.CI(n22993), .I0(n6938[6]), .I1(n597_adj_4073), 
            .CO(n22994));
    SB_LUT4 add_3402_8_lut (.I0(GND_net), .I1(n6938[5]), .I2(n524_adj_4072), 
            .I3(n22992), .O(n6917[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15186_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15186_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3492[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4202));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n6551[20]), .I2(GND_net), 
            .I3(n22703), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17872_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n6823[0]));   // verilog/motorControl.v(34[16:22])
    defparam i17872_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY mult_10_add_1225_23 (.CI(n22703), .I0(n6551[20]), .I1(GND_net), 
            .CO(n22704));
    SB_LUT4 i17874_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n21652));   // verilog/motorControl.v(34[16:22])
    defparam i17874_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3492[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4203));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3402_8 (.CI(n22992), .I0(n6938[5]), .I1(n524_adj_4072), 
            .CO(n22993));
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3492[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4205));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3492[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4206));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_4 (.CI(n22007), .I0(n106[2]), .I1(n155[2]), .CO(n22008));
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3492[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4207));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3402_7_lut (.I0(GND_net), .I1(n6938[4]), .I2(n451_adj_4070), 
            .I3(n22991), .O(n6917[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_7 (.CI(n22991), .I0(n6938[4]), .I1(n451_adj_4070), 
            .CO(n22992));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n6551[19]), .I2(GND_net), 
            .I3(n22702), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n22212), .I0(GND_net), .I1(n1_adj_4303[21]), 
            .CO(n22213));
    SB_LUT4 add_3402_6_lut (.I0(GND_net), .I1(n6938[3]), .I2(n378_adj_4069), 
            .I3(n22990), .O(n6917[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n22702), .I0(n6551[19]), .I1(GND_net), 
            .CO(n22703));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n6551[18]), .I2(GND_net), 
            .I3(n22701), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3492[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4208));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1446 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3392 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [20]), .O(n12_adj_4209));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1446.LUT_INIT = 16'h9c50;
    SB_CARRY add_3402_6 (.CI(n22990), .I0(n6938[3]), .I1(n378_adj_4069), 
            .CO(n22991));
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3492[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4211));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3402_5_lut (.I0(GND_net), .I1(n6938[2]), .I2(n305_adj_4068), 
            .I3(n22989), .O(n6917[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_5 (.CI(n22989), .I0(n6938[2]), .I1(n305_adj_4068), 
            .CO(n22990));
    SB_LUT4 add_3402_4_lut (.I0(GND_net), .I1(n6938[1]), .I2(n232_adj_4067), 
            .I3(n22988), .O(n6917[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3492[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4212));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3402_4 (.CI(n22988), .I0(n6938[1]), .I1(n232_adj_4067), 
            .CO(n22989));
    SB_LUT4 add_3402_3_lut (.I0(GND_net), .I1(n6938[0]), .I2(n159_adj_4066), 
            .I3(n22987), .O(n6917[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_3 (.CI(n22987), .I0(n6938[0]), .I1(n159_adj_4066), 
            .CO(n22988));
    SB_LUT4 add_3402_2_lut (.I0(GND_net), .I1(n17_adj_4065), .I2(n86_adj_4064), 
            .I3(GND_net), .O(n6917[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3492[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4213));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3402_2 (.CI(GND_net), .I0(n17_adj_4065), .I1(n86_adj_4064), 
            .CO(n22987));
    SB_CARRY mult_10_add_1225_21 (.CI(n22701), .I0(n6551[18]), .I1(GND_net), 
            .CO(n22702));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n6551[17]), .I2(GND_net), 
            .I3(n22700), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3401_21_lut (.I0(GND_net), .I1(n6917[18]), .I2(GND_net), 
            .I3(n22986), .O(n6895[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3492[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4214));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3401_20_lut (.I0(GND_net), .I1(n6917[17]), .I2(GND_net), 
            .I3(n22985), .O(n6895[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_20 (.CI(n22985), .I0(n6917[17]), .I1(GND_net), .CO(n22986));
    SB_LUT4 add_3401_19_lut (.I0(GND_net), .I1(n6917[16]), .I2(GND_net), 
            .I3(n22984), .O(n6895[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n22700), .I0(n6551[17]), .I1(GND_net), 
            .CO(n22701));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n6551[16]), .I2(GND_net), 
            .I3(n22699), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_19 (.CI(n22984), .I0(n6917[16]), .I1(GND_net), .CO(n22985));
    SB_CARRY mult_10_add_1225_19 (.CI(n22699), .I0(n6551[16]), .I1(GND_net), 
            .CO(n22700));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4303[20]), .I3(n22211), .O(n41_adj_4215)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3401_18_lut (.I0(GND_net), .I1(n6917[15]), .I2(GND_net), 
            .I3(n22983), .O(n6895[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n6551[15]), .I2(GND_net), 
            .I3(n22698), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n22698), .I0(n6551[15]), .I1(GND_net), 
            .CO(n22699));
    SB_CARRY add_3401_18 (.CI(n22983), .I0(n6917[15]), .I1(GND_net), .CO(n22984));
    SB_LUT4 add_3401_17_lut (.I0(GND_net), .I1(n6917[14]), .I2(GND_net), 
            .I3(n22982), .O(n6895[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n22211), .I0(GND_net), .I1(n1_adj_4303[20]), 
            .CO(n22212));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n6551[14]), .I2(GND_net), 
            .I3(n22697), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_17 (.CI(n22982), .I0(n6917[14]), .I1(GND_net), .CO(n22983));
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3492[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4217));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_17 (.CI(n22697), .I0(n6551[14]), .I1(GND_net), 
            .CO(n22698));
    SB_LUT4 i24325_4_lut (.I0(n21_adj_4217), .I1(n19_adj_4214), .I2(n17_adj_4213), 
            .I3(n9_adj_4212), .O(n29388));
    defparam i24325_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24319_4_lut (.I0(n27_adj_4211), .I1(n15_adj_4208), .I2(n13_adj_4207), 
            .I3(n11_adj_4206), .O(n29382));
    defparam i24319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3401_16_lut (.I0(GND_net), .I1(n6917[13]), .I2(n1105_adj_4062), 
            .I3(n22981), .O(n6895[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_16 (.CI(n22981), .I0(n6917[13]), .I1(n1105_adj_4062), 
            .CO(n22982));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n22006), 
            .O(duty_23__N_3492[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3401_15_lut (.I0(GND_net), .I1(n6917[12]), .I2(n1032_adj_4061), 
            .I3(n22980), .O(n6895[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18023_4_lut (.I0(n7127[2]), .I1(\Ki[4] ), .I2(n6_adj_4139), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [18]), .O(n8_adj_4219));   // verilog/motorControl.v(34[25:36])
    defparam i18023_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n6551[13]), .I2(n1096_adj_4060), 
            .I3(n22696), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n22696), .I0(n6551[13]), .I1(n1096_adj_4060), 
            .CO(n22697));
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_46_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n30965));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_46_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3401_15 (.CI(n22980), .I0(n6917[12]), .I1(n1032_adj_4061), 
            .CO(n22981));
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4205), 
            .I3(GND_net), .O(n12_adj_4220));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24710_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4162), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4146), .O(n29776));
    defparam i24710_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n6551[12]), .I2(n1023_adj_4059), 
            .I3(n22695), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1447 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3392 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [21]), .O(n11_adj_4221));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1447.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4303[19]), .I3(n22210), .O(n39_adj_4222)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_1225_15 (.CI(n22695), .I0(n6551[12]), .I1(n1023_adj_4059), 
            .CO(n22696));
    SB_LUT4 i24708_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n30965), 
            .I2(IntegralLimit[11]), .I3(n29776), .O(n29774));
    defparam i24708_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n6551[11]), .I2(n950_adj_4057), 
            .I3(n22694), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3401_14_lut (.I0(GND_net), .I1(n6917[11]), .I2(n959_adj_4056), 
            .I3(n22979), .O(n6895[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_14 (.CI(n22979), .I0(n6917[11]), .I1(n959_adj_4056), 
            .CO(n22980));
    SB_LUT4 add_3401_13_lut (.I0(GND_net), .I1(n6917[10]), .I2(n886_adj_4055), 
            .I3(n22978), .O(n6895[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_13 (.CI(n22978), .I0(n6917[10]), .I1(n886_adj_4055), 
            .CO(n22979));
    SB_CARRY unary_minus_5_add_3_21 (.CI(n22210), .I0(GND_net), .I1(n1_adj_4303[19]), 
            .CO(n22211));
    SB_LUT4 add_3401_12_lut (.I0(GND_net), .I1(n6917[9]), .I2(n813_adj_4053), 
            .I3(n22977), .O(n6895[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_40_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n30959));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_40_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4207), 
            .I3(GND_net), .O(n10_adj_4223));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4303[18]), .I3(n22209), .O(n37_adj_4224)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n22209), .I0(GND_net), .I1(n1_adj_4303[18]), 
            .CO(n22210));
    SB_CARRY mult_10_add_1225_14 (.CI(n22694), .I0(n6551[11]), .I1(n950_adj_4057), 
            .CO(n22695));
    SB_CARRY add_3401_12 (.CI(n22977), .I0(n6917[9]), .I1(n813_adj_4053), 
            .CO(n22978));
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4220), .I1(n257[17]), .I2(n35_adj_4203), 
            .I3(GND_net), .O(n30_adj_4225));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24392_4_lut (.I0(n27_adj_4226), .I1(n15_adj_4227), .I2(n13_adj_4228), 
            .I3(n11_adj_4229), .O(n29455));
    defparam i24392_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24401_4_lut (.I0(n21_adj_4230), .I1(n19_adj_4231), .I2(n17_adj_4232), 
            .I3(n9_adj_4233), .O(n29464));
    defparam i24401_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_4197), .I3(GND_net), 
            .O(n16_adj_4234));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n6551[10]), .I2(n877_adj_4051), 
            .I3(n22693), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n22693), .I0(n6551[10]), .I1(n877_adj_4051), 
            .CO(n22694));
    SB_LUT4 i24374_2_lut (.I0(n43_adj_4197), .I1(n19_adj_4231), .I2(GND_net), 
            .I3(GND_net), .O(n29437));
    defparam i24374_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4232), .I3(GND_net), 
            .O(n8_adj_4235));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4303[17]), .I3(n22208), .O(n35_adj_4236)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3401_11_lut (.I0(GND_net), .I1(n6917[8]), .I2(n740_adj_4049), 
            .I3(n22976), .O(n6895[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4234), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_4181), .I3(GND_net), 
            .O(n24_adj_4237));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_3401_11 (.CI(n22976), .I0(n6917[8]), .I1(n740_adj_4049), 
            .CO(n22977));
    SB_LUT4 i24601_4_lut (.I0(n13_adj_4207), .I1(n11_adj_4206), .I2(n9_adj_4212), 
            .I3(n29398), .O(n29667));
    defparam i24601_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24597_4_lut (.I0(n19_adj_4214), .I1(n17_adj_4213), .I2(n15_adj_4208), 
            .I3(n29667), .O(n29663));
    defparam i24597_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24932_4_lut (.I0(n25_adj_4200), .I1(n23_adj_4199), .I2(n21_adj_4217), 
            .I3(n29663), .O(n29998));
    defparam i24932_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24765_4_lut (.I0(n31_adj_4202), .I1(n29_adj_4201), .I2(n27_adj_4211), 
            .I3(n29998), .O(n29831));
    defparam i24765_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i18054_4_lut (.I0(n7133[1]), .I1(\Ki[3] ), .I2(n4_adj_4190), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [19]), .O(n6_adj_4238));   // verilog/motorControl.v(34[25:36])
    defparam i18054_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i24992_4_lut (.I0(n37_adj_4198), .I1(n35_adj_4203), .I2(n33_adj_4205), 
            .I3(n29831), .O(n30058));
    defparam i24992_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4196), 
            .I3(GND_net), .O(n16_adj_4239));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24912_3_lut (.I0(n6_adj_4240), .I1(n257[10]), .I2(n21_adj_4217), 
            .I3(GND_net), .O(n29978));   // verilog/motorControl.v(38[19:35])
    defparam i24912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17911_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n6830[0]));   // verilog/motorControl.v(34[16:22])
    defparam i17911_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24913_3_lut (.I0(n29978), .I1(n257[11]), .I2(n23_adj_4199), 
            .I3(GND_net), .O(n29979));   // verilog/motorControl.v(38[19:35])
    defparam i24913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4213), 
            .I3(GND_net), .O(n8_adj_4241));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4239), .I1(n257[22]), .I2(n45_adj_4195), 
            .I3(GND_net), .O(n24_adj_4242));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24305_4_lut (.I0(n43_adj_4196), .I1(n25_adj_4200), .I2(n23_adj_4199), 
            .I3(n29388), .O(n29368));
    defparam i24305_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24805_4_lut (.I0(n24_adj_4242), .I1(n8_adj_4241), .I2(n45_adj_4195), 
            .I3(n29366), .O(n29871));   // verilog/motorControl.v(38[19:35])
    defparam i24805_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24874_3_lut (.I0(n29979), .I1(n257[12]), .I2(n25_adj_4200), 
            .I3(GND_net), .O(n29940));   // verilog/motorControl.v(38[19:35])
    defparam i24874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3492[0]), .I1(n257[1]), 
            .I2(duty_23__N_3492[1]), .I3(n257[0]), .O(n4_adj_4243));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i17913_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n21695));   // verilog/motorControl.v(34[16:22])
    defparam i17913_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i24910_3_lut (.I0(n4_adj_4243), .I1(n257[13]), .I2(n27_adj_4211), 
            .I3(GND_net), .O(n29976));   // verilog/motorControl.v(38[19:35])
    defparam i24910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24911_3_lut (.I0(n29976), .I1(n257[14]), .I2(n29_adj_4201), 
            .I3(GND_net), .O(n29977));   // verilog/motorControl.v(38[19:35])
    defparam i24911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24315_4_lut (.I0(n33_adj_4205), .I1(n31_adj_4202), .I2(n29_adj_4201), 
            .I3(n29382), .O(n29378));
    defparam i24315_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25006_4_lut (.I0(n30_adj_4225), .I1(n10_adj_4223), .I2(n35_adj_4203), 
            .I3(n29376), .O(n30072));   // verilog/motorControl.v(38[19:35])
    defparam i25006_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24876_3_lut (.I0(n29977), .I1(n257[15]), .I2(n31_adj_4202), 
            .I3(GND_net), .O(n29942));   // verilog/motorControl.v(38[19:35])
    defparam i24876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25055_4_lut (.I0(n29942), .I1(n30072), .I2(n35_adj_4203), 
            .I3(n29378), .O(n30121));   // verilog/motorControl.v(38[19:35])
    defparam i25055_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i18089_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3392 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [21]), .O(n21886));   // verilog/motorControl.v(34[25:36])
    defparam i18089_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25056_3_lut (.I0(n30121), .I1(n257[18]), .I2(n37_adj_4198), 
            .I3(GND_net), .O(n30122));   // verilog/motorControl.v(38[19:35])
    defparam i25056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25033_3_lut (.I0(n30122), .I1(n257[19]), .I2(n39_adj_4192), 
            .I3(GND_net), .O(n30099));   // verilog/motorControl.v(38[19:35])
    defparam i25033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24307_4_lut (.I0(n43_adj_4196), .I1(n41_adj_4193), .I2(n39_adj_4192), 
            .I3(n30058), .O(n29370));
    defparam i24307_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24964_4_lut (.I0(n29940), .I1(n29871), .I2(n45_adj_4195), 
            .I3(n29368), .O(n30030));   // verilog/motorControl.v(38[19:35])
    defparam i24964_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3401_10_lut (.I0(GND_net), .I1(n6917[7]), .I2(n667_adj_4048), 
            .I3(n22975), .O(n6895[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_10 (.CI(n22975), .I0(n6917[7]), .I1(n667_adj_4048), 
            .CO(n22976));
    SB_LUT4 add_3401_9_lut (.I0(GND_net), .I1(n6917[6]), .I2(n594), .I3(n22974), 
            .O(n6895[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25025_3_lut (.I0(n30099), .I1(n257[20]), .I2(n41_adj_4193), 
            .I3(GND_net), .O(n40_adj_4244));   // verilog/motorControl.v(38[19:35])
    defparam i25025_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3401_9 (.CI(n22974), .I0(n6917[6]), .I1(n594), .CO(n22975));
    SB_LUT4 add_3401_8_lut (.I0(GND_net), .I1(n6917[5]), .I2(n521), .I3(n22973), 
            .O(n6895[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_8 (.CI(n22973), .I0(n6917[5]), .I1(n521), .CO(n22974));
    SB_LUT4 add_3401_7_lut (.I0(GND_net), .I1(n6917[4]), .I2(n448), .I3(n22972), 
            .O(n6895[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24966_4_lut (.I0(n40_adj_4244), .I1(n30030), .I2(n45_adj_4195), 
            .I3(n29370), .O(n30032));   // verilog/motorControl.v(38[19:35])
    defparam i24966_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3401_7 (.CI(n22972), .I0(n6917[4]), .I1(n448), .CO(n22973));
    SB_LUT4 i24433_2_lut (.I0(n7_adj_4245), .I1(n5_adj_4246), .I2(GND_net), 
            .I3(GND_net), .O(n29496));
    defparam i24433_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24680_4_lut (.I0(n13_adj_4228), .I1(n11_adj_4229), .I2(n9_adj_4233), 
            .I3(n29496), .O(n29746));
    defparam i24680_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24676_4_lut (.I0(n19_adj_4231), .I1(n17_adj_4232), .I2(n15_adj_4227), 
            .I3(n29746), .O(n29742));
    defparam i24676_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24970_4_lut (.I0(n25_adj_4247), .I1(n23_adj_4248), .I2(n21_adj_4230), 
            .I3(n29742), .O(n30036));
    defparam i24970_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24797_4_lut (.I0(n31_adj_4249), .I1(n29_adj_4250), .I2(n27_adj_4226), 
            .I3(n30036), .O(n29863));
    defparam i24797_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24996_4_lut (.I0(n37_adj_4224), .I1(n35_adj_4236), .I2(n33_adj_4251), 
            .I3(n29863), .O(n30062));
    defparam i24996_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3401_6_lut (.I0(GND_net), .I1(n6917[3]), .I2(n375), .I3(n22971), 
            .O(n6895[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n6551[9]), .I2(n804_adj_4047), 
            .I3(n22692), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n22692), .I0(n6551[9]), .I1(n804_adj_4047), 
            .CO(n22693));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n6551[8]), .I2(n731_adj_4046), 
            .I3(n22691), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n22691), .I0(n6551[8]), .I1(n731_adj_4046), 
            .CO(n22692));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n6551[7]), .I2(n658_adj_4043), 
            .I3(n22690), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n22208), .I0(GND_net), .I1(n1_adj_4303[17]), 
            .CO(n22209));
    SB_CARRY add_3401_6 (.CI(n22971), .I0(n6917[3]), .I1(n375), .CO(n22972));
    SB_CARRY mult_10_add_1225_10 (.CI(n22690), .I0(n6551[7]), .I1(n658_adj_4043), 
            .CO(n22691));
    SB_LUT4 add_3401_5_lut (.I0(GND_net), .I1(n6917[2]), .I2(n302), .I3(n22970), 
            .O(n6895[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_3 (.CI(n22006), .I0(n106[1]), .I1(n155[1]), .CO(n22007));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n6551[6]), .I2(n585_adj_4042), 
            .I3(n22689), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_5 (.CI(n22970), .I0(n6917[2]), .I1(n302), .CO(n22971));
    SB_LUT4 add_3401_4_lut (.I0(GND_net), .I1(n6917[1]), .I2(n229), .I3(n22969), 
            .O(n6895[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_4 (.CI(n22969), .I0(n6917[1]), .I1(n229), .CO(n22970));
    SB_LUT4 add_3401_3_lut (.I0(GND_net), .I1(n6917[0]), .I2(n156), .I3(n22968), 
            .O(n6895[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24967_3_lut (.I0(n30032), .I1(duty_23__N_3492[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4252));   // verilog/motorControl.v(38[19:35])
    defparam i24967_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3401_3 (.CI(n22968), .I0(n6917[0]), .I1(n156), .CO(n22969));
    SB_LUT4 add_3401_2_lut (.I0(GND_net), .I1(n14_adj_4040), .I2(n83), 
            .I3(GND_net), .O(n6895[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3401_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3401_2 (.CI(GND_net), .I0(n14_adj_4040), .I1(n83), .CO(n22968));
    SB_LUT4 add_3400_22_lut (.I0(GND_net), .I1(n6895[19]), .I2(GND_net), 
            .I3(n22967), .O(n6872[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3492[0]), .I1(n257[0]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4303[16]), .I3(n22207), .O(n33_adj_4251)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n22207), .I0(GND_net), .I1(n1_adj_4303[16]), 
            .CO(n22208));
    SB_LUT4 i8_4_lut_adj_1448 (.I0(n6_adj_4238), .I1(n11_adj_4221), .I2(n8_adj_4219), 
            .I3(n12_adj_4209), .O(n18_adj_4253));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3467[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3400_21_lut (.I0(GND_net), .I1(n6895[18]), .I2(GND_net), 
            .I3(n22966), .O(n6872[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_21 (.CI(n22966), .I0(n6895[18]), .I1(GND_net), .CO(n22967));
    SB_CARRY mult_10_add_1225_9 (.CI(n22689), .I0(n6551[6]), .I1(n585_adj_4042), 
            .CO(n22690));
    SB_LUT4 add_3400_20_lut (.I0(GND_net), .I1(n6895[17]), .I2(GND_net), 
            .I3(n22965), .O(n6872[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_20 (.CI(n22965), .I0(n6895[17]), .I1(GND_net), .CO(n22966));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n6551[5]), .I2(n512_adj_4038), 
            .I3(n22688), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_8 (.CI(n22688), .I0(n6551[5]), .I1(n512_adj_4038), 
            .CO(n22689));
    SB_LUT4 add_3400_19_lut (.I0(GND_net), .I1(n6895[16]), .I2(GND_net), 
            .I3(n22964), .O(n6872[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n6551[4]), .I2(n439_adj_4037), 
            .I3(n22687), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n22687), .I0(n6551[4]), .I1(n439_adj_4037), 
            .CO(n22688));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n6551[3]), .I2(n366_adj_4036), 
            .I3(n22686), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_19 (.CI(n22964), .I0(n6895[16]), .I1(GND_net), .CO(n22965));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4303[15]), .I3(n22206), .O(n31_adj_4249)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3400_18_lut (.I0(GND_net), .I1(n6895[15]), .I2(GND_net), 
            .I3(n22963), .O(n6872[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n22686), .I0(n6551[3]), .I1(n366_adj_4036), 
            .CO(n22687));
    SB_CARRY add_3400_18 (.CI(n22963), .I0(n6895[15]), .I1(GND_net), .CO(n22964));
    SB_LUT4 add_3400_17_lut (.I0(GND_net), .I1(n6895[14]), .I2(GND_net), 
            .I3(n22962), .O(n6872[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_17 (.CI(n22962), .I0(n6895[14]), .I1(GND_net), .CO(n22963));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n6551[2]), .I2(n293_adj_4034), 
            .I3(n22685), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_16_lut (.I0(GND_net), .I1(n6895[13]), .I2(n1102), 
            .I3(n22961), .O(n6872[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n22685), .I0(n6551[2]), .I1(n293_adj_4034), 
            .CO(n22686));
    SB_CARRY add_3400_16 (.CI(n22961), .I0(n6895[13]), .I1(n1102), .CO(n22962));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n6551[1]), .I2(n220_adj_4033), 
            .I3(n22684), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_15_lut (.I0(GND_net), .I1(n6895[12]), .I2(n1029), 
            .I3(n22960), .O(n6872[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_15 (.CI(n22960), .I0(n6895[12]), .I1(n1029), .CO(n22961));
    SB_CARRY mult_10_add_1225_4 (.CI(n22684), .I0(n6551[1]), .I1(n220_adj_4033), 
            .CO(n22685));
    SB_LUT4 add_3400_14_lut (.I0(GND_net), .I1(n6895[11]), .I2(n956), 
            .I3(n22959), .O(n6872[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n6551[0]), .I2(n147_adj_4032), 
            .I3(n22683), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_14 (.CI(n22959), .I0(n6895[11]), .I1(n956), .CO(n22960));
    SB_CARRY mult_10_add_1225_3 (.CI(n22683), .I0(n6551[0]), .I1(n147_adj_4032), 
            .CO(n22684));
    SB_LUT4 add_3400_13_lut (.I0(GND_net), .I1(n6895[10]), .I2(n883), 
            .I3(n22958), .O(n6872[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3492[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_13 (.CI(n22958), .I0(n6895[10]), .I1(n883), .CO(n22959));
    SB_LUT4 add_3400_12_lut (.I0(GND_net), .I1(n6895[9]), .I2(n810), .I3(n22957), 
            .O(n6872[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_12 (.CI(n22957), .I0(n6895[9]), .I1(n810), .CO(n22958));
    SB_LUT4 add_3400_11_lut (.I0(GND_net), .I1(n6895[8]), .I2(n737), .I3(n22956), 
            .O(n6872[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1449 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3392 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3392 [22]), .O(n13_adj_4254));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut_adj_1449.LUT_INIT = 16'h6ca0;
    SB_CARRY add_3400_11 (.CI(n22956), .I0(n6895[8]), .I1(n737), .CO(n22957));
    SB_LUT4 add_3400_10_lut (.I0(GND_net), .I1(n6895[7]), .I2(n664), .I3(n22955), 
            .O(n6872[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_10 (.CI(n22955), .I0(n6895[7]), .I1(n664), .CO(n22956));
    SB_LUT4 add_3400_9_lut (.I0(GND_net), .I1(n6895[6]), .I2(n591), .I3(n22954), 
            .O(n6872[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_9 (.CI(n22954), .I0(n6895[6]), .I1(n591), .CO(n22955));
    SB_LUT4 add_3400_8_lut (.I0(GND_net), .I1(n6895[5]), .I2(n518), .I3(n22953), 
            .O(n6872[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_8 (.CI(n22953), .I0(n6895[5]), .I1(n518), .CO(n22954));
    SB_LUT4 add_3400_7_lut (.I0(GND_net), .I1(n6895[4]), .I2(n445), .I3(n22952), 
            .O(n6872[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1450 (.I0(n13_adj_4254), .I1(n18_adj_4253), .I2(n21886), 
            .I3(n4_adj_4255), .O(n27839));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_CARRY add_3400_7 (.CI(n22952), .I0(n6895[4]), .I1(n445), .CO(n22953));
    SB_LUT4 add_3400_6_lut (.I0(GND_net), .I1(n6895[3]), .I2(n372), .I3(n22951), 
            .O(n6872[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_6 (.CI(n22951), .I0(n6895[3]), .I1(n372), .CO(n22952));
    SB_LUT4 i24714_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n30983), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4145), .O(n29780));
    defparam i24714_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_33_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n30952));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24702_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n30952), 
            .I2(IntegralLimit[14]), .I3(n29780), .O(n29768));
    defparam i24702_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_28_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n30947));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_28_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4256));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24446_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n29510));
    defparam i24446_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_51_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n30970));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_51_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4257));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4031), .I2(n74_adj_4030), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4256), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4258));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4031), .I1(n74_adj_4030), 
            .CO(n22683));
    SB_LUT4 add_3400_5_lut (.I0(GND_net), .I1(n6895[2]), .I2(n299), .I3(n22950), 
            .O(n6872[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_5 (.CI(n22950), .I0(n6895[2]), .I1(n299), .CO(n22951));
    SB_LUT4 i24895_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n30965), 
            .I2(IntegralLimit[11]), .I3(n29778), .O(n29961));
    defparam i24895_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_3377_23_lut (.I0(GND_net), .I1(n6575[20]), .I2(GND_net), 
            .I3(n22682), .O(n6551[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_22_lut (.I0(GND_net), .I1(n6575[19]), .I2(GND_net), 
            .I3(n22681), .O(n6551[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24454_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n30959), 
            .I2(IntegralLimit[13]), .I3(n29961), .O(n29518));
    defparam i24454_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_3400_4_lut (.I0(GND_net), .I1(n6895[1]), .I2(n226), .I3(n22949), 
            .O(n6872[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_31_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n30950));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3400_4 (.CI(n22949), .I0(n6895[1]), .I1(n226), .CO(n22950));
    SB_LUT4 add_3400_3_lut (.I0(GND_net), .I1(n6895[0]), .I2(n153), .I3(n22948), 
            .O(n6872[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_3 (.CI(n22948), .I0(n6895[0]), .I1(n153), .CO(n22949));
    SB_LUT4 add_3400_2_lut (.I0(GND_net), .I1(n11_adj_4029), .I2(n80), 
            .I3(GND_net), .O(n6872[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_2 (.CI(GND_net), .I0(n11_adj_4029), .I1(n80), .CO(n22948));
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n22006));
    SB_CARRY add_560_4 (.CI(n21946), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n2552[2]), .CO(n21947));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3392 [23]), 
            .I1(n6848[21]), .I2(GND_net), .I3(n22947), .O(n5002[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24823_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n30950), 
            .I2(IntegralLimit[15]), .I3(n29518), .O(n29889));
    defparam i24823_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_57_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n30976));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_57_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24974_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n30976), 
            .I2(IntegralLimit[17]), .I3(n29889), .O(n30040));
    defparam i24974_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n6848[20]), .I2(GND_net), 
            .I3(n22946), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n22946), .I0(n6848[20]), .I1(GND_net), 
            .CO(n22947));
    SB_CARRY add_3377_22 (.CI(n22681), .I0(n6575[19]), .I1(GND_net), .CO(n22682));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n6848[19]), .I2(GND_net), 
            .I3(n22945), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n22945), .I0(n6848[19]), .I1(GND_net), 
            .CO(n22946));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n6848[18]), .I2(GND_net), 
            .I3(n22944), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n22944), .I0(n6848[18]), .I1(GND_net), 
            .CO(n22945));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n22206), .I0(GND_net), .I1(n1_adj_4303[15]), 
            .CO(n22207));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n6848[17]), .I2(GND_net), 
            .I3(n22943), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4303[14]), .I3(n22205), .O(n29_adj_4250)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_560_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n2552[1]), .I3(n21945), .O(\PID_CONTROLLER.integral_23__N_3392 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n22943), .I0(n6848[17]), .I1(GND_net), 
            .CO(n22944));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n6848[16]), .I2(GND_net), 
            .I3(n22942), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_21_lut (.I0(GND_net), .I1(n6575[18]), .I2(GND_net), 
            .I3(n22680), .O(n6551[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_21 (.CI(n22680), .I0(n6575[18]), .I1(GND_net), .CO(n22681));
    SB_LUT4 add_3377_20_lut (.I0(GND_net), .I1(n6575[17]), .I2(GND_net), 
            .I3(n22679), .O(n6551[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_20 (.CI(n22679), .I0(n6575[17]), .I1(GND_net), .CO(n22680));
    SB_LUT4 add_3377_19_lut (.I0(GND_net), .I1(n6575[16]), .I2(GND_net), 
            .I3(n22678), .O(n6551[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_19 (.CI(n22678), .I0(n6575[16]), .I1(GND_net), .CO(n22679));
    SB_LUT4 add_3377_18_lut (.I0(GND_net), .I1(n6575[15]), .I2(GND_net), 
            .I3(n22677), .O(n6551[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n22205), .I0(GND_net), .I1(n1_adj_4303[14]), 
            .CO(n22206));
    SB_CARRY mult_11_add_1225_19 (.CI(n22942), .I0(n6848[16]), .I1(GND_net), 
            .CO(n22943));
    SB_CARRY add_3377_18 (.CI(n22677), .I0(n6575[15]), .I1(GND_net), .CO(n22678));
    SB_LUT4 add_3377_17_lut (.I0(GND_net), .I1(n6575[14]), .I2(GND_net), 
            .I3(n22676), .O(n6551[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_17 (.CI(n22676), .I0(n6575[14]), .I1(GND_net), .CO(n22677));
    SB_LUT4 add_3377_16_lut (.I0(GND_net), .I1(n6575[13]), .I2(n1099_adj_4027), 
            .I3(n22675), .O(n6551[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_16 (.CI(n22675), .I0(n6575[13]), .I1(n1099_adj_4027), 
            .CO(n22676));
    SB_LUT4 add_3377_15_lut (.I0(GND_net), .I1(n6575[12]), .I2(n1026_adj_4026), 
            .I3(n22674), .O(n6551[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_15 (.CI(n22674), .I0(n6575[12]), .I1(n1026_adj_4026), 
            .CO(n22675));
    SB_LUT4 add_3377_14_lut (.I0(GND_net), .I1(n6575[11]), .I2(n953_adj_4025), 
            .I3(n22673), .O(n6551[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_14 (.CI(n22673), .I0(n6575[11]), .I1(n953_adj_4025), 
            .CO(n22674));
    SB_LUT4 add_3377_13_lut (.I0(GND_net), .I1(n6575[10]), .I2(n880_adj_4024), 
            .I3(n22672), .O(n6551[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_13 (.CI(n22672), .I0(n6575[10]), .I1(n880_adj_4024), 
            .CO(n22673));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n6848[15]), .I2(GND_net), 
            .I3(n22941), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_3 (.CI(n21945), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n2552[1]), .CO(n21946));
    SB_CARRY mult_11_add_1225_18 (.CI(n22941), .I0(n6848[15]), .I1(GND_net), 
            .CO(n22942));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n6848[14]), .I2(GND_net), 
            .I3(n22940), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_12_lut (.I0(GND_net), .I1(n6575[9]), .I2(n807_adj_4023), 
            .I3(n22671), .O(n6551[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n22940), .I0(n6848[14]), .I1(GND_net), 
            .CO(n22941));
    SB_CARRY add_3377_12 (.CI(n22671), .I0(n6575[9]), .I1(n807_adj_4023), 
            .CO(n22672));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n6848[13]), .I2(n1096), 
            .I3(n22939), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n22939), .I0(n6848[13]), .I1(n1096), 
            .CO(n22940));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n6848[12]), .I2(n1023), 
            .I3(n22938), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_11_lut (.I0(GND_net), .I1(n6575[8]), .I2(n734_adj_4022), 
            .I3(n22670), .O(n6551[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_11 (.CI(n22670), .I0(n6575[8]), .I1(n734_adj_4022), 
            .CO(n22671));
    SB_LUT4 add_3377_10_lut (.I0(GND_net), .I1(n6575[7]), .I2(n661_adj_4021), 
            .I3(n22669), .O(n6551[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n22938), .I0(n6848[12]), .I1(n1023), 
            .CO(n22939));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n6848[11]), .I2(n950), 
            .I3(n22937), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n22937), .I0(n6848[11]), .I1(n950), 
            .CO(n22938));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4303[13]), .I3(n22204), .O(n27_adj_4226)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n6848[10]), .I2(n877), 
            .I3(n22936), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_10 (.CI(n22669), .I0(n6575[7]), .I1(n661_adj_4021), 
            .CO(n22670));
    SB_LUT4 add_3377_9_lut (.I0(GND_net), .I1(n6575[6]), .I2(n588_adj_4019), 
            .I3(n22668), .O(n6551[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_9 (.CI(n22668), .I0(n6575[6]), .I1(n588_adj_4019), 
            .CO(n22669));
    SB_CARRY mult_11_add_1225_13 (.CI(n22936), .I0(n6848[10]), .I1(n877), 
            .CO(n22937));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n22204), .I0(GND_net), .I1(n1_adj_4303[13]), 
            .CO(n22205));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4303[12]), .I3(n22203), .O(n25_adj_4247)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n22203), .I0(GND_net), .I1(n1_adj_4303[12]), 
            .CO(n22204));
    SB_LUT4 add_560_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n2552[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3392 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_8_lut (.I0(GND_net), .I1(n6575[5]), .I2(n515_adj_4017), 
            .I3(n22667), .O(n6551[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_8 (.CI(n22667), .I0(n6575[5]), .I1(n515_adj_4017), 
            .CO(n22668));
    SB_LUT4 add_3377_7_lut (.I0(GND_net), .I1(n6575[4]), .I2(n442_adj_4016), 
            .I3(n22666), .O(n6551[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_7 (.CI(n22666), .I0(n6575[4]), .I1(n442_adj_4016), 
            .CO(n22667));
    SB_LUT4 add_3377_6_lut (.I0(GND_net), .I1(n6575[3]), .I2(n369_adj_4015), 
            .I3(n22665), .O(n6551[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_6 (.CI(n22665), .I0(n6575[3]), .I1(n369_adj_4015), 
            .CO(n22666));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n6848[9]), .I2(n804), 
            .I3(n22935), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_5_lut (.I0(GND_net), .I1(n6575[2]), .I2(n296_adj_4013), 
            .I3(n22664), .O(n6551[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n22935), .I0(n6848[9]), .I1(n804), 
            .CO(n22936));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n6848[8]), .I2(n731), 
            .I3(n22934), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n22934), .I0(n6848[8]), .I1(n731), 
            .CO(n22935));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n6848[7]), .I2(n658), 
            .I3(n22933), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n22933), .I0(n6848[7]), .I1(n658), 
            .CO(n22934));
    SB_CARRY add_3377_5 (.CI(n22664), .I0(n6575[2]), .I1(n296_adj_4013), 
            .CO(n22665));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n6848[6]), .I2(n585), 
            .I3(n22932), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n22932), .I0(n6848[6]), .I1(n585), 
            .CO(n22933));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n6848[5]), .I2(n512), 
            .I3(n22931), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n22931), .I0(n6848[5]), .I1(n512), 
            .CO(n22932));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n6848[4]), .I2(n439), 
            .I3(n22930), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n22930), .I0(n6848[4]), .I1(n439), 
            .CO(n22931));
    SB_CARRY add_560_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n2552[0]), .CO(n21945));
    SB_LUT4 add_3377_4_lut (.I0(GND_net), .I1(n6575[1]), .I2(n223_adj_4012), 
            .I3(n22663), .O(n6551[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4303[11]), .I3(n22202), .O(n23_adj_4248)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n6848[3]), .I2(n366), 
            .I3(n22929), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n22929), .I0(n6848[3]), .I1(n366), 
            .CO(n22930));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n6848[2]), .I2(n293), 
            .I3(n22928), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n22928), .I0(n6848[2]), .I1(n293), 
            .CO(n22929));
    SB_CARRY add_3377_4 (.CI(n22663), .I0(n6575[1]), .I1(n223_adj_4012), 
            .CO(n22664));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n6848[1]), .I2(n220), 
            .I3(n22927), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n22927), .I0(n6848[1]), .I1(n220), 
            .CO(n22928));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n6848[0]), .I2(n147_adj_4010), 
            .I3(n22926), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n22926), .I0(n6848[0]), .I1(n147_adj_4010), 
            .CO(n22927));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4009), .I2(n74), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4009), .I1(n74), 
            .CO(n22926));
    SB_LUT4 add_3399_23_lut (.I0(GND_net), .I1(n6872[20]), .I2(GND_net), 
            .I3(n22925), .O(n6848[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_3_lut (.I0(GND_net), .I1(n6575[0]), .I2(n150_adj_4008), 
            .I3(n22662), .O(n6551[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3399_22_lut (.I0(GND_net), .I1(n6872[19]), .I2(GND_net), 
            .I3(n22924), .O(n6848[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_22 (.CI(n22924), .I0(n6872[19]), .I1(GND_net), .CO(n22925));
    SB_LUT4 add_3399_21_lut (.I0(GND_net), .I1(n6872[18]), .I2(GND_net), 
            .I3(n22923), .O(n6848[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_21 (.CI(n22923), .I0(n6872[18]), .I1(GND_net), .CO(n22924));
    SB_LUT4 add_3399_20_lut (.I0(GND_net), .I1(n6872[17]), .I2(GND_net), 
            .I3(n22922), .O(n6848[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_20 (.CI(n22922), .I0(n6872[17]), .I1(GND_net), .CO(n22923));
    SB_LUT4 add_3399_19_lut (.I0(GND_net), .I1(n6872[16]), .I2(GND_net), 
            .I3(n22921), .O(n6848[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_19 (.CI(n22921), .I0(n6872[16]), .I1(GND_net), .CO(n22922));
    SB_LUT4 add_3399_18_lut (.I0(GND_net), .I1(n6872[15]), .I2(GND_net), 
            .I3(n22920), .O(n6848[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_3 (.CI(n22662), .I0(n6575[0]), .I1(n150_adj_4008), 
            .CO(n22663));
    SB_CARRY add_3399_18 (.CI(n22920), .I0(n6872[15]), .I1(GND_net), .CO(n22921));
    SB_LUT4 add_3399_17_lut (.I0(GND_net), .I1(n6872[14]), .I2(GND_net), 
            .I3(n22919), .O(n6848[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_17 (.CI(n22919), .I0(n6872[14]), .I1(GND_net), .CO(n22920));
    SB_LUT4 add_3377_2_lut (.I0(GND_net), .I1(n8_adj_4007), .I2(n77_adj_4005), 
            .I3(GND_net), .O(n6551[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3399_16_lut (.I0(GND_net), .I1(n6872[13]), .I2(n1099), 
            .I3(n22918), .O(n6848[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_2 (.CI(GND_net), .I0(n8_adj_4007), .I1(n77_adj_4005), 
            .CO(n22662));
    SB_CARRY add_3399_16 (.CI(n22918), .I0(n6872[13]), .I1(n1099), .CO(n22919));
    SB_LUT4 add_3399_15_lut (.I0(GND_net), .I1(n6872[12]), .I2(n1026), 
            .I3(n22917), .O(n6848[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_22_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n30941));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_22_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25028_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n30941), 
            .I2(IntegralLimit[19]), .I3(n30040), .O(n30094));
    defparam i25028_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_19_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n30938));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4263));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24435_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n29498));
    defparam i24435_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_3399_15 (.CI(n22917), .I0(n6872[12]), .I1(n1026), .CO(n22918));
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4263), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4264));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3399_14_lut (.I0(GND_net), .I1(n6872[11]), .I2(n953), 
            .I3(n22916), .O(n6848[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4265));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3399_14 (.CI(n22916), .I0(n6872[11]), .I1(n953), .CO(n22917));
    SB_LUT4 i24843_3_lut (.I0(n6_adj_4265), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n29909));   // verilog/motorControl.v(31[10:34])
    defparam i24843_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3399_13_lut (.I0(GND_net), .I1(n6872[10]), .I2(n880), 
            .I3(n22915), .O(n6848[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24844_3_lut (.I0(n29909), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n29910));   // verilog/motorControl.v(31[10:34])
    defparam i24844_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3399_13 (.CI(n22915), .I0(n6872[10]), .I1(n880), .CO(n22916));
    SB_LUT4 i24437_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n30959), 
            .I2(IntegralLimit[21]), .I3(n29774), .O(n29500));
    defparam i24437_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_3399_12_lut (.I0(GND_net), .I1(n6872[9]), .I2(n807), .I3(n22914), 
            .O(n6848[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_12 (.CI(n22914), .I0(n6872[9]), .I1(n807), .CO(n22915));
    SB_LUT4 i24799_4_lut (.I0(n24_adj_4264), .I1(n8_adj_4266), .I2(n30936), 
            .I3(n29498), .O(n29865));   // verilog/motorControl.v(31[10:34])
    defparam i24799_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3399_11_lut (.I0(GND_net), .I1(n6872[8]), .I2(n734), .I3(n22913), 
            .O(n6848[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24656_3_lut (.I0(n29910), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n29722));   // verilog/motorControl.v(31[10:34])
    defparam i24656_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3399_11 (.CI(n22913), .I0(n6872[8]), .I1(n734), .CO(n22914));
    SB_LUT4 add_3399_10_lut (.I0(GND_net), .I1(n6872[7]), .I2(n661), .I3(n22912), 
            .O(n6848[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_10 (.CI(n22912), .I0(n6872[7]), .I1(n661), .CO(n22913));
    SB_LUT4 add_3399_9_lut (.I0(GND_net), .I1(n6872[6]), .I2(n588), .I3(n22911), 
            .O(n6848[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_9 (.CI(n22911), .I0(n6872[6]), .I1(n588), .CO(n22912));
    SB_LUT4 add_3399_8_lut (.I0(GND_net), .I1(n6872[5]), .I2(n515), .I3(n22910), 
            .O(n6848[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_8 (.CI(n22910), .I0(n6872[5]), .I1(n515), .CO(n22911));
    SB_LUT4 add_3399_7_lut (.I0(GND_net), .I1(n6872[4]), .I2(n442), .I3(n22909), 
            .O(n6848[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_7 (.CI(n22909), .I0(n6872[4]), .I1(n442), .CO(n22910));
    SB_LUT4 add_3399_6_lut (.I0(GND_net), .I1(n6872[3]), .I2(n369), .I3(n22908), 
            .O(n6848[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_6 (.CI(n22908), .I0(n6872[3]), .I1(n369), .CO(n22909));
    SB_LUT4 add_3399_5_lut (.I0(GND_net), .I1(n6872[2]), .I2(n296), .I3(n22907), 
            .O(n6848[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_5 (.CI(n22907), .I0(n6872[2]), .I1(n296), .CO(n22908));
    SB_LUT4 add_3399_4_lut (.I0(GND_net), .I1(n6872[1]), .I2(n223), .I3(n22906), 
            .O(n6848[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_4 (.CI(n22906), .I0(n6872[1]), .I1(n223), .CO(n22907));
    SB_LUT4 add_3399_3_lut (.I0(GND_net), .I1(n6872[0]), .I2(n150), .I3(n22905), 
            .O(n6848[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_3 (.CI(n22905), .I0(n6872[0]), .I1(n150), .CO(n22906));
    SB_LUT4 add_3399_2_lut (.I0(GND_net), .I1(n8_adj_4002), .I2(n77), 
            .I3(GND_net), .O(n6848[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n22202), .I0(GND_net), .I1(n1_adj_4303[11]), 
            .CO(n22203));
    SB_CARRY add_3399_2 (.CI(GND_net), .I0(n8_adj_4002), .I1(n77), .CO(n22905));
    SB_LUT4 add_3393_7_lut (.I0(GND_net), .I1(n27634), .I2(n490_adj_3992), 
            .I3(n22904), .O(n6815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3393_6_lut (.I0(GND_net), .I1(n6823[3]), .I2(n417_adj_3960), 
            .I3(n22903), .O(n6815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_6 (.CI(n22903), .I0(n6823[3]), .I1(n417_adj_3960), 
            .CO(n22904));
    SB_LUT4 add_3393_5_lut (.I0(GND_net), .I1(n6823[2]), .I2(n344_adj_3940), 
            .I3(n22902), .O(n6815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_5 (.CI(n22902), .I0(n6823[2]), .I1(n344_adj_3940), 
            .CO(n22903));
    SB_LUT4 add_3393_4_lut (.I0(GND_net), .I1(n6823[1]), .I2(n271_adj_3925), 
            .I3(n22901), .O(n6815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_4 (.CI(n22901), .I0(n6823[1]), .I1(n271_adj_3925), 
            .CO(n22902));
    SB_LUT4 add_3393_3_lut (.I0(GND_net), .I1(n6823[0]), .I2(n198_adj_3921), 
            .I3(n22900), .O(n6815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_3 (.CI(n22900), .I0(n6823[0]), .I1(n198_adj_3921), 
            .CO(n22901));
    SB_LUT4 add_3393_2_lut (.I0(GND_net), .I1(n56_adj_3918), .I2(n125_adj_3907), 
            .I3(GND_net), .O(n6815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_2 (.CI(GND_net), .I0(n56_adj_3918), .I1(n125_adj_3907), 
            .CO(n22900));
    SB_LUT4 add_3392_8_lut (.I0(GND_net), .I1(n6815[5]), .I2(n560_adj_3902), 
            .I3(n22899), .O(n6806[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3392_7_lut (.I0(GND_net), .I1(n6815[4]), .I2(n487_adj_3898), 
            .I3(n22898), .O(n6806[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4303[10]), .I3(n22201), .O(n21_adj_4230)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3392_7 (.CI(n22898), .I0(n6815[4]), .I1(n487_adj_3898), 
            .CO(n22899));
    SB_LUT4 add_3392_6_lut (.I0(GND_net), .I1(n6815[3]), .I2(n414), .I3(n22897), 
            .O(n6806[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_6 (.CI(n22897), .I0(n6815[3]), .I1(n414), .CO(n22898));
    SB_LUT4 add_3392_5_lut (.I0(GND_net), .I1(n6815[2]), .I2(n341), .I3(n22896), 
            .O(n6806[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_5 (.CI(n22896), .I0(n6815[2]), .I1(n341), .CO(n22897));
    SB_LUT4 add_560_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n2552[6]), .I3(n21950), .O(\PID_CONTROLLER.integral_23__N_3392 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3443 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4267), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4268));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i24942_3_lut (.I0(n4_adj_4268), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27_adj_4226), .I3(GND_net), .O(n30008));   // verilog/motorControl.v(31[38:63])
    defparam i24942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24943_3_lut (.I0(n30008), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4250), .I3(GND_net), .O(n30009));   // verilog/motorControl.v(31[38:63])
    defparam i24943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_4251), .I3(GND_net), 
            .O(n12_adj_4269));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24384_2_lut (.I0(n33_adj_4251), .I1(n15_adj_4227), .I2(GND_net), 
            .I3(GND_net), .O(n29447));
    defparam i24384_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4228), .I3(GND_net), 
            .O(n10_adj_4270));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4269), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4236), .I3(GND_net), 
            .O(n30_adj_4271));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24386_4_lut (.I0(n33_adj_4251), .I1(n31_adj_4249), .I2(n29_adj_4250), 
            .I3(n29455), .O(n29449));
    defparam i24386_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i25002_4_lut (.I0(n30_adj_4271), .I1(n10_adj_4270), .I2(n35_adj_4236), 
            .I3(n29447), .O(n30068));   // verilog/motorControl.v(31[38:63])
    defparam i25002_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24864_3_lut (.I0(n30009), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_4249), .I3(GND_net), .O(n29930));   // verilog/motorControl.v(31[38:63])
    defparam i24864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25051_4_lut (.I0(n29930), .I1(n30068), .I2(n35_adj_4236), 
            .I3(n29449), .O(n30117));   // verilog/motorControl.v(31[38:63])
    defparam i25051_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25052_3_lut (.I0(n30117), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_4224), .I3(GND_net), .O(n30118));   // verilog/motorControl.v(31[38:63])
    defparam i25052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25037_3_lut (.I0(n30118), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_4222), .I3(GND_net), .O(n30103));   // verilog/motorControl.v(31[38:63])
    defparam i25037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4245), .I3(GND_net), 
            .O(n6_adj_4272));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_3392_4_lut (.I0(GND_net), .I1(n6815[1]), .I2(n268), .I3(n22895), 
            .O(n6806[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_4 (.CI(n22895), .I0(n6815[1]), .I1(n268), .CO(n22896));
    SB_LUT4 add_3392_3_lut (.I0(GND_net), .I1(n6815[0]), .I2(n195_adj_3888), 
            .I3(n22894), .O(n6806[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_3 (.CI(n22894), .I0(n6815[0]), .I1(n195_adj_3888), 
            .CO(n22895));
    SB_LUT4 add_3392_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n6806[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n22894));
    SB_LUT4 add_3391_9_lut (.I0(GND_net), .I1(n6806[6]), .I2(n630), .I3(n22893), 
            .O(n6796[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3391_8_lut (.I0(GND_net), .I1(n6806[5]), .I2(n557), .I3(n22892), 
            .O(n6796[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4179));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3391_8 (.CI(n22892), .I0(n6806[5]), .I1(n557), .CO(n22893));
    SB_LUT4 add_3391_7_lut (.I0(GND_net), .I1(n6806[4]), .I2(n484), .I3(n22891), 
            .O(n6796[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_7 (.CI(n22891), .I0(n6806[4]), .I1(n484), .CO(n22892));
    SB_LUT4 add_3391_6_lut (.I0(GND_net), .I1(n6806[3]), .I2(n411), .I3(n22890), 
            .O(n6796[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_6 (.CI(n22890), .I0(n6806[3]), .I1(n411), .CO(n22891));
    SB_LUT4 add_3391_5_lut (.I0(GND_net), .I1(n6806[2]), .I2(n338), .I3(n22889), 
            .O(n6796[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_5 (.CI(n22889), .I0(n6806[2]), .I1(n338), .CO(n22890));
    SB_LUT4 add_3391_4_lut (.I0(GND_net), .I1(n6806[1]), .I2(n265), .I3(n22888), 
            .O(n6796[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_4 (.CI(n22888), .I0(n6806[1]), .I1(n265), .CO(n22889));
    SB_LUT4 add_3391_3_lut (.I0(GND_net), .I1(n6806[0]), .I2(n192), .I3(n22887), 
            .O(n6796[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_3 (.CI(n22887), .I0(n6806[0]), .I1(n192), .CO(n22888));
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4303[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4178));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15184_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15184_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3391_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n6796[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n22887));
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4176));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4175));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_10_lut (.I0(GND_net), .I1(n6796[7]), .I2(n700), .I3(n22886), 
            .O(n6785[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4173));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_9_lut (.I0(GND_net), .I1(n6796[6]), .I2(n627), .I3(n22885), 
            .O(n6785[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_9 (.CI(n22885), .I0(n6796[6]), .I1(n627), .CO(n22886));
    SB_LUT4 add_3390_8_lut (.I0(GND_net), .I1(n6796[5]), .I2(n554), .I3(n22884), 
            .O(n6785[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_8 (.CI(n22884), .I0(n6796[5]), .I1(n554), .CO(n22885));
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4169));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4163));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_7_lut (.I0(GND_net), .I1(n6796[4]), .I2(n481), .I3(n22883), 
            .O(n6785[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_7 (.CI(n22883), .I0(n6796[4]), .I1(n481), .CO(n22884));
    SB_LUT4 add_3390_6_lut (.I0(GND_net), .I1(n6796[3]), .I2(n408), .I3(n22882), 
            .O(n6785[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_6 (.CI(n22882), .I0(n6796[3]), .I1(n408), .CO(n22883));
    SB_LUT4 add_3390_5_lut (.I0(GND_net), .I1(n6796[2]), .I2(n335), .I3(n22881), 
            .O(n6785[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4157));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3390_5 (.CI(n22881), .I0(n6796[2]), .I1(n335), .CO(n22882));
    SB_LUT4 add_3390_4_lut (.I0(GND_net), .I1(n6796[1]), .I2(n262), .I3(n22880), 
            .O(n6785[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_4 (.CI(n22880), .I0(n6796[1]), .I1(n262), .CO(n22881));
    SB_LUT4 add_3390_3_lut (.I0(GND_net), .I1(n6796[0]), .I2(n189), .I3(n22879), 
            .O(n6785[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_3 (.CI(n22879), .I0(n6796[0]), .I1(n189), .CO(n22880));
    SB_LUT4 add_3390_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n6785[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n22879));
    SB_LUT4 add_3389_11_lut (.I0(GND_net), .I1(n6785[8]), .I2(n770), .I3(n22878), 
            .O(n6773[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_10_lut (.I0(GND_net), .I1(n6785[7]), .I2(n697), .I3(n22877), 
            .O(n6773[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_10 (.CI(n22877), .I0(n6785[7]), .I1(n697), .CO(n22878));
    SB_LUT4 add_3389_9_lut (.I0(GND_net), .I1(n6785[6]), .I2(n624), .I3(n22876), 
            .O(n6773[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_9 (.CI(n22876), .I0(n6785[6]), .I1(n624), .CO(n22877));
    SB_LUT4 add_3389_8_lut (.I0(GND_net), .I1(n6785[5]), .I2(n551), .I3(n22875), 
            .O(n6773[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_8 (.CI(n22875), .I0(n6785[5]), .I1(n551), .CO(n22876));
    SB_LUT4 add_3389_7_lut (.I0(GND_net), .I1(n6785[4]), .I2(n478), .I3(n22874), 
            .O(n6773[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_7 (.CI(n22874), .I0(n6785[4]), .I1(n478), .CO(n22875));
    SB_LUT4 add_3389_6_lut (.I0(GND_net), .I1(n6785[3]), .I2(n405), .I3(n22873), 
            .O(n6773[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_6 (.CI(n22873), .I0(n6785[3]), .I1(n405), .CO(n22874));
    SB_LUT4 add_3389_5_lut (.I0(GND_net), .I1(n6785[2]), .I2(n332), .I3(n22872), 
            .O(n6773[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_5 (.CI(n22872), .I0(n6785[2]), .I1(n332), .CO(n22873));
    SB_LUT4 add_3389_4_lut (.I0(GND_net), .I1(n6785[1]), .I2(n259), .I3(n22871), 
            .O(n6773[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_4 (.CI(n22871), .I0(n6785[1]), .I1(n259), .CO(n22872));
    SB_LUT4 add_3389_3_lut (.I0(GND_net), .I1(n6785[0]), .I2(n186), .I3(n22870), 
            .O(n6773[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_3 (.CI(n22870), .I0(n6785[0]), .I1(n186), .CO(n22871));
    SB_LUT4 add_3389_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n6773[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n22870));
    SB_LUT4 add_3388_12_lut (.I0(GND_net), .I1(n6773[9]), .I2(n840), .I3(n22869), 
            .O(n6760[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3388_11_lut (.I0(GND_net), .I1(n6773[8]), .I2(n767), .I3(n22868), 
            .O(n6760[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_11 (.CI(n22868), .I0(n6773[8]), .I1(n767), .CO(n22869));
    SB_LUT4 add_3388_10_lut (.I0(GND_net), .I1(n6773[7]), .I2(n694), .I3(n22867), 
            .O(n6760[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_10 (.CI(n22867), .I0(n6773[7]), .I1(n694), .CO(n22868));
    SB_LUT4 add_3388_9_lut (.I0(GND_net), .I1(n6773[6]), .I2(n621), .I3(n22866), 
            .O(n6760[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_9 (.CI(n22866), .I0(n6773[6]), .I1(n621), .CO(n22867));
    SB_LUT4 add_3388_8_lut (.I0(GND_net), .I1(n6773[5]), .I2(n548), .I3(n22865), 
            .O(n6760[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_8 (.CI(n22865), .I0(n6773[5]), .I1(n548), .CO(n22866));
    SB_LUT4 add_3388_7_lut (.I0(GND_net), .I1(n6773[4]), .I2(n475), .I3(n22864), 
            .O(n6760[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_7 (.CI(n22864), .I0(n6773[4]), .I1(n475), .CO(n22865));
    SB_LUT4 add_3388_6_lut (.I0(GND_net), .I1(n6773[3]), .I2(n402), .I3(n22863), 
            .O(n6760[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_6 (.CI(n22863), .I0(n6773[3]), .I1(n402), .CO(n22864));
    SB_LUT4 add_3388_5_lut (.I0(GND_net), .I1(n6773[2]), .I2(n329), .I3(n22862), 
            .O(n6760[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_5 (.CI(n22862), .I0(n6773[2]), .I1(n329), .CO(n22863));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n22201), .I0(GND_net), .I1(n1_adj_4303[10]), 
            .CO(n22202));
    SB_LUT4 i24835_3_lut (.I0(n6_adj_4272), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4230), .I3(GND_net), .O(n29901));   // verilog/motorControl.v(31[38:63])
    defparam i24835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24836_3_lut (.I0(n29901), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4248), .I3(GND_net), .O(n29902));   // verilog/motorControl.v(31[38:63])
    defparam i24836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24376_4_lut (.I0(n43_adj_4197), .I1(n25_adj_4247), .I2(n23_adj_4248), 
            .I3(n29464), .O(n29439));
    defparam i24376_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24801_4_lut (.I0(n24_adj_4237), .I1(n8_adj_4235), .I2(n45_adj_4181), 
            .I3(n29437), .O(n29867));   // verilog/motorControl.v(31[38:63])
    defparam i24801_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24666_3_lut (.I0(n29902), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4247), .I3(GND_net), .O(n29732));   // verilog/motorControl.v(31[38:63])
    defparam i24666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24378_4_lut (.I0(n43_adj_4197), .I1(n41_adj_4215), .I2(n39_adj_4222), 
            .I3(n30062), .O(n29441));
    defparam i24378_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24952_4_lut (.I0(n29732), .I1(n29867), .I2(n45_adj_4181), 
            .I3(n29439), .O(n30018));   // verilog/motorControl.v(31[38:63])
    defparam i24952_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25021_3_lut (.I0(n30103), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4215), .I3(GND_net), .O(n40_adj_4273));   // verilog/motorControl.v(31[38:63])
    defparam i25021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24954_4_lut (.I0(n40_adj_4273), .I1(n30018), .I2(n45_adj_4181), 
            .I3(n29441), .O(n30020));   // verilog/motorControl.v(31[38:63])
    defparam i24954_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4155));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4274));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i24841_3_lut (.I0(n4_adj_4274), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n29907));   // verilog/motorControl.v(31[10:34])
    defparam i24841_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24842_3_lut (.I0(n29907), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n29908));   // verilog/motorControl.v(31[10:34])
    defparam i24842_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24448_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n30947), 
            .I2(IntegralLimit[16]), .I3(n29768), .O(n29512));
    defparam i24448_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i15185_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15185_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15189_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15189_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_4_lut (.I0(GND_net), .I1(n6773[1]), .I2(n256), .I3(n22861), 
            .O(n6760[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_4 (.CI(n22861), .I0(n6773[1]), .I1(n256), .CO(n22862));
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4148));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_3_lut (.I0(GND_net), .I1(n6773[0]), .I2(n183), .I3(n22860), 
            .O(n6760[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_3 (.CI(n22860), .I0(n6773[0]), .I1(n183), .CO(n22861));
    SB_LUT4 add_3388_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n6760[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n22860));
    SB_LUT4 add_3387_13_lut (.I0(GND_net), .I1(n6760[10]), .I2(n910), 
            .I3(n22859), .O(n6746[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_12_lut (.I0(GND_net), .I1(n6760[9]), .I2(n837), .I3(n22858), 
            .O(n6746[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_12 (.CI(n22858), .I0(n6760[9]), .I1(n837), .CO(n22859));
    SB_LUT4 add_3387_11_lut (.I0(GND_net), .I1(n6760[8]), .I2(n764), .I3(n22857), 
            .O(n6746[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_11 (.CI(n22857), .I0(n6760[8]), .I1(n764), .CO(n22858));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4303[9]), .I3(n22200), .O(n19_adj_4231)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3387_10_lut (.I0(GND_net), .I1(n6760[7]), .I2(n691), .I3(n22856), 
            .O(n6746[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_10 (.CI(n22856), .I0(n6760[7]), .I1(n691), .CO(n22857));
    SB_LUT4 add_3387_9_lut (.I0(GND_net), .I1(n6760[6]), .I2(n618), .I3(n22855), 
            .O(n6746[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4126));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_9 (.CI(n22855), .I0(n6760[6]), .I1(n618), .CO(n22856));
    SB_LUT4 add_3387_8_lut (.I0(GND_net), .I1(n6760[5]), .I2(n545), .I3(n22854), 
            .O(n6746[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_8 (.CI(n22854), .I0(n6760[5]), .I1(n545), .CO(n22855));
    SB_LUT4 add_3387_7_lut (.I0(GND_net), .I1(n6760[4]), .I2(n472), .I3(n22853), 
            .O(n6746[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_7 (.CI(n22853), .I0(n6760[4]), .I1(n472), .CO(n22854));
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3387_6_lut (.I0(GND_net), .I1(n6760[3]), .I2(n399), .I3(n22852), 
            .O(n6746[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_6 (.CI(n22852), .I0(n6760[3]), .I1(n399), .CO(n22853));
    SB_LUT4 add_3387_5_lut (.I0(GND_net), .I1(n6760[2]), .I2(n326), .I3(n22851), 
            .O(n6746[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_5 (.CI(n22851), .I0(n6760[2]), .I1(n326), .CO(n22852));
    SB_LUT4 add_3387_4_lut (.I0(GND_net), .I1(n6760[1]), .I2(n253), .I3(n22850), 
            .O(n6746[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_4 (.CI(n22850), .I0(n6760[1]), .I1(n253), .CO(n22851));
    SB_LUT4 add_3387_3_lut (.I0(GND_net), .I1(n6760[0]), .I2(n180), .I3(n22849), 
            .O(n6746[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_3 (.CI(n22849), .I0(n6760[0]), .I1(n180), .CO(n22850));
    SB_LUT4 add_3387_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n6746[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n22849));
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3386_14_lut (.I0(GND_net), .I1(n6746[11]), .I2(n980), 
            .I3(n22848), .O(n6731[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3386_13_lut (.I0(GND_net), .I1(n6746[10]), .I2(n907), 
            .I3(n22847), .O(n6731[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_13 (.CI(n22847), .I0(n6746[10]), .I1(n907), .CO(n22848));
    SB_LUT4 add_3386_12_lut (.I0(GND_net), .I1(n6746[9]), .I2(n834), .I3(n22846), 
            .O(n6731[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_12 (.CI(n22846), .I0(n6746[9]), .I1(n834), .CO(n22847));
    SB_LUT4 add_3386_11_lut (.I0(GND_net), .I1(n6746[8]), .I2(n761), .I3(n22845), 
            .O(n6731[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_11 (.CI(n22845), .I0(n6746[8]), .I1(n761), .CO(n22846));
    SB_LUT4 add_3386_10_lut (.I0(GND_net), .I1(n6746[7]), .I2(n688), .I3(n22844), 
            .O(n6731[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24986_4_lut (.I0(n30_adj_4258), .I1(n10_adj_4257), .I2(n30970), 
            .I3(n29510), .O(n30052));   // verilog/motorControl.v(31[10:34])
    defparam i24986_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24658_3_lut (.I0(n29908), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n29724));   // verilog/motorControl.v(31[10:34])
    defparam i24658_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3386_10 (.CI(n22844), .I0(n6746[7]), .I1(n688), .CO(n22845));
    SB_LUT4 i25038_4_lut (.I0(n29724), .I1(n30052), .I2(n30970), .I3(n29512), 
            .O(n30104));   // verilog/motorControl.v(31[10:34])
    defparam i25038_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25039_3_lut (.I0(n30104), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n30105));   // verilog/motorControl.v(31[10:34])
    defparam i25039_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25013_3_lut (.I0(n30105), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n30079));   // verilog/motorControl.v(31[10:34])
    defparam i25013_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24439_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n30938), 
            .I2(IntegralLimit[21]), .I3(n30094), .O(n29502));
    defparam i24439_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_17_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n30936));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24948_4_lut (.I0(n29722), .I1(n29865), .I2(n30936), .I3(n29500), 
            .O(n30014));   // verilog/motorControl.v(31[10:34])
    defparam i24948_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24664_3_lut (.I0(n30079), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n29730));   // verilog/motorControl.v(31[10:34])
    defparam i24664_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24955_3_lut (.I0(n30020), .I1(\PID_CONTROLLER.integral_23__N_3443 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3442 ));   // verilog/motorControl.v(31[38:63])
    defparam i24955_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24998_4_lut (.I0(n29730), .I1(n30014), .I2(n30936), .I3(n29502), 
            .O(n30064));   // verilog/motorControl.v(31[10:34])
    defparam i24998_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_9_lut (.I0(GND_net), .I1(n6746[6]), .I2(n615), .I3(n22843), 
            .O(n6731[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_9 (.CI(n22843), .I0(n6746[6]), .I1(n615), .CO(n22844));
    SB_LUT4 add_3386_8_lut (.I0(GND_net), .I1(n6746[5]), .I2(n542), .I3(n22842), 
            .O(n6731[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_8 (.CI(n22842), .I0(n6746[5]), .I1(n542), .CO(n22843));
    SB_LUT4 add_3386_7_lut (.I0(GND_net), .I1(n6746[4]), .I2(n469), .I3(n22841), 
            .O(n6731[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_7 (.CI(n22841), .I0(n6746[4]), .I1(n469), .CO(n22842));
    SB_LUT4 add_3386_6_lut (.I0(GND_net), .I1(n6746[3]), .I2(n396), .I3(n22840), 
            .O(n6731[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_6 (.CI(n22840), .I0(n6746[3]), .I1(n396), .CO(n22841));
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_5_lut (.I0(GND_net), .I1(n6746[2]), .I2(n323), .I3(n22839), 
            .O(n6731[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_5 (.CI(n22839), .I0(n6746[2]), .I1(n323), .CO(n22840));
    SB_LUT4 add_3386_4_lut (.I0(GND_net), .I1(n6746[1]), .I2(n250), .I3(n22838), 
            .O(n6731[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n22200), .I0(GND_net), .I1(n1_adj_4303[9]), 
            .CO(n22201));
    SB_CARRY add_3386_4 (.CI(n22838), .I0(n6746[1]), .I1(n250), .CO(n22839));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4303[8]), .I3(n22199), .O(n17_adj_4232)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3386_3_lut (.I0(GND_net), .I1(n6746[0]), .I2(n177), .I3(n22837), 
            .O(n6731[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n22199), .I0(GND_net), .I1(n1_adj_4303[8]), 
            .CO(n22200));
    SB_CARRY add_3386_3 (.CI(n22837), .I0(n6746[0]), .I1(n177), .CO(n22838));
    SB_LUT4 add_3386_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n6731[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n22837));
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4115));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_15_lut (.I0(GND_net), .I1(n6731[12]), .I2(n1050), 
            .I3(n22836), .O(n6715[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3385_14_lut (.I0(GND_net), .I1(n6731[11]), .I2(n977), 
            .I3(n22835), .O(n6715[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_14 (.CI(n22835), .I0(n6731[11]), .I1(n977), .CO(n22836));
    SB_LUT4 add_3385_13_lut (.I0(GND_net), .I1(n6731[10]), .I2(n904), 
            .I3(n22834), .O(n6715[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_830_4_lut  (.I0(n30064), .I1(\PID_CONTROLLER.integral_23__N_3442 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3440 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_830_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4303[7]), .I3(n22198), .O(n15_adj_4227)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n22198), .I0(GND_net), .I1(n1_adj_4303[7]), 
            .CO(n22199));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4303[6]), .I3(n22197), .O(n13_adj_4228)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4112));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4109));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4106));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4095));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4091));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4071));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4014));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4003));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_3991));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_3990));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3988));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3987));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_3986));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_3985));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3385_13 (.CI(n22834), .I0(n6731[10]), .I1(n904), .CO(n22835));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n22197), .I0(GND_net), .I1(n1_adj_4303[6]), 
            .CO(n22198));
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_3983));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4303[5]), .I3(n22196), .O(n11_adj_4229)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n22196), .I0(GND_net), .I1(n1_adj_4303[5]), 
            .CO(n22197));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4303[4]), .I3(n22195), .O(n9_adj_4233)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n22195), .I0(GND_net), .I1(n1_adj_4303[4]), 
            .CO(n22196));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4303[3]), .I3(n22194), .O(n7_adj_4245)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3385_12_lut (.I0(GND_net), .I1(n6731[9]), .I2(n831), .I3(n22833), 
            .O(n6715[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n22194), .I0(GND_net), .I1(n1_adj_4303[3]), 
            .CO(n22195));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4303[2]), .I3(n22193), .O(n5_adj_4246)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n22193), .I0(GND_net), .I1(n1_adj_4303[2]), 
            .CO(n22194));
    SB_CARRY add_3385_12 (.CI(n22833), .I0(n6731[9]), .I1(n831), .CO(n22834));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4303[1]), .I3(n22192), .O(n3_adj_4267)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n22192), .I0(GND_net), .I1(n1_adj_4303[1]), 
            .CO(n22193));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4303[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3443 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4303[0]), 
            .CO(n22192));
    SB_LUT4 i15187_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15187_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n22191), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3385_11_lut (.I0(GND_net), .I1(n6731[8]), .I2(n758), .I3(n22832), 
            .O(n6715[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_11 (.CI(n22832), .I0(n6731[8]), .I1(n758), .CO(n22833));
    SB_LUT4 add_3385_10_lut (.I0(GND_net), .I1(n6731[7]), .I2(n685), .I3(n22831), 
            .O(n6715[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_10 (.CI(n22831), .I0(n6731[7]), .I1(n685), .CO(n22832));
    SB_LUT4 add_3385_9_lut (.I0(GND_net), .I1(n6731[6]), .I2(n612), .I3(n22830), 
            .O(n6715[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n22190), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_9 (.CI(n22830), .I0(n6731[6]), .I1(n612), .CO(n22831));
    SB_LUT4 add_3385_8_lut (.I0(GND_net), .I1(n6731[5]), .I2(n539), .I3(n22829), 
            .O(n6715[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_8 (.CI(n22829), .I0(n6731[5]), .I1(n539), .CO(n22830));
    SB_LUT4 add_3385_7_lut (.I0(GND_net), .I1(n6731[4]), .I2(n466), .I3(n22828), 
            .O(n6715[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_7 (.CI(n22828), .I0(n6731[4]), .I1(n466), .CO(n22829));
    SB_CARRY sub_3_add_2_24 (.CI(n22190), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n22191));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n22189), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_23 (.CI(n22189), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n22190));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n22188), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3385_6_lut (.I0(GND_net), .I1(n6731[3]), .I2(n393), .I3(n22827), 
            .O(n6715[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n22188), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n22189));
    SB_CARRY add_3385_6 (.CI(n22827), .I0(n6731[3]), .I1(n393), .CO(n22828));
    SB_LUT4 add_3385_5_lut (.I0(GND_net), .I1(n6731[2]), .I2(n320), .I3(n22826), 
            .O(n6715[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_3982));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3385_5 (.CI(n22826), .I0(n6731[2]), .I1(n320), .CO(n22827));
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_3981));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_4_lut (.I0(GND_net), .I1(n6731[1]), .I2(n247), .I3(n22825), 
            .O(n6715[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_4 (.CI(n22825), .I0(n6731[1]), .I1(n247), .CO(n22826));
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n22187), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n22187), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n22188));
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n22186), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_3980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_3_lut (.I0(GND_net), .I1(n6731[0]), .I2(n174), .I3(n22824), 
            .O(n6715[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n22186), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n22187));
    SB_CARRY add_3385_3 (.CI(n22824), .I0(n6731[0]), .I1(n174), .CO(n22825));
    SB_LUT4 add_3385_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n6715[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n22824));
    SB_LUT4 add_3384_16_lut (.I0(GND_net), .I1(n6715[13]), .I2(n1120), 
            .I3(n22823), .O(n6698[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3384_15_lut (.I0(GND_net), .I1(n6715[12]), .I2(n1047), 
            .I3(n22822), .O(n6698[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_15 (.CI(n22822), .I0(n6715[12]), .I1(n1047), .CO(n22823));
    SB_LUT4 add_3384_14_lut (.I0(GND_net), .I1(n6715[11]), .I2(n974), 
            .I3(n22821), .O(n6698[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_14 (.CI(n22821), .I0(n6715[11]), .I1(n974), .CO(n22822));
    SB_LUT4 add_3384_13_lut (.I0(GND_net), .I1(n6715[10]), .I2(n901), 
            .I3(n22820), .O(n6698[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_13 (.CI(n22820), .I0(n6715[10]), .I1(n901), .CO(n22821));
    SB_LUT4 add_3384_12_lut (.I0(GND_net), .I1(n6715[9]), .I2(n828), .I3(n22819), 
            .O(n6698[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_12 (.CI(n22819), .I0(n6715[9]), .I1(n828), .CO(n22820));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n22185), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3384_11_lut (.I0(GND_net), .I1(n6715[8]), .I2(n755), .I3(n22818), 
            .O(n6698[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n22185), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n22186));
    SB_CARRY add_3384_11 (.CI(n22818), .I0(n6715[8]), .I1(n755), .CO(n22819));
    SB_LUT4 add_3384_10_lut (.I0(GND_net), .I1(n6715[7]), .I2(n682), .I3(n22817), 
            .O(n6698[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_10 (.CI(n22817), .I0(n6715[7]), .I1(n682), .CO(n22818));
    SB_LUT4 add_3384_9_lut (.I0(GND_net), .I1(n6715[6]), .I2(n609), .I3(n22816), 
            .O(n6698[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_9 (.CI(n22816), .I0(n6715[6]), .I1(n609), .CO(n22817));
    SB_LUT4 add_3384_8_lut (.I0(GND_net), .I1(n6715[5]), .I2(n536), .I3(n22815), 
            .O(n6698[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_8 (.CI(n22815), .I0(n6715[5]), .I1(n536), .CO(n22816));
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_3979));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3384_7_lut (.I0(GND_net), .I1(n6715[4]), .I2(n463), .I3(n22814), 
            .O(n6698[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n22184), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n22184), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n22185));
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n22183), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_3978));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_3977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_3976));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_3975));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_3974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_3973));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_17 (.CI(n22183), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n22184));
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3972));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n22182), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n22182), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n22183));
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3384_7 (.CI(n22814), .I0(n6715[4]), .I1(n463), .CO(n22815));
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_3970));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n22181), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n22181), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n22182));
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n22180), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n22180), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n22181));
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_3969));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n22179), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n22179), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n22180));
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n22178), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_3968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_3967));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_3966));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_3965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_3964));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3384_6_lut (.I0(GND_net), .I1(n6715[3]), .I2(n390_adj_4133), 
            .I3(n22813), .O(n6698[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_3963));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3384_6 (.CI(n22813), .I0(n6715[3]), .I1(n390_adj_4133), 
            .CO(n22814));
    SB_LUT4 add_3384_5_lut (.I0(GND_net), .I1(n6715[2]), .I2(n317_adj_4132), 
            .I3(n22812), .O(n6698[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_3962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3384_5 (.CI(n22812), .I0(n6715[2]), .I1(n317_adj_4132), 
            .CO(n22813));
    SB_LUT4 add_3384_4_lut (.I0(GND_net), .I1(n6715[1]), .I2(n244_adj_4131), 
            .I3(n22811), .O(n6698[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_4 (.CI(n22811), .I0(n6715[1]), .I1(n244_adj_4131), 
            .CO(n22812));
    SB_LUT4 add_3384_3_lut (.I0(GND_net), .I1(n6715[0]), .I2(n171_adj_4130), 
            .I3(n22810), .O(n6698[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_3 (.CI(n22810), .I0(n6715[0]), .I1(n171_adj_4130), 
            .CO(n22811));
    SB_LUT4 add_3384_2_lut (.I0(GND_net), .I1(n29_adj_4129), .I2(n98_adj_4128), 
            .I3(GND_net), .O(n6698[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_2 (.CI(GND_net), .I0(n29_adj_4129), .I1(n98_adj_4128), 
            .CO(n22810));
    SB_LUT4 add_3383_17_lut (.I0(GND_net), .I1(n6698[14]), .I2(GND_net), 
            .I3(n22809), .O(n6680[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_3961));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_3959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_3958));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_16_lut (.I0(GND_net), .I1(n6698[13]), .I2(n1117_adj_4127), 
            .I3(n22808), .O(n6680[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_16 (.CI(n22808), .I0(n6698[13]), .I1(n1117_adj_4127), 
            .CO(n22809));
    SB_LUT4 add_3383_15_lut (.I0(GND_net), .I1(n6698[12]), .I2(n1044_adj_4125), 
            .I3(n22807), .O(n6680[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_15 (.CI(n22807), .I0(n6698[12]), .I1(n1044_adj_4125), 
            .CO(n22808));
    SB_LUT4 add_3383_14_lut (.I0(GND_net), .I1(n6698[11]), .I2(n971_adj_4124), 
            .I3(n22806), .O(n6680[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3957));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3383_14 (.CI(n22806), .I0(n6698[11]), .I1(n971_adj_4124), 
            .CO(n22807));
    SB_LUT4 add_3383_13_lut (.I0(GND_net), .I1(n6698[10]), .I2(n898_adj_4123), 
            .I3(n22805), .O(n6680[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_13 (.CI(n22805), .I0(n6698[10]), .I1(n898_adj_4123), 
            .CO(n22806));
    SB_LUT4 add_3383_12_lut (.I0(GND_net), .I1(n6698[9]), .I2(n825_adj_4122), 
            .I3(n22804), .O(n6680[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_12 (.CI(n22804), .I0(n6698[9]), .I1(n825_adj_4122), 
            .CO(n22805));
    SB_LUT4 add_3383_11_lut (.I0(GND_net), .I1(n6698[8]), .I2(n752_adj_4120), 
            .I3(n22803), .O(n6680[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_11 (.CI(n22803), .I0(n6698[8]), .I1(n752_adj_4120), 
            .CO(n22804));
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_10_lut (.I0(GND_net), .I1(n6698[7]), .I2(n679_adj_4119), 
            .I3(n22802), .O(n6680[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_10 (.CI(n22802), .I0(n6698[7]), .I1(n679_adj_4119), 
            .CO(n22803));
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3955));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_9_lut (.I0(GND_net), .I1(n6698[6]), .I2(n606), .I3(n22801), 
            .O(n6680[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_9 (.CI(n22801), .I0(n6698[6]), .I1(n606), .CO(n22802));
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_3954));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_8_lut (.I0(GND_net), .I1(n6698[5]), .I2(n533), .I3(n22800), 
            .O(n6680[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_8 (.CI(n22800), .I0(n6698[5]), .I1(n533), .CO(n22801));
    SB_LUT4 add_3383_7_lut (.I0(GND_net), .I1(n6698[4]), .I2(n460), .I3(n22799), 
            .O(n6680[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_7 (.CI(n22799), .I0(n6698[4]), .I1(n460), .CO(n22800));
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_3953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_6_lut (.I0(GND_net), .I1(n6698[3]), .I2(n387), .I3(n22798), 
            .O(n6680[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_6 (.CI(n22798), .I0(n6698[3]), .I1(n387), .CO(n22799));
    SB_LUT4 add_3383_5_lut (.I0(GND_net), .I1(n6698[2]), .I2(n314), .I3(n22797), 
            .O(n6680[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_5 (.CI(n22797), .I0(n6698[2]), .I1(n314), .CO(n22798));
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_3952));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_4_lut (.I0(GND_net), .I1(n6698[1]), .I2(n241), .I3(n22796), 
            .O(n6680[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_12 (.CI(n22178), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n22179));
    SB_CARRY add_3383_4 (.CI(n22796), .I0(n6698[1]), .I1(n241), .CO(n22797));
    SB_LUT4 i15197_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3383_3_lut (.I0(GND_net), .I1(n6698[0]), .I2(n168), .I3(n22795), 
            .O(n6680[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_3 (.CI(n22795), .I0(n6698[0]), .I1(n168), .CO(n22796));
    SB_LUT4 add_3383_2_lut (.I0(GND_net), .I1(n26_adj_4101), .I2(n95), 
            .I3(GND_net), .O(n6680[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3383_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3383_2 (.CI(GND_net), .I0(n26_adj_4101), .I1(n95), .CO(n22795));
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_3951));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3382_18_lut (.I0(GND_net), .I1(n6680[15]), .I2(GND_net), 
            .I3(n22794), .O(n6661[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_17_lut (.I0(GND_net), .I1(n6680[14]), .I2(GND_net), 
            .I3(n22793), .O(n6661[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_3950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_17 (.CI(n22793), .I0(n6680[14]), .I1(GND_net), .CO(n22794));
    SB_LUT4 add_3382_16_lut (.I0(GND_net), .I1(n6680[13]), .I2(n1114), 
            .I3(n22792), .O(n6661[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_16 (.CI(n22792), .I0(n6680[13]), .I1(n1114), .CO(n22793));
    SB_LUT4 add_3382_15_lut (.I0(GND_net), .I1(n6680[12]), .I2(n1041), 
            .I3(n22791), .O(n6661[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_3949));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_3948));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_3947));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_3946));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_3945));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3944));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3943));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3942));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3941));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_3939));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_3938));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_3937));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_3936));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_3935));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_3934));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_3933));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_3932));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3931));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3930));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3929));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_15 (.CI(n22791), .I0(n6680[12]), .I1(n1041), .CO(n22792));
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3928));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3382_14_lut (.I0(GND_net), .I1(n6680[11]), .I2(n968), 
            .I3(n22790), .O(n6661[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_14 (.CI(n22790), .I0(n6680[11]), .I1(n968), .CO(n22791));
    SB_LUT4 add_3382_13_lut (.I0(GND_net), .I1(n6680[10]), .I2(n895), 
            .I3(n22789), .O(n6661[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3927));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_13 (.CI(n22789), .I0(n6680[10]), .I1(n895), .CO(n22790));
    SB_LUT4 add_3382_12_lut (.I0(GND_net), .I1(n6680[9]), .I2(n822), .I3(n22788), 
            .O(n6661[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3926));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_12 (.CI(n22788), .I0(n6680[9]), .I1(n822), .CO(n22789));
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3924));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3382_11_lut (.I0(GND_net), .I1(n6680[8]), .I2(n749), .I3(n22787), 
            .O(n6661[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_11 (.CI(n22787), .I0(n6680[8]), .I1(n749), .CO(n22788));
    SB_LUT4 add_3382_10_lut (.I0(GND_net), .I1(n6680[7]), .I2(n676), .I3(n22786), 
            .O(n6661[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_10 (.CI(n22786), .I0(n6680[7]), .I1(n676), .CO(n22787));
    SB_LUT4 add_3382_9_lut (.I0(GND_net), .I1(n6680[6]), .I2(n603), .I3(n22785), 
            .O(n6661[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3923));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_9 (.CI(n22785), .I0(n6680[6]), .I1(n603), .CO(n22786));
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n22177), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_8_lut (.I0(GND_net), .I1(n6680[5]), .I2(n530), .I3(n22784), 
            .O(n6661[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_8 (.CI(n22784), .I0(n6680[5]), .I1(n530), .CO(n22785));
    SB_LUT4 add_3382_7_lut (.I0(GND_net), .I1(n6680[4]), .I2(n457), .I3(n22783), 
            .O(n6661[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_7 (.CI(n22783), .I0(n6680[4]), .I1(n457), .CO(n22784));
    SB_LUT4 add_3382_6_lut (.I0(GND_net), .I1(n6680[3]), .I2(n384), .I3(n22782), 
            .O(n6661[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_6 (.CI(n22782), .I0(n6680[3]), .I1(n384), .CO(n22783));
    SB_LUT4 add_3382_5_lut (.I0(GND_net), .I1(n6680[2]), .I2(n311), .I3(n22781), 
            .O(n6661[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_5 (.CI(n22781), .I0(n6680[2]), .I1(n311), .CO(n22782));
    SB_LUT4 add_3382_4_lut (.I0(GND_net), .I1(n6680[1]), .I2(n238), .I3(n22780), 
            .O(n6661[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_3922));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_3920));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_3919));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_4 (.CI(n22780), .I0(n6680[1]), .I1(n238), .CO(n22781));
    SB_LUT4 add_3382_3_lut (.I0(GND_net), .I1(n6680[0]), .I2(n165), .I3(n22779), 
            .O(n6661[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_3 (.CI(n22779), .I0(n6680[0]), .I1(n165), .CO(n22780));
    SB_LUT4 add_3382_2_lut (.I0(GND_net), .I1(n23_adj_4045), .I2(n92), 
            .I3(GND_net), .O(n6661[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_2 (.CI(GND_net), .I0(n23_adj_4045), .I1(n92), .CO(n22779));
    SB_LUT4 add_3381_19_lut (.I0(GND_net), .I1(n6661[16]), .I2(GND_net), 
            .I3(n22778), .O(n6641[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3381_18_lut (.I0(GND_net), .I1(n6661[15]), .I2(GND_net), 
            .I3(n22777), .O(n6641[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3917));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15198_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15199_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15199_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3381_18 (.CI(n22777), .I0(n6661[15]), .I1(GND_net), .CO(n22778));
    SB_LUT4 add_3381_17_lut (.I0(GND_net), .I1(n6661[14]), .I2(GND_net), 
            .I3(n22776), .O(n6641[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_17 (.CI(n22776), .I0(n6661[14]), .I1(GND_net), .CO(n22777));
    SB_LUT4 add_3381_16_lut (.I0(GND_net), .I1(n6661[13]), .I2(n1111), 
            .I3(n22775), .O(n6641[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_16 (.CI(n22775), .I0(n6661[13]), .I1(n1111), .CO(n22776));
    SB_LUT4 add_3381_15_lut (.I0(GND_net), .I1(n6661[12]), .I2(n1038), 
            .I3(n22774), .O(n6641[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_15 (.CI(n22774), .I0(n6661[12]), .I1(n1038), .CO(n22775));
    SB_LUT4 add_3381_14_lut (.I0(GND_net), .I1(n6661[11]), .I2(n965), 
            .I3(n22773), .O(n6641[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_14 (.CI(n22773), .I0(n6661[11]), .I1(n965), .CO(n22774));
    SB_LUT4 add_3381_13_lut (.I0(GND_net), .I1(n6661[10]), .I2(n892), 
            .I3(n22772), .O(n6641[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_13 (.CI(n22772), .I0(n6661[10]), .I1(n892), .CO(n22773));
    SB_LUT4 add_3381_12_lut (.I0(GND_net), .I1(n6661[9]), .I2(n819), .I3(n22771), 
            .O(n6641[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_12 (.CI(n22771), .I0(n6661[9]), .I1(n819), .CO(n22772));
    SB_LUT4 add_3381_11_lut (.I0(GND_net), .I1(n6661[8]), .I2(n746), .I3(n22770), 
            .O(n6641[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_11 (.CI(n22770), .I0(n6661[8]), .I1(n746), .CO(n22771));
    SB_CARRY sub_3_add_2_11 (.CI(n22177), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n22178));
    SB_LUT4 i15200_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3492[23]), .I1(n257[23]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n22176), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3467[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_10 (.CI(n22176), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n22177));
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3492[22]), .I1(n257[22]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3381_10_lut (.I0(GND_net), .I1(n6661[7]), .I2(n673), .I3(n22769), 
            .O(n6641[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n22175), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_10 (.CI(n22769), .I0(n6661[7]), .I1(n673), .CO(n22770));
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3467[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3916));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3492[21]), .I1(n257[21]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3381_9_lut (.I0(GND_net), .I1(n6661[6]), .I2(n600), .I3(n22768), 
            .O(n6641[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_9 (.CI(n22768), .I0(n6661[6]), .I1(n600), .CO(n22769));
    SB_LUT4 add_3381_8_lut (.I0(GND_net), .I1(n6661[5]), .I2(n527), .I3(n22767), 
            .O(n6641[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_8 (.CI(n22767), .I0(n6661[5]), .I1(n527), .CO(n22768));
    SB_LUT4 add_3381_7_lut (.I0(GND_net), .I1(n6661[4]), .I2(n454), .I3(n22766), 
            .O(n6641[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_7 (.CI(n22766), .I0(n6661[4]), .I1(n454), .CO(n22767));
    SB_LUT4 add_3381_6_lut (.I0(GND_net), .I1(n6661[3]), .I2(n381), .I3(n22765), 
            .O(n6641[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3467[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_9 (.CI(n22175), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n22176));
    SB_CARRY add_3381_6 (.CI(n22765), .I0(n6661[3]), .I1(n381), .CO(n22766));
    SB_LUT4 add_3381_5_lut (.I0(GND_net), .I1(n6661[2]), .I2(n308), .I3(n22764), 
            .O(n6641[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3492[20]), .I1(n257[20]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3915));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3467[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3492[19]), .I1(n257[19]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3467[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3492[18]), .I1(n257[18]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3467[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3492[17]), .I1(n257[17]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3467[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3492[16]), .I1(n257[16]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3467[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3492[15]), .I1(n257[15]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3467[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3492[14]), .I1(n257[14]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3467[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3492[13]), .I1(n257[13]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3467[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3492[12]), .I1(n257[12]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3467[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3492[11]), .I1(n257[11]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3467[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3492[10]), .I1(n257[10]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3467[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3492[9]), .I1(n257[9]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3467[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3381_5 (.CI(n22764), .I0(n6661[2]), .I1(n308), .CO(n22765));
    SB_LUT4 add_3381_4_lut (.I0(GND_net), .I1(n6661[1]), .I2(n235), .I3(n22763), 
            .O(n6641[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3492[8]), .I1(n257[8]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3467[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3492[7]), .I1(n257[7]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3467[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3492[6]), .I1(n257[6]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3467[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3492[5]), .I1(n257[5]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3467[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3492[4]), .I1(n257[4]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3467[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3381_4 (.CI(n22763), .I0(n6661[1]), .I1(n235), .CO(n22764));
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3492[3]), .I1(n257[3]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3381_3_lut (.I0(GND_net), .I1(n6661[0]), .I2(n162), .I3(n22762), 
            .O(n6641[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3467[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15190_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15190_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15201_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15202_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15203_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15204_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4275));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3381_3 (.CI(n22762), .I0(n6661[0]), .I1(n162), .CO(n22763));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n22174), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3914));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3381_2_lut (.I0(GND_net), .I1(n20_adj_4276), .I2(n89_adj_4277), 
            .I3(GND_net), .O(n6641[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3381_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3381_2 (.CI(GND_net), .I0(n20_adj_4276), .I1(n89_adj_4277), 
            .CO(n22762));
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3492[2]), .I1(n257[2]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3467[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3380_20_lut (.I0(GND_net), .I1(n6641[17]), .I2(GND_net), 
            .I3(n22761), .O(n6620[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3380_19_lut (.I0(GND_net), .I1(n6641[16]), .I2(GND_net), 
            .I3(n22760), .O(n6620[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_19 (.CI(n22760), .I0(n6641[16]), .I1(GND_net), .CO(n22761));
    SB_LUT4 add_3380_18_lut (.I0(GND_net), .I1(n6641[15]), .I2(GND_net), 
            .I3(n22759), .O(n6620[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_18 (.CI(n22759), .I0(n6641[15]), .I1(GND_net), .CO(n22760));
    SB_LUT4 add_3380_17_lut (.I0(GND_net), .I1(n6641[14]), .I2(GND_net), 
            .I3(n22758), .O(n6620[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_17 (.CI(n22758), .I0(n6641[14]), .I1(GND_net), .CO(n22759));
    SB_LUT4 add_3380_16_lut (.I0(GND_net), .I1(n6641[13]), .I2(n1108_adj_4278), 
            .I3(n22757), .O(n6620[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_8 (.CI(n22174), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n22175));
    SB_CARRY add_3380_16 (.CI(n22757), .I0(n6641[13]), .I1(n1108_adj_4278), 
            .CO(n22758));
    SB_LUT4 add_3380_15_lut (.I0(GND_net), .I1(n6641[12]), .I2(n1035_adj_4279), 
            .I3(n22756), .O(n6620[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_15 (.CI(n22756), .I0(n6641[12]), .I1(n1035_adj_4279), 
            .CO(n22757));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n22173), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3380_14_lut (.I0(GND_net), .I1(n6641[11]), .I2(n962_adj_4280), 
            .I3(n22755), .O(n6620[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3368[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_3380_14 (.CI(n22755), .I0(n6641[11]), .I1(n962_adj_4280), 
            .CO(n22756));
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4281));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4146));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4282));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3380_13_lut (.I0(GND_net), .I1(n6641[10]), .I2(n889_adj_4282), 
            .I3(n22754), .O(n6620[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3492[1]), .I1(n257[1]), .I2(n256_adj_4252), 
            .I3(GND_net), .O(duty_23__N_3467[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3467[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3491), .I3(GND_net), .O(duty_23__N_3368[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4145));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4162));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_3_add_2_7 (.CI(n22173), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n22174));
    SB_CARRY add_3380_13 (.CI(n22754), .I0(n6641[10]), .I1(n889_adj_4282), 
            .CO(n22755));
    SB_LUT4 add_3380_12_lut (.I0(GND_net), .I1(n6641[9]), .I2(n816_adj_4281), 
            .I3(n22753), .O(n6620[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_12 (.CI(n22753), .I0(n6641[9]), .I1(n816_adj_4281), 
            .CO(n22754));
    SB_LUT4 add_3380_9_lut (.I0(GND_net), .I1(n6641[6]), .I2(n597), .I3(n22750), 
            .O(n6620[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n22172), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n22172), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n22173));
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n22171), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_3913));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3368[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_3_add_2_5 (.CI(n22171), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n22172));
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n22170), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3380_11_lut (.I0(GND_net), .I1(n6641[8]), .I2(n743_adj_4275), 
            .I3(n22752), .O(n6620[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n2552[23]), .I3(n21967), .O(\PID_CONTROLLER.integral_23__N_3392 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n2552[22]), .I3(n21966), .O(\PID_CONTROLLER.integral_23__N_3392 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_24 (.CI(n21966), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n2552[22]), .CO(n21967));
    SB_CARRY sub_3_add_2_4 (.CI(n22170), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n22171));
    SB_LUT4 add_560_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n2552[21]), .I3(n21965), .O(\PID_CONTROLLER.integral_23__N_3392 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_23 (.CI(n21965), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n2552[21]), .CO(n21966));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n22169), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n2552[20]), .I3(n21964), .O(\PID_CONTROLLER.integral_23__N_3392 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n22169), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n22170));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_22 (.CI(n21964), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n2552[20]), .CO(n21965));
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n22169));
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_3912));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_560_11 (.CI(n21953), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n2552[9]), .CO(n21954));
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3368[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3368[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3368[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3368[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3368[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3368[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3368[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3368[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3368[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3368[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3368[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3368[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3368[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3368[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3368[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3368[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3368[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3368[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3368[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3368[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3368[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3392 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15191_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15191_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_560_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n2552[19]), .I3(n21963), .O(\PID_CONTROLLER.integral_23__N_3392 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_3911));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4280));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_3910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15192_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15192_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4304[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_560_21 (.CI(n21963), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n2552[19]), .CO(n21964));
    SB_LUT4 add_560_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n2552[18]), .I3(n21962), .O(\PID_CONTROLLER.integral_23__N_3392 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4279));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4278));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_560_20 (.CI(n21962), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n2552[18]), .CO(n21963));
    SB_LUT4 add_560_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n2552[17]), .I3(n21961), .O(\PID_CONTROLLER.integral_23__N_3392 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24335_3_lut_4_lut (.I0(duty_23__N_3492[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3492[2]), .O(n29398));   // verilog/motorControl.v(38[19:35])
    defparam i24335_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3492[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4240));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_3909));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_3908));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_560_19 (.CI(n21961), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n2552[17]), .CO(n21962));
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n4998[0]), .I2(n5002[0]), 
            .I3(n22028), .O(duty_23__N_3492[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n22027), .O(duty_23__N_3492[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n22027), .I0(n106[22]), .I1(n155[22]), .CO(n22028));
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n22026), .O(duty_23__N_3492[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n2552[16]), .I3(n21960), .O(\PID_CONTROLLER.integral_23__N_3392 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3906));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3905));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18015_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [18]), 
            .I2(n4_adj_4301), .I3(n7127[1]), .O(n6_adj_4139));   // verilog/motorControl.v(34[25:36])
    defparam i18015_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1451 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [18]), 
            .I2(n7127[1]), .I3(n4_adj_4301), .O(n7120[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1451.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3903));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_23 (.CI(n22026), .I0(n106[21]), .I1(n155[21]), .CO(n22027));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n22025), .O(duty_23__N_3492[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_18 (.CI(n21960), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n2552[16]), .CO(n21961));
    SB_LUT4 add_560_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n2552[15]), .I3(n21959), .O(\PID_CONTROLLER.integral_23__N_3392 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24372_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3492[3]), 
            .I2(duty_23__N_3492[2]), .I3(PWMLimit[2]), .O(n29435));   // verilog/motorControl.v(36[10:25])
    defparam i24372_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_3901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_831_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3492[3]), 
            .I2(duty_23__N_3492[2]), .I3(GND_net), .O(n6_adj_4185));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i2_3_lut_4_lut_adj_1452 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [18]), 
            .I2(n7127[0]), .I3(n21784), .O(n7120[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1452.LUT_INIT = 16'h8778;
    SB_LUT4 i18007_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [18]), 
            .I2(n21784), .I3(n7127[0]), .O(n4_adj_4301));   // verilog/motorControl.v(34[25:36])
    defparam i18007_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i17996_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3392 [18]), .I3(\Ki[1] ), 
            .O(n21784));   // verilog/motorControl.v(34[25:36])
    defparam i17996_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i17994_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3392 [18]), .I3(\Ki[1] ), 
            .O(n7120[0]));   // verilog/motorControl.v(34[25:36])
    defparam i17994_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4266));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15193_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15193_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_22 (.CI(n22025), .I0(n106[20]), .I1(n155[20]), .CO(n22026));
    SB_CARRY add_560_17 (.CI(n21959), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n2552[15]), .CO(n21960));
    SB_LUT4 add_560_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n2552[14]), .I3(n21958), .O(\PID_CONTROLLER.integral_23__N_3392 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n22024), .O(duty_23__N_3492[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24303_2_lut_4_lut (.I0(duty_23__N_3492[21]), .I1(n257[21]), 
            .I2(duty_23__N_3492[9]), .I3(n257[9]), .O(n29366));
    defparam i24303_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i24313_2_lut_4_lut (.I0(duty_23__N_3492[16]), .I1(n257[16]), 
            .I2(duty_23__N_3492[7]), .I3(n257[7]), .O(n29376));
    defparam i24313_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4277));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4276));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_21 (.CI(n22024), .I0(n106[19]), .I1(n155[19]), .CO(n22025));
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n22023), .O(duty_23__N_3492[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_20 (.CI(n22023), .I0(n106[18]), .I1(n155[18]), .CO(n22024));
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n22022), .O(duty_23__N_3492[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_16 (.CI(n21958), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n2552[14]), .CO(n21959));
    SB_LUT4 i18077_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [20]), 
            .I2(n21861), .I3(n7138[0]), .O(n4_adj_4255));   // verilog/motorControl.v(34[25:36])
    defparam i18077_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_560_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n2552[13]), .I3(n21957), .O(\PID_CONTROLLER.integral_23__N_3392 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1453 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [20]), 
            .I2(n7138[0]), .I3(n21861), .O(n7133[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1453.LUT_INIT = 16'h8778;
    SB_CARRY add_12_19 (.CI(n22022), .I0(n106[17]), .I1(n155[17]), .CO(n22023));
    SB_LUT4 i2_3_lut_4_lut_adj_1454 (.I0(n62), .I1(n131), .I2(n7133[0]), 
            .I3(n204), .O(n7127[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1454.LUT_INIT = 16'h8778;
    SB_LUT4 i18046_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n7133[0]), 
            .O(n4_adj_4190));   // verilog/motorControl.v(34[25:36])
    defparam i18046_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i18066_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3392 [20]), .I3(\Ki[1] ), 
            .O(n21861));   // verilog/motorControl.v(34[25:36])
    defparam i18066_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i18064_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3392 [20]), .I3(\Ki[1] ), 
            .O(n7133[0]));   // verilog/motorControl.v(34[25:36])
    defparam i18064_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i15194_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15194_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24337_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3492[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3492[9]), .O(n29400));
    defparam i24337_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n22021), .O(duty_23__N_3492[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_15 (.CI(n21957), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n2552[13]), .CO(n21958));
    SB_LUT4 add_560_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n2552[12]), .I3(n21956), .O(\PID_CONTROLLER.integral_23__N_3392 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24348_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3492[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3492[7]), .O(n29411));
    defparam i24348_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_12_18 (.CI(n22021), .I0(n106[16]), .I1(n155[16]), .CO(n22022));
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n22020), .O(duty_23__N_3492[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_17 (.CI(n22020), .I0(n106[15]), .I1(n155[15]), .CO(n22021));
    SB_CARRY add_3380_11 (.CI(n22752), .I0(n6641[8]), .I1(n743_adj_4275), 
            .CO(n22753));
    SB_LUT4 add_3380_10_lut (.I0(GND_net), .I1(n6641[7]), .I2(n670_adj_4302), 
            .I3(n22751), .O(n6620[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3380_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3380_10 (.CI(n22751), .I0(n6641[7]), .I1(n670_adj_4302), 
            .CO(n22752));
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n22019), .O(duty_23__N_3492[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n22019), .I0(n106[14]), .I1(n155[14]), .CO(n22020));
    SB_LUT4 i15195_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3440 ), 
            .I2(GND_net), .I3(GND_net), .O(n2552[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i15195_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18033_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3392 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3392 [19]), 
            .O(n7127[0]));   // verilog/motorControl.v(34[25:36])
    defparam i18033_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n22018), .O(duty_23__N_3492[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n22018), .I0(n106[13]), .I1(n155[13]), .CO(n22019));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n22017), .O(duty_23__N_3492[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_14 (.CI(n21956), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n2552[12]), .CO(n21957));
    SB_CARRY add_12_14 (.CI(n22017), .I0(n106[12]), .I1(n155[12]), .CO(n22018));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n22016), .O(duty_23__N_3492[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[23]), 
            .I3(n22237), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n2552[11]), .I3(n21955), .O(\PID_CONTROLLER.integral_23__N_3392 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[22]), 
            .I3(n22236), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n22236), .I0(GND_net), .I1(n1_adj_4304[22]), 
            .CO(n22237));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[21]), 
            .I3(n22235), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n22235), .I0(GND_net), .I1(n1_adj_4304[21]), 
            .CO(n22236));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[20]), 
            .I3(n22234), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n22234), .I0(GND_net), .I1(n1_adj_4304[20]), 
            .CO(n22235));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[19]), 
            .I3(n22233), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n22233), .I0(GND_net), .I1(n1_adj_4304[19]), 
            .CO(n22234));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[18]), 
            .I3(n22232), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n22232), .I0(GND_net), .I1(n1_adj_4304[18]), 
            .CO(n22233));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[17]), 
            .I3(n22231), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n22231), .I0(GND_net), .I1(n1_adj_4304[17]), 
            .CO(n22232));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[16]), 
            .I3(n22230), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n22230), .I0(GND_net), .I1(n1_adj_4304[16]), 
            .CO(n22231));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[15]), 
            .I3(n22229), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n22229), .I0(GND_net), .I1(n1_adj_4304[15]), 
            .CO(n22230));
    SB_CARRY add_560_13 (.CI(n21955), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n2552[11]), .CO(n21956));
    SB_LUT4 add_560_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n2552[10]), .I3(n21954), .O(\PID_CONTROLLER.integral_23__N_3392 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[14]), 
            .I3(n22228), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n22228), .I0(GND_net), .I1(n1_adj_4304[14]), 
            .CO(n22229));
    SB_CARRY add_12_13 (.CI(n22016), .I0(n106[11]), .I1(n155[11]), .CO(n22017));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[13]), 
            .I3(n22227), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_12 (.CI(n21954), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n2552[10]), .CO(n21955));
    SB_LUT4 add_560_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n2552[9]), .I3(n21953), .O(\PID_CONTROLLER.integral_23__N_3392 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_9 (.CI(n21951), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n2552[7]), .CO(n21952));
    SB_CARRY unary_minus_16_add_3_15 (.CI(n22227), .I0(GND_net), .I1(n1_adj_4304[13]), 
            .CO(n22228));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[12]), 
            .I3(n22226), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n22226), .I0(GND_net), .I1(n1_adj_4304[12]), 
            .CO(n22227));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[11]), 
            .I3(n22225), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n22225), .I0(GND_net), .I1(n1_adj_4304[11]), 
            .CO(n22226));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[10]), 
            .I3(n22224), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n22224), .I0(GND_net), .I1(n1_adj_4304[10]), 
            .CO(n22225));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[9]), 
            .I3(n22223), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n22223), .I0(GND_net), .I1(n1_adj_4304[9]), 
            .CO(n22224));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[8]), 
            .I3(n22222), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n22222), .I0(GND_net), .I1(n1_adj_4304[8]), 
            .CO(n22223));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[7]), 
            .I3(n22221), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n22015), .O(duty_23__N_3492[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n22221), .I0(GND_net), .I1(n1_adj_4304[7]), 
            .CO(n22222));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[6]), 
            .I3(n22220), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n22220), .I0(GND_net), .I1(n1_adj_4304[6]), 
            .CO(n22221));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4304[5]), 
            .I3(n22219), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n22015), .I0(n106[10]), .I1(n155[10]), .CO(n22016));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n22014), 
            .O(duty_23__N_3492[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n22014), .I0(n106[9]), .I1(n155[9]), .CO(n22015));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n22013), 
            .O(duty_23__N_3492[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n29954, VCC_net, INHA_c, clk32MHz, n13407, GND_net, 
            n13405, \pwm_counter[6] , \pwm_counter[8] , \pwm_counter[7] , 
            \pwm_counter[13] , \pwm_counter[10] , \pwm_counter[9] , \pwm_counter[17] , 
            \pwm_counter[22] , \pwm_counter[14] , \pwm_counter[18] , \pwm_counter[21] , 
            \pwm_counter[16] , \pwm_counter[12] , \pwm_counter[15] , \pwm_counter[19] , 
            \pwm_counter[11] , \pwm_counter[20] , \pwm_counter[31] , \pwm_counter[0] , 
            \pwm_counter[5] , \pwm_counter[4] , \pwm_counter[3] , \pwm_counter[2] , 
            \pwm_counter[1] ) /* synthesis syn_module_defined=1 */ ;
    input n29954;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n13407;
    input GND_net;
    output n13405;
    output \pwm_counter[6] ;
    output \pwm_counter[8] ;
    output \pwm_counter[7] ;
    output \pwm_counter[13] ;
    output \pwm_counter[10] ;
    output \pwm_counter[9] ;
    output \pwm_counter[17] ;
    output \pwm_counter[22] ;
    output \pwm_counter[14] ;
    output \pwm_counter[18] ;
    output \pwm_counter[21] ;
    output \pwm_counter[16] ;
    output \pwm_counter[12] ;
    output \pwm_counter[15] ;
    output \pwm_counter[19] ;
    output \pwm_counter[11] ;
    output \pwm_counter[20] ;
    output \pwm_counter[31] ;
    output \pwm_counter[0] ;
    output \pwm_counter[5] ;
    output \pwm_counter[4] ;
    output \pwm_counter[3] ;
    output \pwm_counter[2] ;
    output \pwm_counter[1] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n10, n14, n27151, n18, n24, n22, n26, n21, pwm_counter_31__N_531;
    wire [31:0]n133;
    
    wire n22404, n22403, n22402, n22401, n22400, n22399, n22398, 
        n22397, n22396, n22395, n22394, n22393, n22392, n22391, 
        n22390, n22389, n22388, n22387, n22386, n22385, n22384, 
        n22383, n22382, n22381, n22380, n22379, n22378, n22377, 
        n22376, n22375, n22374;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n29954), 
            .R(n13407));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[29]), .I2(pwm_counter[25]), 
            .I3(pwm_counter[26]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(pwm_counter[30]), .I1(n14), .I2(n10), .I3(pwm_counter[24]), 
            .O(n13405));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(\pwm_counter[6] ), .I1(\pwm_counter[8] ), .I2(\pwm_counter[7] ), 
            .I3(GND_net), .O(n27151));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n27151), .I1(\pwm_counter[13] ), .I2(\pwm_counter[10] ), 
            .I3(\pwm_counter[9] ), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(\pwm_counter[17] ), .I1(\pwm_counter[22] ), .I2(\pwm_counter[14] ), 
            .I3(\pwm_counter[18] ), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(\pwm_counter[21] ), .I1(n13405), .I2(\pwm_counter[16] ), 
            .I3(\pwm_counter[12] ), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(\pwm_counter[15] ), .I1(n24), .I2(n18), .I3(\pwm_counter[19] ), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(\pwm_counter[11] ), .I1(\pwm_counter[20] ), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14975_4_lut (.I0(n21), .I1(\pwm_counter[31] ), .I2(n26), 
            .I3(n22), .O(pwm_counter_31__N_531));   // verilog/pwm.v(18[8:40])
    defparam i14975_4_lut.LUT_INIT = 16'h3332;
    SB_DFFSR pwm_counter_1123__i0 (.Q(\pwm_counter[0] ), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1123_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[31] ), 
            .I3(n22404), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1123_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n22403), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_32 (.CI(n22403), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n22404));
    SB_LUT4 pwm_counter_1123_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n22402), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_31 (.CI(n22402), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n22403));
    SB_LUT4 pwm_counter_1123_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n22401), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_30 (.CI(n22401), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n22402));
    SB_LUT4 pwm_counter_1123_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n22400), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_29 (.CI(n22400), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n22401));
    SB_LUT4 pwm_counter_1123_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n22399), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_28 (.CI(n22399), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n22400));
    SB_LUT4 pwm_counter_1123_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n22398), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_27 (.CI(n22398), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n22399));
    SB_LUT4 pwm_counter_1123_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n22397), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_26 (.CI(n22397), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n22398));
    SB_LUT4 pwm_counter_1123_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n22396), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_25 (.CI(n22396), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n22397));
    SB_LUT4 pwm_counter_1123_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[22] ), 
            .I3(n22395), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_24 (.CI(n22395), .I0(GND_net), .I1(\pwm_counter[22] ), 
            .CO(n22396));
    SB_LUT4 pwm_counter_1123_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[21] ), 
            .I3(n22394), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_23 (.CI(n22394), .I0(GND_net), .I1(\pwm_counter[21] ), 
            .CO(n22395));
    SB_LUT4 pwm_counter_1123_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[20] ), 
            .I3(n22393), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_22 (.CI(n22393), .I0(GND_net), .I1(\pwm_counter[20] ), 
            .CO(n22394));
    SB_LUT4 pwm_counter_1123_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[19] ), 
            .I3(n22392), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_21 (.CI(n22392), .I0(GND_net), .I1(\pwm_counter[19] ), 
            .CO(n22393));
    SB_LUT4 pwm_counter_1123_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[18] ), 
            .I3(n22391), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_20 (.CI(n22391), .I0(GND_net), .I1(\pwm_counter[18] ), 
            .CO(n22392));
    SB_LUT4 pwm_counter_1123_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[17] ), 
            .I3(n22390), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_19 (.CI(n22390), .I0(GND_net), .I1(\pwm_counter[17] ), 
            .CO(n22391));
    SB_LUT4 pwm_counter_1123_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[16] ), 
            .I3(n22389), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_18 (.CI(n22389), .I0(GND_net), .I1(\pwm_counter[16] ), 
            .CO(n22390));
    SB_LUT4 pwm_counter_1123_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[15] ), 
            .I3(n22388), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_17 (.CI(n22388), .I0(GND_net), .I1(\pwm_counter[15] ), 
            .CO(n22389));
    SB_LUT4 pwm_counter_1123_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[14] ), 
            .I3(n22387), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_16 (.CI(n22387), .I0(GND_net), .I1(\pwm_counter[14] ), 
            .CO(n22388));
    SB_LUT4 pwm_counter_1123_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[13] ), 
            .I3(n22386), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_15 (.CI(n22386), .I0(GND_net), .I1(\pwm_counter[13] ), 
            .CO(n22387));
    SB_LUT4 pwm_counter_1123_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[12] ), 
            .I3(n22385), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_14 (.CI(n22385), .I0(GND_net), .I1(\pwm_counter[12] ), 
            .CO(n22386));
    SB_LUT4 pwm_counter_1123_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[11] ), 
            .I3(n22384), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_13 (.CI(n22384), .I0(GND_net), .I1(\pwm_counter[11] ), 
            .CO(n22385));
    SB_LUT4 pwm_counter_1123_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[10] ), 
            .I3(n22383), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_12 (.CI(n22383), .I0(GND_net), .I1(\pwm_counter[10] ), 
            .CO(n22384));
    SB_LUT4 pwm_counter_1123_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[9] ), 
            .I3(n22382), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_11 (.CI(n22382), .I0(GND_net), .I1(\pwm_counter[9] ), 
            .CO(n22383));
    SB_LUT4 pwm_counter_1123_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[8] ), 
            .I3(n22381), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_10 (.CI(n22381), .I0(GND_net), .I1(\pwm_counter[8] ), 
            .CO(n22382));
    SB_LUT4 pwm_counter_1123_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[7] ), 
            .I3(n22380), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_9 (.CI(n22380), .I0(GND_net), .I1(\pwm_counter[7] ), 
            .CO(n22381));
    SB_LUT4 pwm_counter_1123_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[6] ), 
            .I3(n22379), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_8 (.CI(n22379), .I0(GND_net), .I1(\pwm_counter[6] ), 
            .CO(n22380));
    SB_LUT4 pwm_counter_1123_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[5] ), 
            .I3(n22378), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_7 (.CI(n22378), .I0(GND_net), .I1(\pwm_counter[5] ), 
            .CO(n22379));
    SB_LUT4 pwm_counter_1123_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[4] ), 
            .I3(n22377), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_6 (.CI(n22377), .I0(GND_net), .I1(\pwm_counter[4] ), 
            .CO(n22378));
    SB_LUT4 pwm_counter_1123_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[3] ), 
            .I3(n22376), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_5 (.CI(n22376), .I0(GND_net), .I1(\pwm_counter[3] ), 
            .CO(n22377));
    SB_LUT4 pwm_counter_1123_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[2] ), 
            .I3(n22375), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_4 (.CI(n22375), .I0(GND_net), .I1(\pwm_counter[2] ), 
            .CO(n22376));
    SB_LUT4 pwm_counter_1123_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[1] ), 
            .I3(n22374), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_3 (.CI(n22374), .I0(GND_net), .I1(\pwm_counter[1] ), 
            .CO(n22375));
    SB_LUT4 pwm_counter_1123_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1123_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1123_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\pwm_counter[0] ), 
            .CO(n22374));
    SB_DFFSR pwm_counter_1123__i1 (.Q(\pwm_counter[1] ), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i2 (.Q(\pwm_counter[2] ), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i3 (.Q(\pwm_counter[3] ), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i4 (.Q(\pwm_counter[4] ), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i5 (.Q(\pwm_counter[5] ), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i6 (.Q(\pwm_counter[6] ), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i7 (.Q(\pwm_counter[7] ), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i8 (.Q(\pwm_counter[8] ), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i9 (.Q(\pwm_counter[9] ), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i10 (.Q(\pwm_counter[10] ), .C(clk32MHz), 
            .D(n133[10]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i11 (.Q(\pwm_counter[11] ), .C(clk32MHz), 
            .D(n133[11]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i12 (.Q(\pwm_counter[12] ), .C(clk32MHz), 
            .D(n133[12]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i13 (.Q(\pwm_counter[13] ), .C(clk32MHz), 
            .D(n133[13]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i14 (.Q(\pwm_counter[14] ), .C(clk32MHz), 
            .D(n133[14]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i15 (.Q(\pwm_counter[15] ), .C(clk32MHz), 
            .D(n133[15]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i16 (.Q(\pwm_counter[16] ), .C(clk32MHz), 
            .D(n133[16]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i17 (.Q(\pwm_counter[17] ), .C(clk32MHz), 
            .D(n133[17]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i18 (.Q(\pwm_counter[18] ), .C(clk32MHz), 
            .D(n133[18]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i19 (.Q(\pwm_counter[19] ), .C(clk32MHz), 
            .D(n133[19]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i20 (.Q(\pwm_counter[20] ), .C(clk32MHz), 
            .D(n133[20]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i21 (.Q(\pwm_counter[21] ), .C(clk32MHz), 
            .D(n133[21]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i22 (.Q(\pwm_counter[22] ), .C(clk32MHz), 
            .D(n133[22]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1123__i31 (.Q(\pwm_counter[31] ), .C(clk32MHz), 
            .D(n133[31]), .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    
endmodule
//
// Verilog Description of module coms
//

module coms (GND_net, \data_out_frame[25] , rx_data, setpoint, clk32MHz, 
            n14885, IntegralLimit, n14884, n14883, n10896, \data_in_frame[1] , 
            \data_in_frame[2] , n4141, \data_in_frame[3] , \data_out_frame[23] , 
            \data_out_frame[20] , \data_out_frame[16] , \data_out_frame[17] , 
            \data_out_frame[18] , \data_out_frame[19] , \data_out_frame[5] , 
            \data_out_frame[6] , \data_out_frame[7] , n14882, \data_in_frame[6] , 
            \data_in_frame[8] , n14881, n14880, n14879, \data_in_frame[5] , 
            n14878, \data_in_frame[4] , n14877, n14876, rx_data_ready, 
            n14875, n14874, \data_out_frame[15] , n14873, \data_out_frame[12] , 
            \data_out_frame[10] , \data_out_frame[9] , \data_out_frame[13] , 
            \data_out_frame[24] , n2252, \data_in[1] , \data_in[0] , 
            \data_in[2] , \data_in[3] , n63, n3, \data_in_frame[9] , 
            \data_in_frame[11] , \data_in_frame[10] , \data_in_frame[13] , 
            \FRAME_MATCHER.state_31__N_2380[2] , \data_in_frame[12] , n4137, 
            \data_out_frame[14] , \data_out_frame[11] , \data_out_frame[8] , 
            \data_out_frame[27][0] , n4, tx_active, n14641, n24343, 
            n1, DE_c, n26748, n7, n7_adj_3, LED_c, n5, n26399, 
            n14833, PWMLimit, n14832, control_mode, n28285, n30820, 
            n15337, n15336, n15335, n15334, n15333, n15332, n15331, 
            n15330, n15329, n15328, n15327, n15326, n15325, n15324, 
            n15323, n15322, n15321, n15320, n15319, n15318, n15317, 
            n15316, n15315, n15314, n15313, n15312, n15311, n15310, 
            n15309, n15308, n15132, neopxl_color, n15131, n15130, 
            n15129, n15128, n15127, n15126, n15125, n15124, n15123, 
            n15122, n15121, n15120, n15119, n15118, n15117, n15116, 
            n15115, n15114, n15113, n15112, n15111, n15110, n15109, 
            n15108, n15107, n15106, n15105, n15104, n15103, n15102, 
            n15101, n15100, n15099, n15098, n15097, n15096, n15095, 
            n15094, n15093, n15092, n15091, n15090, n15089, n15088, 
            n15087, n15086, n15085, n15084, n15083, n15082, n15081, 
            n15080, n15079, n15077, n15076, n15075, n15074, n15073, 
            n15072, n15071, n15070, n15069, n15068, n15067, n15066, 
            n15065, n15064, n15063, n15062, n15061, n15060, n15059, 
            n15058, n15057, n15056, n15055, n15054, n15053, n15052, 
            n15051, n15050, n15049, n15048, n15047, n15046, n15045, 
            n15044, n15043, n15042, n15041, n15040, n15039, n15038, 
            n15037, n15036, n15035, n15034, n15033, n15032, n15031, 
            n15030, n15029, n15028, n15027, n15026, n15025, n15024, 
            n15023, n15022, n15021, n15020, n27156, n15019, n15018, 
            n15017, n15016, n15015, n15014, n15013, n15012, n15011, 
            n15010, n15009, n15008, n15007, n15006, n15005, n15004, 
            n15003, n15002, n15001, n15000, n14999, n14998, n14997, 
            n14996, n14995, n14994, n14993, n14992, n14991, n14990, 
            n14989, n14830, n14829, \Ki[0] , n14828, \Kp[0] , n14827, 
            n14988, n14987, n14986, n14985, n14984, n14983, n14982, 
            n14818, n14981, n14980, n14979, n14978, n14977, n14976, 
            n14975, n14974, n14973, n14972, n14971, n14970, n14969, 
            n14968, n14967, n14966, n14965, n14964, n14963, n14962, 
            n14961, n14960, n14959, n14958, n14957, n14956, \Ki[15] , 
            n14955, \Ki[14] , n14954, \Ki[13] , n14953, \Ki[12] , 
            n14952, \Ki[11] , n14951, \Ki[10] , n14950, \Ki[9] , 
            n14949, \Ki[8] , n14948, \Ki[7] , n14947, \Ki[6] , n14946, 
            \Ki[5] , n14945, \Ki[4] , n14944, \Ki[3] , n14943, \Ki[2] , 
            n14942, \Ki[1] , n14941, \Kp[15] , n14940, \Kp[14] , 
            n14939, \Kp[13] , n14938, \Kp[12] , n14937, \Kp[11] , 
            n14936, \Kp[10] , n14935, \Kp[9] , n14934, \Kp[8] , 
            n14933, \Kp[7] , n14932, \Kp[6] , n14931, \Kp[5] , n14930, 
            \Kp[4] , n14929, \Kp[3] , n14928, \Kp[2] , n14927, \Kp[1] , 
            n14926, n14925, n14924, n14923, n14922, n14921, n14920, 
            n14919, n14918, n14917, n14916, n14915, n14914, n14913, 
            n14912, n14911, n14910, n14909, n14908, n14907, n14906, 
            n14905, n14904, n14903, n14902, n14901, \displacement[1] , 
            n14900, n14899, n14898, n14897, n14896, n14895, n14894, 
            n14893, n14892, n14891, n14890, n14889, n14888, n14887, 
            n14886, n26856, n26880, r_SM_Main, \r_SM_Main_2__N_3333[1] , 
            tx_o, n14872, VCC_net, \r_Bit_Index[0] , n7375, n14835, 
            n4_adj_4, n30875, tx_enable, n14672, n14766, \r_SM_Main_2__N_3262[2] , 
            r_SM_Main_adj_12, n26029, r_Rx_Data, RX_N_2, \r_Bit_Index[0]_adj_8 , 
            n13551, n4_adj_9, n15342, n25777, n15346, n18789, n4_adj_10, 
            n4_adj_11, n13556, n14826, n14825, n14824, n14823, n14822, 
            n14821, n14820) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [7:0]\data_out_frame[25] ;
    output [7:0]rx_data;
    output [23:0]setpoint;
    input clk32MHz;
    input n14885;
    output [23:0]IntegralLimit;
    input n14884;
    input n14883;
    output n10896;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output n4141;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    input n14882;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[8] ;
    input n14881;
    input n14880;
    input n14879;
    output [7:0]\data_in_frame[5] ;
    input n14878;
    output [7:0]\data_in_frame[4] ;
    input n14877;
    input n14876;
    output rx_data_ready;
    input n14875;
    input n14874;
    output [7:0]\data_out_frame[15] ;
    input n14873;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[24] ;
    output n2252;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    output n63;
    output n3;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[13] ;
    output \FRAME_MATCHER.state_31__N_2380[2] ;
    output [7:0]\data_in_frame[12] ;
    output n4137;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[8] ;
    output \data_out_frame[27][0] ;
    output n4;
    output tx_active;
    output n14641;
    output n24343;
    output n1;
    output DE_c;
    output n26748;
    output n7;
    output n7_adj_3;
    output LED_c;
    output n5;
    output n26399;
    input n14833;
    output [23:0]PWMLimit;
    input n14832;
    output [7:0]control_mode;
    input n28285;
    input n30820;
    input n15337;
    input n15336;
    input n15335;
    input n15334;
    input n15333;
    input n15332;
    input n15331;
    input n15330;
    input n15329;
    input n15328;
    input n15327;
    input n15326;
    input n15325;
    input n15324;
    input n15323;
    input n15322;
    input n15321;
    input n15320;
    input n15319;
    input n15318;
    input n15317;
    input n15316;
    input n15315;
    input n15314;
    input n15313;
    input n15312;
    input n15311;
    input n15310;
    input n15309;
    input n15308;
    input n15132;
    output [23:0]neopxl_color;
    input n15131;
    input n15130;
    input n15129;
    input n15128;
    input n15127;
    input n15126;
    input n15125;
    input n15124;
    input n15123;
    input n15122;
    input n15121;
    input n15120;
    input n15119;
    input n15118;
    input n15117;
    input n15116;
    input n15115;
    input n15114;
    input n15113;
    input n15112;
    input n15111;
    input n15110;
    input n15109;
    input n15108;
    input n15107;
    input n15106;
    input n15105;
    input n15104;
    input n15103;
    input n15102;
    input n15101;
    input n15100;
    input n15099;
    input n15098;
    input n15097;
    input n15096;
    input n15095;
    input n15094;
    input n15093;
    input n15092;
    input n15091;
    input n15090;
    input n15089;
    input n15088;
    input n15087;
    input n15086;
    input n15085;
    input n15084;
    input n15083;
    input n15082;
    input n15081;
    input n15080;
    input n15079;
    input n15077;
    input n15076;
    input n15075;
    input n15074;
    input n15073;
    input n15072;
    input n15071;
    input n15070;
    input n15069;
    input n15068;
    input n15067;
    input n15066;
    input n15065;
    input n15064;
    input n15063;
    input n15062;
    input n15061;
    input n15060;
    input n15059;
    input n15058;
    input n15057;
    input n15056;
    input n15055;
    input n15054;
    input n15053;
    input n15052;
    input n15051;
    input n15050;
    input n15049;
    input n15048;
    input n15047;
    input n15046;
    input n15045;
    input n15044;
    input n15043;
    input n15042;
    input n15041;
    input n15040;
    input n15039;
    input n15038;
    input n15037;
    input n15036;
    input n15035;
    input n15034;
    input n15033;
    input n15032;
    input n15031;
    input n15030;
    input n15029;
    input n15028;
    input n15027;
    input n15026;
    input n15025;
    input n15024;
    input n15023;
    input n15022;
    input n15021;
    input n15020;
    output n27156;
    input n15019;
    input n15018;
    input n15017;
    input n15016;
    input n15015;
    input n15014;
    input n15013;
    input n15012;
    input n15011;
    input n15010;
    input n15009;
    input n15008;
    input n15007;
    input n15006;
    input n15005;
    input n15004;
    input n15003;
    input n15002;
    input n15001;
    input n15000;
    input n14999;
    input n14998;
    input n14997;
    input n14996;
    input n14995;
    input n14994;
    input n14993;
    input n14992;
    input n14991;
    input n14990;
    input n14989;
    input n14830;
    input n14829;
    output \Ki[0] ;
    input n14828;
    output \Kp[0] ;
    input n14827;
    input n14988;
    input n14987;
    input n14986;
    input n14985;
    input n14984;
    input n14983;
    input n14982;
    input n14818;
    input n14981;
    input n14980;
    input n14979;
    input n14978;
    input n14977;
    input n14976;
    input n14975;
    input n14974;
    input n14973;
    input n14972;
    input n14971;
    input n14970;
    input n14969;
    input n14968;
    input n14967;
    input n14966;
    input n14965;
    input n14964;
    input n14963;
    input n14962;
    input n14961;
    input n14960;
    input n14959;
    input n14958;
    input n14957;
    input n14956;
    output \Ki[15] ;
    input n14955;
    output \Ki[14] ;
    input n14954;
    output \Ki[13] ;
    input n14953;
    output \Ki[12] ;
    input n14952;
    output \Ki[11] ;
    input n14951;
    output \Ki[10] ;
    input n14950;
    output \Ki[9] ;
    input n14949;
    output \Ki[8] ;
    input n14948;
    output \Ki[7] ;
    input n14947;
    output \Ki[6] ;
    input n14946;
    output \Ki[5] ;
    input n14945;
    output \Ki[4] ;
    input n14944;
    output \Ki[3] ;
    input n14943;
    output \Ki[2] ;
    input n14942;
    output \Ki[1] ;
    input n14941;
    output \Kp[15] ;
    input n14940;
    output \Kp[14] ;
    input n14939;
    output \Kp[13] ;
    input n14938;
    output \Kp[12] ;
    input n14937;
    output \Kp[11] ;
    input n14936;
    output \Kp[10] ;
    input n14935;
    output \Kp[9] ;
    input n14934;
    output \Kp[8] ;
    input n14933;
    output \Kp[7] ;
    input n14932;
    output \Kp[6] ;
    input n14931;
    output \Kp[5] ;
    input n14930;
    output \Kp[4] ;
    input n14929;
    output \Kp[3] ;
    input n14928;
    output \Kp[2] ;
    input n14927;
    output \Kp[1] ;
    input n14926;
    input n14925;
    input n14924;
    input n14923;
    input n14922;
    input n14921;
    input n14920;
    input n14919;
    input n14918;
    input n14917;
    input n14916;
    input n14915;
    input n14914;
    input n14913;
    input n14912;
    input n14911;
    input n14910;
    input n14909;
    input n14908;
    input n14907;
    input n14906;
    input n14905;
    input n14904;
    input n14903;
    input n14902;
    input n14901;
    input \displacement[1] ;
    input n14900;
    input n14899;
    input n14898;
    input n14897;
    input n14896;
    input n14895;
    input n14894;
    input n14893;
    input n14892;
    input n14891;
    input n14890;
    input n14889;
    input n14888;
    input n14887;
    input n14886;
    output n26856;
    output n26880;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3333[1] ;
    output tx_o;
    input n14872;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n7375;
    input n14835;
    output n4_adj_4;
    input n30875;
    output tx_enable;
    output n14672;
    output n14766;
    output \r_SM_Main_2__N_3262[2] ;
    output [2:0]r_SM_Main_adj_12;
    input n26029;
    output r_Rx_Data;
    input RX_N_2;
    output \r_Bit_Index[0]_adj_8 ;
    output n13551;
    output n4_adj_9;
    input n15342;
    input n25777;
    input n15346;
    output n18789;
    output n4_adj_10;
    output n4_adj_11;
    output n13556;
    input n14826;
    input n14825;
    input n14824;
    input n14823;
    input n14822;
    input n14821;
    input n14820;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n17125, n17129, n7_c, n24756, n26377, n27865, n27162, 
        n26136, n26476;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n18, n19251, n26035;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n15193;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n2272, n3_c, n3_adj_3581, n3_adj_3582, n3_adj_3583, n3_adj_3584, 
        n3_adj_3585, n3939, n14593, n2, n3_adj_3586, n3_adj_3587, 
        n21982, n21983, n3_adj_3588, n3_adj_3589, n3_adj_3590, n3_adj_3591, 
        n3_adj_3592, n3_adj_3593, n3_adj_3594, n3_adj_3595, n3_adj_3596;
    wire [31:0]\FRAME_MATCHER.state_31__N_2444 ;
    
    wire n19405, n3_adj_3597, n3_adj_3598, n3_adj_3599, n3_adj_3600, 
        n3_adj_3601, n3_adj_3602, n3_adj_3603, n3_adj_3604, n3_adj_3605, 
        n3_adj_3606, n3_adj_3607, n3_adj_3608, n3_adj_3609, n3_adj_3610, 
        n3_adj_3611;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n3938, n3962, n3961, n3960, n3959, n3958, n3957, n3956, 
        n3955;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n3954, n3953, n3952, n25968, n31, n6, n3951, n4_c, 
        n3950, n3949, n3948, n3947;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n3946, n3945, n3944, n3943, n3942, n3941, n3940;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n29240, n29239, n16, n17, n29237, n29236, n16_adj_3612, 
        n17_adj_3613, n29230, n29229, n16_adj_3614, n17_adj_3615, 
        n29224, n29223, n16_adj_3616, n17_adj_3617, n29221, n29220, 
        n16_adj_3618, n17_adj_3619, n29218, n29217, n6_adj_3620, n5_c, 
        n29157, n7_adj_3621, n30448, n30436, n14, n30502, n29216, 
        n6_adj_3622, n5_adj_3623, n7_adj_3624, n30442, n30478, n14_adj_3625, 
        n30508, n29219, n6_adj_3626, n5_adj_3627, n7_adj_3628, n30430, 
        n30346, n14_adj_3629, n30286, n29222, n2_adj_3630, n21981, 
        n1656, n16_adj_3631, n17_adj_3632, n29227, n29226, n15194, 
        n15195, n8, n15180, n29573, n5_adj_3633, n7_adj_3634, n30424, 
        n30550, n14_adj_3635, n30292, n29225, n29567, n5_adj_3636, 
        n7_adj_3637, n30418, n30568, n14_adj_3638, n30298, n29228, 
        n6_adj_3639, n5_adj_3640, n7_adj_3641, n30412, n30394, n14_adj_3642, 
        n30322, n29231, n29545, n5_adj_3643, n7_adj_3644, n15181, 
        n30472, n30382, n14_adj_3645, n30340, n29238, n15182, n23683, 
        n26389, n29590, n5_adj_3646, n7_adj_3647, n30466, n30454, 
        n14_adj_3648, n30490, n29274;
    wire [7:0]\data_out_frame[20]_c ;   // verilog/coms.v(97[12:26])
    
    wire n8_adj_3649, n30496, n29799, n15183, n15184, n15185, n15186, 
        n15187, n14279, n26482, n26157, n14273, n8_adj_3650, n15172, 
        n15173, n28358, n28168;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n24052, n26, n15174, n15175, n24618, n27443, n13813, 
        n6_adj_3651, Kp_23__N_656, n28018, n26262, n22, n15176, 
        n28354, n26964, n26206, n28380, n27416, n26624, n21, n27369, 
        n29, n26145, n6_adj_3652, n14111, n31_adj_3653, n15177, 
        n15178, n15179, n14192, n26113, Kp_23__N_816, n10649, n26353, 
        n26256, n23699, n24006;
    wire [0:0]n2786;
    wire [2:0]r_SM_Main_2__N_3336;
    
    wire n26052, n2_adj_3654, n21980, \FRAME_MATCHER.rx_data_ready_prev , 
        n25509, n25725;
    wire [7:0]n8825;
    
    wire n14614, n14738, n26102, n26674, n26464, n14_adj_3655, n6_adj_3656, 
        n26486, n10, n26116, n26110, n24620, n24605, n23661, n26373, 
        n24770, n26303, n26568, n26402, n26347, n24737, n13970, 
        n10_adj_3657, n27637, n24614, n26413, n2_adj_3658, n21979, 
        n26269, n27993, n26442, n24722, n26099, n2_adj_3659, n21978, 
        n2_adj_3660, n21977, n27795, n23765, n27602, n13816, n23877, 
        n27731, n26217, n23715, n26350, n3_adj_3661, n26074, n25549, 
        n25555, n25561, n25567, n25573, n25579, n25585, n25591, 
        n25597, n25603, n25609, n25631, n25643;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n6_adj_3662, n25521, n2_adj_3663, n2_adj_3664, n25695, n8_adj_3665, 
        n13538, n4452, n25671, n25693, n25691, n25689, n8_adj_3666, 
        n15164, n18723, n18721, n15165, n15166, n13503, n15, n1_c, 
        n15167, n18719, n13541, n13535, n18_adj_3667, n25687, n28376, 
        n12, n17879, n10_adj_3668, n15168, n23166, n25685, n2_adj_3669, 
        n21976, n97, n22005, n10_adj_3670, n18_adj_3671, n16_adj_3672, 
        n20, n13402, n14_adj_3673, n9, n7_adj_3674, n16_adj_3675, 
        n17_adj_3676, n25683, n63_c, n7_adj_3677, n18_adj_3678, n2_adj_3679, 
        n21975, n28382, n25681, n12_adj_3680, n63_adj_3681, n82, 
        n22004, n5_adj_3682, n771, n18717, n7_adj_3683, n18713, 
        n8604;
    wire [31:0]\FRAME_MATCHER.state_31__N_2380 ;
    
    wire n7_adj_3684, n88, n28, n26_adj_3686, n27, n25, n28207, 
        n18_adj_3687, n25679, n16_adj_3688, n7_adj_3689, n20_adj_3690, 
        n25677, n13372, n15169, n8_adj_3691, n3303, n25675, n25673, 
        n2_adj_3692, n21974, n7_adj_3693, n15170, n4_adj_3695, n25663, 
        n7_adj_3696, n15171, n25669, n101, n112, n25481, n8_adj_3697, 
        n15156, n22003, n15157, n19229, n15158, n26154, n13826, 
        n130, n2_adj_3698, n23168, n27344, tx_transmit_N_3233, n19227, 
        n26051, n13, n29270, n15159, n19225, n22002, n8_adj_3699, 
        n15160, n15161, n8_adj_3700, n23172, n8_adj_3701, n8_adj_3702, 
        n2_adj_3703, n21973, n8_adj_3704, n22001, n19223, n25459, 
        n8_adj_3705, n26334, n26544;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n26380, n13_adj_3706, n15162, n26362, n18732, n26044, n14289, 
        n26500, n34, n39, n2_adj_3707, n21972, n15163, n8_adj_3708, 
        n15148, n83, n13604, n15149, n26278, Kp_23__N_650, n15150, 
        n2_adj_3709, n21971, n22000, n15151, n26209, n14224, n6_adj_3710, 
        Kp_23__N_915, n26244, n6_adj_3711, n15152, n6_adj_3712, n15153, 
        n14294, n15154, n12779, n10_adj_3713, Kp_23__N_708, n23701, 
        n26457, n14403, n26106, n28350, n2_adj_3714, n21970, n8_adj_3715, 
        n15155;
    wire [31:0]n92;
    
    wire n8_adj_3716, n15140, n26559, n26581, n26343, n26649, n10_adj_3717, 
        n14_adj_3718;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n26636, n9_adj_3719, n24641, n23804, n26405, n7_adj_3720, 
        n15141, n17197, n17173, n21999, n26571, n26214, n6_adj_3721, 
        Kp_23__N_1026, n26526, n26547, n15142, n26445, n26645, n14149, 
        n14429, n23657, n10_adj_3722, n14_adj_3723, n26596, n24179, 
        n27569, n23779, n26203, n26190, n24616, n28_adj_3724, n26259, 
        n26655, n26_adj_3725, n23828, n26609, n26689, n27_adj_3726, 
        n26699, n25_adj_3727, n26565, n27426, n10_adj_3728, n23841, 
        Kp_23__N_1237, n24653, n6_adj_3729, n24728, n26409, n26337, 
        n24735, n24639, n26421, n13253, n14315, n26275, n26395, 
        n10_adj_3730, n13670, n14309, n24637, n23621, n26418, n13882, 
        n13890, n23477, n26529, n15_adj_3731, n14_adj_3732, n14098, 
        n6_adj_3733, n26340, n24599, n10_adj_3734, n4_adj_3735, n26132, 
        n15133, n14503, n26415, n23681, n15134, n15135, n15136, 
        n10_adj_3736, n15137, n15138, n15139, n4_adj_3737, n20_adj_3738, 
        n28_adj_3739, n26184, n12_adj_3740, n24659, n26_adj_3741, 
        n13685, n26196, n14140, n27_adj_3742, n26180, n24719, n25_adj_3743, 
        n11166, n26492, n6_adj_3744, n26033, n18_adj_3745, n14831, 
        n24635, n26556, n16_adj_3746, n20_adj_3747, n26057, n26079, 
        n6_adj_3748, n26129, n14432, n18866, n10_adj_3749, n26233, 
        n10_adj_3750, n21564, n6_adj_3751, n14524, n2_adj_3752, n14_adj_3753, 
        n10_adj_3754, n13915, n26250, n13804, n26272, n16570, n24622, 
        n11, n14196, n15143, n9_adj_3755, n12_adj_3756, n2_adj_3757, 
        n21969, n26170, n10_adj_3758, Kp_23__N_1002, n26630, n23794, 
        n13867, n26089, n26140, n12_adj_3759, n23664, n26587, Kp_23__N_1256, 
        n26671, n26575, n14_adj_3760, n10_adj_3761, n26658, n26590, 
        n14_adj_3762, n10_adj_3763, n23708, n42, n26308, n24689, 
        n57, n36, n26328, n26_adj_3764, n40, n38, n15144, n26652, 
        n26423, n37, n27143, n66, n64, n38_adj_3765, n65, n26520, 
        n63_adj_3766, n60, n43, n14485, n62, n26517, n61, n72, 
        n24414, n67, n24206, n13719, n14_adj_3767, n26292, n13904, 
        n26553, n8_adj_3768, n26436, n6_adj_3769, n27074, n26227, 
        n13921, n10_adj_3770, n26086, n14_adj_3771, n26247, n12_adj_3772, 
        Kp_23__N_1283, n14152, n12_adj_3773, n26541, n26433, n12002, 
        n14_adj_3774, n10_adj_3775, n26661, n26693, n26538, n8_adj_3776, 
        n26480, n26331, n10_adj_3777, n8_adj_3778, n12_adj_3779, n27630, 
        n12_adj_3780, n14_adj_3781, n9_adj_3782, n30565, n30559;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n30304, n30553, n30547, n30310, n30541, n30316, n30535, 
        n30526, n30529, n30523, n133, n27310, n30328, n30517, 
        n27889, n14_adj_3783, n4_adj_3784, n26987, n30334, n30511;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n30505, n30499, n6_adj_3785, n30493, n30487, n30475, n26495, 
        n10_adj_3786, n30469, n30463, n30451, n30445, n13178, n4_adj_3787, 
        n30439, n14_adj_3788, n30433, n26677, n30427, n26454, n30421, 
        n30415, n30409, n26151, n26164, n30391, n14446, n26461, 
        n30379, n6_adj_3789, n30352, n30361, n2_adj_3790, n21998, 
        n30349, n30343, n30, n30337, n34_adj_3791, n30331, n32, 
        n30325, n33, n30319, n31_adj_3792, n30313, n30307, n30301, 
        n15300, n15301, n2_adj_3793, n2_adj_3794, n21997, n15302, 
        n15303, n15304, n15305, n15306, n15307, n15145, n13998, 
        n14360, n23654, n807, n2_adj_3796, n2_adj_3797, n2_adj_3798, 
        n2_adj_3799, n2_adj_3800, n2_adj_3801, n2_adj_3802, n2_adj_3803, 
        n2_adj_3804, n2_adj_3805, n2_adj_3806, n2_adj_3807, n2_adj_3808, 
        n2_adj_3809, n2_adj_3810, n21968, n17_adj_3811, n16_adj_3812, 
        n4_adj_3813, n15292, n15146, n28031, n27106, n27586, n26125, 
        n27190, n26401, n27494, n26427, n26524, n26255, n27842, 
        n15293, n15147, n15294, n161, n13872, n15295, n15296, 
        n25515, n25667, n15297, n15298, n15299, n62_adj_3815, n27319, 
        n135, n26359, n6_adj_3816, n14002, n10_adj_3817, n6_adj_3818, 
        n26467, n10_adj_3819, n26167, n21996, n26126, n26120, n6_adj_3820, 
        n6_adj_3821, n26287, n26323, n11_adj_3822, n6_adj_3823, n26448, 
        n26223, n13990, n23458, n26367, n7_adj_3824, n27708, n14506, 
        n27647, n23796, n26535, n8_adj_3826, n15284, n15285, n15286, 
        n15287, n10_adj_3827, n27710, n26426, n15288, n24055, n27908, 
        n26253, n15289, n24632, n15290, n15291, n60_adj_3828, n21995, 
        n30295, n21994, n15276, n24657, n8_adj_3830, n15277, n26489, 
        n15278, n15279, n15280, n15281, n28332, n30_adj_3831, n28_adj_3832, 
        n29_adj_3833, n27_adj_3834, n15282, n28244, n15283, n21993, 
        n15268, n15269, n15270, n15271, n15272, n15273, n15274, 
        n15275, n23800, n23771, n26523, n15260, n26508, n24645, 
        n26281, n26284, n26230, n10_adj_3836, n26386, n26174, n13291, 
        n13_adj_3837, n26175, n15261, n26297, n13221, n15262, n26593, 
        n52, n59, n26696, n24630, n26642, n56, n26633, n26702, 
        n26502, n54, n26241, n14240, n23824, n55, n15263, n26356, 
        n26683, n53, n26236, n26093, n58, n64_adj_3838, n57_adj_3839, 
        n65_adj_3840, n13726, n15264, n26187, n8_adj_3841, n12_adj_3842, 
        n26_adj_3843, n24375, n23761, n15265, n12_adj_3844, n15266, 
        n48, n26562, n46, n26300, n47, n26314, n45, n15267, 
        n26289, n44, n43_adj_3845, n21992, n15252, n15253, n15254, 
        n54_adj_3846, n49, n15255, n21991, n15256, n14501, n24674, 
        n27564, n26123, n15257, n15258, n24601, n26550, n15259, 
        n15244, n24607, n21990, n15245, n15251, n15250, n15249, 
        n26317, n15246, n14336, n26505, n8_adj_3847, n13788, n7_adj_3848, 
        n15248, n15247, n15243, n15242, n15241, n15240, n15239, 
        n15238, n15237, n15236, n15235, n15234, n15233, n15232, 
        n15231, n15230, n15229, n15228, n15227, n15226, n15225, 
        n15224, n15223, n15222, n15221, n15220, n15219, n15218, 
        n15217, n15216, n15215, n15214, n15213, n15212, n15211, 
        n15210, n15209, n15208, n15207, n15206, n15205, n15204, 
        n15203, n15202, n15201, n15200, n15199, n15198, n15197, 
        n15196, n15192, n15191, n15190, n15189, n15188, n26680, 
        n26615, n15_adj_3849, n13974, n12_adj_3850, n4_adj_3851, n26600, 
        n12_adj_3852, n12_adj_3853, n26668, n13_adj_3854, n30289, 
        n28172, n26311, n13236, n26621, n26320, n15078, n7_adj_3855, 
        n26532, n21989, n14011, n14_adj_3856, n15_adj_3857, n26618, 
        n14_adj_3858, n24314, n26200, n21988, n26639, n26470, n8_adj_3859, 
        n24463, n7_adj_3860, n8_adj_3861, n26193, n6_adj_3862, n26511, 
        n16_adj_3863, n26584, n26686, n17_adj_3864, n27507, n26603, 
        n14_adj_3865, n26083, n21987, n26665, n8_adj_3866, n21986, 
        n26211, n12_adj_3867, n26612, n10_adj_3868, n30283, n6_adj_3869, 
        n26514, n21985, n12_adj_3870, n21984, n15_adj_3871;
    
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n17125), .I2(GND_net), 
            .I3(GND_net), .O(n17129));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(n7_c), .I1(\data_out_frame[25] [7]), .I2(n24756), 
            .I3(n26377), .O(n27865));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(n27162), .I1(n26136), .I2(n26476), .I3(\data_in_frame[20] [5]), 
            .O(n18));
    defparam i2_4_lut.LUT_INIT = 16'hbeeb;
    SB_LUT4 i11388_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n15193));
    defparam i11388_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_292_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_c));
    defparam select_292_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3581));
    defparam select_292_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3582));
    defparam select_292_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3583));
    defparam select_292_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3584));
    defparam select_292_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3585));
    defparam select_292_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n14593), .D(n3939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n14885));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_292_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3587));
    defparam select_292_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_17 (.CI(n21982), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n21983));
    SB_LUT4 select_292_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3588));
    defparam select_292_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3589));
    defparam select_292_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3590));
    defparam select_292_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3591));
    defparam select_292_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3592));
    defparam select_292_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3593));
    defparam select_292_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n14884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n14883));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_292_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3594));
    defparam select_292_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3595));
    defparam select_292_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3596));
    defparam select_292_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(\FRAME_MATCHER.state_31__N_2444 [3]), .I1(n19405), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n10896));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 select_292_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3597));
    defparam select_292_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3598));
    defparam select_292_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3599));
    defparam select_292_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3600));
    defparam select_292_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3601));
    defparam select_292_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3602));
    defparam select_292_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3603));
    defparam select_292_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3604));
    defparam select_292_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3605));
    defparam select_292_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3606));
    defparam select_292_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3607));
    defparam select_292_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3608));
    defparam select_292_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3609));
    defparam select_292_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3610));
    defparam select_292_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_292_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3611));
    defparam select_292_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_984_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n3938), .I3(GND_net), .O(n3962));
    defparam mux_984_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n3938), .I3(GND_net), .O(n3961));
    defparam mux_984_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n3938), .I3(GND_net), .O(n3960));
    defparam mux_984_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n3938), .I3(GND_net), .O(n3959));
    defparam mux_984_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n3938), .I3(GND_net), .O(n3958));
    defparam mux_984_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n3938), .I3(GND_net), .O(n3957));
    defparam mux_984_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n3938), .I3(GND_net), .O(n3956));
    defparam mux_984_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n3938), .I3(GND_net), .O(n3955));
    defparam mux_984_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n3938), .I3(GND_net), .O(n3954));
    defparam mux_984_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_292_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2272), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3586));
    defparam select_292_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_984_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n3938), .I3(GND_net), .O(n3953));
    defparam mux_984_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n3938), .I3(GND_net), .O(n3952));
    defparam mux_984_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_836 (.I0(n25968), .I1(n31), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i1_2_lut_adj_836.LUT_INIT = 16'h2222;
    SB_LUT4 mux_984_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n3938), .I3(GND_net), .O(n3951));
    defparam mux_984_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_837 (.I0(\FRAME_MATCHER.state [2]), .I1(n17129), 
            .I2(n4_c), .I3(n6), .O(n4141));
    defparam i4_4_lut_adj_837.LUT_INIT = 16'h0200;
    SB_LUT4 mux_984_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n3938), .I3(GND_net), .O(n3950));
    defparam mux_984_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n3938), .I3(GND_net), .O(n3949));
    defparam mux_984_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n3938), .I3(GND_net), .O(n3948));
    defparam mux_984_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n3938), .I3(GND_net), .O(n3947));
    defparam mux_984_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n3938), .I3(GND_net), .O(n3946));
    defparam mux_984_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n3938), .I3(GND_net), .O(n3945));
    defparam mux_984_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n3938), .I3(GND_net), .O(n3944));
    defparam mux_984_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n3938), .I3(GND_net), .O(n3943));
    defparam mux_984_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n3938), .I3(GND_net), .O(n3942));
    defparam mux_984_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n3938), .I3(GND_net), .O(n3941));
    defparam mux_984_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_984_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n3938), .I3(GND_net), .O(n3940));
    defparam mux_984_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24480_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29240));
    defparam i24480_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24483_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29239));
    defparam i24483_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24496_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29237));
    defparam i24496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24286_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29236));
    defparam i24286_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3612));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3613));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24501_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29230));
    defparam i24501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24505_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29229));
    defparam i24505_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3614));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3615));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24511_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29224));
    defparam i24511_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24513_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29223));
    defparam i24513_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12778_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n16_adj_3616));   // verilog/coms.v(102[12:33])
    defparam i12778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3617));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24516_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29221));
    defparam i24516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24518_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29220));
    defparam i24518_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3618));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3619));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24520_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29218));
    defparam i24520_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24522_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29217));
    defparam i24522_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3620));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hb0b3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut (.I0(n5_c), .I1(n6_adj_3620), 
            .I2(n29157), .I3(GND_net), .O(n7_adj_3621));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1568646_i1_3_lut (.I0(n30448), .I1(n30436), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14));
    defparam i1568646_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24247_2_lut (.I0(n30502), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29216));
    defparam i24247_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3622));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3623));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_adj_3623), 
            .I1(n6_adj_3622), .I2(n29157), .I3(GND_net), .O(n7_adj_3624));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1569249_i1_3_lut (.I0(n30442), .I1(n30478), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3625));
    defparam i1569249_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24521_2_lut (.I0(n30508), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29219));
    defparam i24521_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3626));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3627));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_3627), 
            .I1(n6_adj_3626), .I2(n29157), .I3(GND_net), .O(n7_adj_3628));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1569852_i1_3_lut (.I0(n30430), .I1(n30346), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3629));
    defparam i1569852_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24517_2_lut (.I0(n30286), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29222));
    defparam i24517_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_43_16_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n21981), .O(n2_adj_3630)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n14882));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3631));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3632));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24507_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29227));
    defparam i24507_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24510_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29226));
    defparam i24510_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11389_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n15194));
    defparam i11389_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11390_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n15195));
    defparam i11390_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11375_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n15180));
    defparam i11375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n29573));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3633));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_3633), 
            .I1(byte_transmit_counter[0]), .I2(n29157), .I3(n29573), .O(n7_adj_3634));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1570455_i1_3_lut (.I0(n30424), .I1(n30550), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3635));
    defparam i1570455_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24512_2_lut (.I0(n30292), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29225));
    defparam i24512_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24502_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29567));   // verilog/coms.v(106[34:55])
    defparam i24502_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3636));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_3636), 
            .I1(n29567), .I2(n29157), .I3(byte_transmit_counter[0]), .O(n7_adj_3637));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1571058_i1_3_lut (.I0(n30418), .I1(n30568), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3638));
    defparam i1571058_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24509_2_lut (.I0(n30298), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29228));
    defparam i24509_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i6_3_lut (.I0(\data_out_frame[5] [7]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n6_adj_3639));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3640));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut (.I0(n5_adj_3640), 
            .I1(n6_adj_3639), .I2(n29157), .I3(GND_net), .O(n7_adj_3641));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1571661_i1_3_lut (.I0(n30412), .I1(n30394), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3642));
    defparam i1571661_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24504_2_lut (.I0(n30322), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29231));
    defparam i24504_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_3_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n29545));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3643));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_4_lut (.I0(n5_adj_3643), 
            .I1(byte_transmit_counter[0]), .I2(n29157), .I3(n29545), .O(n7_adj_3644));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i11376_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n15181));
    defparam i11376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1572867_i1_3_lut (.I0(n30472), .I1(n30382), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3645));
    defparam i1572867_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24497_2_lut (.I0(n30340), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29238));
    defparam i24497_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_16 (.CI(n21981), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n21982));
    SB_LUT4 i11377_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n15182));
    defparam i11377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_838 (.I0(\data_in_frame[8] [1]), .I1(n23683), .I2(GND_net), 
            .I3(GND_net), .O(n26389));
    defparam i1_2_lut_adj_838.LUT_INIT = 16'h6666;
    SB_LUT4 i24073_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n29157));   // verilog/coms.v(106[34:55])
    defparam i24073_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24524_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n29590));   // verilog/coms.v(106[34:55])
    defparam i24524_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3646));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_4_lut (.I0(n5_adj_3646), 
            .I1(n29590), .I2(n29157), .I3(byte_transmit_counter[0]), .O(n7_adj_3647));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_4_lut.LUT_INIT = 16'haca0;
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n14881));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1568043_i1_3_lut (.I0(n30466), .I1(n30454), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3648));
    defparam i1568043_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24262_2_lut (.I0(n30490), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29274));   // verilog/coms.v(106[34:55])
    defparam i24262_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[20]_c [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(byte_transmit_counter[1]), 
            .O(n8_adj_3649));   // verilog/coms.v(106[34:55])
    defparam i22_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i24733_3_lut (.I0(n30496), .I1(n8_adj_3649), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n29799));
    defparam i24733_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n14880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n14879));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11378_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n15183));
    defparam i11378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11379_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n15184));
    defparam i11379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11380_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n15185));
    defparam i11380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11381_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n15186));
    defparam i11381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11382_3_lut_4_lut (.I0(n8), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n15187));
    defparam i11382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut (.I0(n14279), .I1(n26482), .I2(n26157), .I3(\data_in_frame[1] [6]), 
            .O(n14273));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11367_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n15172));
    defparam i11367_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11368_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n15173));
    defparam i11368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut (.I0(n28358), .I1(n28168), .I2(\data_in_frame[21] [1]), 
            .I3(n24052), .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'h7ff7;
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n14878));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11369_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n15174));
    defparam i11369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11370_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n15175));
    defparam i11370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_839 (.I0(\data_in_frame[21] [0]), .I1(n24052), 
            .I2(n24618), .I3(GND_net), .O(n27443));
    defparam i2_3_lut_adj_839.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_840 (.I0(\data_in_frame[1] [5]), .I1(n13813), .I2(\data_in_frame[3] [7]), 
            .I3(n6_adj_3651), .O(Kp_23__N_656));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_840.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n28018), .I1(\data_in_frame[21] [2]), .I2(n26262), 
            .I3(n24618), .O(n22));
    defparam i6_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i11371_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n15176));
    defparam i11371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23317_4_lut (.I0(\data_in_frame[21] [4]), .I1(n28354), .I2(n26964), 
            .I3(n26206), .O(n28380));
    defparam i23317_4_lut.LUT_INIT = 16'h4080;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[20] [4]), .I1(n27416), .I2(n26476), 
            .I3(n26624), .O(n21));
    defparam i5_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i13_4_lut (.I0(n27443), .I1(n26), .I2(n18), .I3(n27369), 
            .O(n29));
    defparam i13_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i4_4_lut_adj_841 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[4] [3]), 
            .I2(n26145), .I3(n6_adj_3652), .O(n14111));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_841.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n29), .I1(n21), .I2(n28380), .I3(n22), .O(n31_adj_3653));
    defparam i15_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i11372_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n15177));
    defparam i11372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11373_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n15178));
    defparam i11373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11374_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n15179));
    defparam i11374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_842 (.I0(n14192), .I1(n26113), .I2(\data_in_frame[4] [3]), 
            .I3(GND_net), .O(Kp_23__N_816));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_842.LUT_INIT = 16'h9696;
    SB_LUT4 i1571_3_lut (.I0(n31_adj_3653), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n10649));
    defparam i1571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_843 (.I0(n26353), .I1(n26256), .I2(\data_in_frame[1] [4]), 
            .I3(n23699), .O(n24006));
    defparam i3_4_lut_adj_843.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n14877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n14876));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3336[0]), .C(clk32MHz), 
            .D(n2786[0]), .R(n26052));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_15_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n21980), .O(n2_adj_3654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
            .D(n25509), .S(n25725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n14875));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n14614), .D(n8825[7]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n14874));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(n26102), .O(n26674));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(n26464), .I3(\data_out_frame[15] [7]), .O(n14_adj_3655));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_844 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[7] [0]), 
            .I2(\data_in_frame[4] [4]), .I3(n6_adj_3656), .O(n26486));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_844.LUT_INIT = 16'h6996;
    SB_CARRY add_43_15 (.CI(n21980), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n21981));
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n14873));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[12] [2]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n10));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_845 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[12] [2]), 
            .I2(\data_out_frame[10] [1]), .I3(n26116), .O(n26110));
    defparam i2_3_lut_4_lut_adj_845.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_846 (.I0(n24620), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[18] [6]), .I3(\data_out_frame[20] [7]), 
            .O(n24605));
    defparam i2_3_lut_4_lut_adj_846.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut (.I0(n23661), .I1(n26373), .I2(n24770), .I3(n26303), 
            .O(n26568));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(n23661), .I1(n26373), .I2(\data_out_frame[19] [6]), 
            .I3(GND_net), .O(n26402));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n14614), .D(n8825[6]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n14614), .D(n8825[5]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_847 (.I0(n23661), .I1(n26373), .I2(n26347), 
            .I3(GND_net), .O(n24737));
    defparam i1_2_lut_3_lut_adj_847.LUT_INIT = 16'h6969;
    SB_LUT4 i5_3_lut_4_lut_adj_848 (.I0(\data_out_frame[17] [6]), .I1(n13970), 
            .I2(\data_out_frame[15] [6]), .I3(n10_adj_3657), .O(n27637));
    defparam i5_3_lut_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_849 (.I0(\data_out_frame[17] [6]), .I1(n13970), 
            .I2(n24614), .I3(GND_net), .O(n26413));
    defparam i1_2_lut_3_lut_adj_849.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_14_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n21979), .O(n2_adj_3658)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_14 (.CI(n21979), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n21980));
    SB_LUT4 i1_2_lut_4_lut (.I0(n26269), .I1(\data_out_frame[9] [2]), .I2(n27993), 
            .I3(n26442), .O(n24722));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_850 (.I0(n26269), .I1(\data_out_frame[9] [2]), 
            .I2(n27993), .I3(\data_out_frame[13] [5]), .O(n26099));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_13_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n21978), .O(n2_adj_3659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_13 (.CI(n21978), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n21979));
    SB_LUT4 add_43_12_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n21977), .O(n2_adj_3660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_851 (.I0(n24737), .I1(n27795), .I2(n23765), 
            .I3(\data_out_frame[24] [3]), .O(n27602));
    defparam i2_3_lut_4_lut_adj_851.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_852 (.I0(n24737), .I1(n27795), .I2(n13816), 
            .I3(n23877), .O(n27731));
    defparam i2_3_lut_4_lut_adj_852.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_853 (.I0(n26217), .I1(n23715), .I2(\data_out_frame[23] [0]), 
            .I3(\data_out_frame[19] [0]), .O(n26350));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_853.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_854 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n25549));
    defparam i1_2_lut_3_lut_adj_854.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_855 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n25555));
    defparam i1_2_lut_3_lut_adj_855.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_856 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n25561));
    defparam i1_2_lut_3_lut_adj_856.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_857 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n25567));
    defparam i1_2_lut_3_lut_adj_857.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_858 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n25573));
    defparam i1_2_lut_3_lut_adj_858.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_859 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n25579));
    defparam i1_2_lut_3_lut_adj_859.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_860 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n25585));
    defparam i1_2_lut_3_lut_adj_860.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_861 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n25591));
    defparam i1_2_lut_3_lut_adj_861.LUT_INIT = 16'he0e0;
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n14614), .D(n8825[4]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_862 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n25597));
    defparam i1_2_lut_3_lut_adj_862.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_863 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n25603));
    defparam i1_2_lut_3_lut_adj_863.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_864 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n25609));
    defparam i1_2_lut_3_lut_adj_864.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_865 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n25631));
    defparam i1_2_lut_3_lut_adj_865.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_866 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n25643));
    defparam i1_2_lut_3_lut_adj_866.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_867 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3662));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_868 (.I0(n3_adj_3661), .I1(n26074), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n25521));
    defparam i1_2_lut_3_lut_adj_868.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_12 (.CI(n21977), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n21978));
    SB_LUT4 i1_2_lut_3_lut_adj_869 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [31]), .I3(GND_net), .O(n25695));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_869.LUT_INIT = 16'he0e0;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n14614), .D(n8825[3]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15002_4_lut (.I0(n8_adj_3665), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n13538), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i15002_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_3_lut_adj_870 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [30]), .I3(GND_net), .O(n25671));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_870.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_871 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [29]), .I3(GND_net), .O(n25693));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_871.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_872 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [28]), .I3(GND_net), .O(n25691));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_872.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_873 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [27]), .I3(GND_net), .O(n25689));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_873.LUT_INIT = 16'he0e0;
    SB_LUT4 i11359_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n15164));
    defparam i11359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_874 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [26]), .I3(GND_net), .O(n18723));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_874.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_875 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [25]), .I3(GND_net), .O(n18721));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_875.LUT_INIT = 16'he0e0;
    SB_LUT4 i11360_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n15165));
    defparam i11360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11361_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n15166));
    defparam i11361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_876 (.I0(n1656), .I1(n13503), .I2(n15), .I3(n1_c), 
            .O(n2252));
    defparam i3_4_lut_adj_876.LUT_INIT = 16'h0040;
    SB_LUT4 i11362_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n15167));
    defparam i11362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_877 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [24]), .I3(GND_net), .O(n18719));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_877.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut (.I0(n13541), .I1(\data_in[1] [6]), .I2(\data_in[0] [1]), 
            .I3(n13535), .O(n18_adj_3667));
    defparam i7_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_878 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [23]), .I3(GND_net), .O(n25687));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_878.LUT_INIT = 16'he0e0;
    SB_LUT4 i23313_4_lut (.I0(\data_in[2] [0]), .I1(\data_in[1] [3]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n28376));
    defparam i23313_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_879 (.I0(n28376), .I1(\data_in[2] [5]), .I2(n18_adj_3667), 
            .I3(n12), .O(n17879));
    defparam i10_4_lut_adj_879.LUT_INIT = 16'hfff7;
    SB_LUT4 i4_4_lut_adj_880 (.I0(\data_in[1] [0]), .I1(\data_in[0] [6]), 
            .I2(\data_in[1] [4]), .I3(\data_in[0] [3]), .O(n10_adj_3668));
    defparam i4_4_lut_adj_880.LUT_INIT = 16'hfdff;
    SB_LUT4 i11363_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n15168));
    defparam i11363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18116_2_lut_3_lut (.I0(n2_adj_3663), .I1(n2_adj_3664), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n23166));   // verilog/coms.v(115[11:12])
    defparam i18116_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_881 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [21]), .I3(GND_net), .O(n25685));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_881.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_11_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n21976), .O(n2_adj_3669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_882 (.I0(\data_in[3] [0]), .I1(\data_in[2] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n97));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_adj_882.LUT_INIT = 16'hdddd;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n22005), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_883 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3670));
    defparam i4_4_lut_adj_883.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut (.I0(\data_in[3] [4]), .I1(n10_adj_3670), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n13535));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i7_4_lut_adj_884 (.I0(\data_in[1] [3]), .I1(n13535), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n18_adj_3671));
    defparam i7_4_lut_adj_884.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(\data_in[3] [7]), .I1(\data_in[0] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_3672));
    defparam i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i9_4_lut (.I0(\data_in[0] [5]), .I1(n18_adj_3671), .I2(\data_in[2] [5]), 
            .I3(\data_in[2] [6]), .O(n20));
    defparam i9_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i10_4_lut_adj_885 (.I0(\data_in[1] [6]), .I1(n20), .I2(n16_adj_3672), 
            .I3(\data_in[2] [0]), .O(n13402));
    defparam i10_4_lut_adj_885.LUT_INIT = 16'hfffd;
    SB_LUT4 i6_4_lut_adj_886 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3673));
    defparam i6_4_lut_adj_886.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_887 (.I0(\data_in[3] [3]), .I1(\data_in[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_887.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_888 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [20]), .I3(GND_net), .O(n7_adj_3674));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_888.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_889 (.I0(n9), .I1(n14_adj_3673), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [1]), .O(n13541));
    defparam i7_4_lut_adj_889.LUT_INIT = 16'hffef;
    SB_LUT4 i6_4_lut_adj_890 (.I0(\data_in[2] [2]), .I1(\data_in[0] [6]), 
            .I2(n13541), .I3(n13402), .O(n16_adj_3675));
    defparam i6_4_lut_adj_890.LUT_INIT = 16'hfffb;
    SB_LUT4 i7_4_lut_adj_891 (.I0(\data_in[3] [0]), .I1(\data_in[1] [5]), 
            .I2(\data_in[2] [4]), .I3(\data_in[1] [0]), .O(n17_adj_3676));
    defparam i7_4_lut_adj_891.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_892 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [19]), .I3(GND_net), .O(n25683));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_892.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_4_lut_adj_893 (.I0(n17_adj_3676), .I1(\data_in[0] [3]), .I2(n16_adj_3675), 
            .I3(\data_in[1] [4]), .O(n63_c));
    defparam i9_4_lut_adj_893.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_894 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [18]), .I3(GND_net), .O(n7_adj_3677));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_894.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_895 (.I0(n13402), .I1(\data_in[3] [6]), .I2(\data_in[0] [2]), 
            .I3(\data_in[0] [7]), .O(n18_adj_3678));
    defparam i7_4_lut_adj_895.LUT_INIT = 16'hffef;
    SB_CARRY add_43_11 (.CI(n21976), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n21977));
    SB_LUT4 add_43_10_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n21975), .O(n2_adj_3679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i23319_4_lut (.I0(\data_in[3] [3]), .I1(\data_in[2] [3]), .I2(\data_in[3] [1]), 
            .I3(\data_in[3] [5]), .O(n28382));
    defparam i23319_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_896 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [17]), .I3(GND_net), .O(n25681));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_896.LUT_INIT = 16'he0e0;
    SB_LUT4 i10_4_lut_adj_897 (.I0(n28382), .I1(\data_in[2] [1]), .I2(n18_adj_3678), 
            .I3(n12_adj_3680), .O(n63_adj_3681));
    defparam i10_4_lut_adj_897.LUT_INIT = 16'hfff7;
    SB_LUT4 i3_4_lut_adj_898 (.I0(\data_in[3] [7]), .I1(n97), .I2(\data_in[0] [5]), 
            .I3(n17879), .O(n82));   // verilog/coms.v(95[12:19])
    defparam i3_4_lut_adj_898.LUT_INIT = 16'hffef;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n22004), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n14614), .D(n8825[2]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14956_4_lut (.I0(n5_adj_3682), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i14956_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_3_lut_adj_899 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [16]), .I3(GND_net), .O(n18717));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_899.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_900 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [15]), .I3(GND_net), .O(n7_adj_3683));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_900.LUT_INIT = 16'he0e0;
    SB_LUT4 i14924_2_lut_3_lut (.I0(n2_adj_3663), .I1(n2_adj_3664), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n18713));   // verilog/coms.v(115[11:12])
    defparam i14924_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i15099_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n8604), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2380 [0]));
    defparam i15099_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut_adj_901 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [13]), .I3(GND_net), .O(n7_adj_3684));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_901.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_902 (.I0(\FRAME_MATCHER.state [1]), .I1(n88), .I2(n17125), 
            .I3(\FRAME_MATCHER.state [3]), .O(n63));   // verilog/coms.v(201[5:24])
    defparam i3_4_lut_adj_902.LUT_INIT = 16'hfeff;
    SB_LUT4 i12_4_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [21]), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_903 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [29]), .O(n26_adj_3686));
    defparam i10_4_lut_adj_903.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i [23]), 
            .I2(\FRAME_MATCHER.i [17]), .I3(\FRAME_MATCHER.i [25]), .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_904 (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [6]), .O(n25));
    defparam i9_4_lut_adj_904.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_905 (.I0(n25), .I1(n27), .I2(n26_adj_3686), 
            .I3(n28), .O(n28207));
    defparam i15_4_lut_adj_905.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_906 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [7]), .O(n18_adj_3687));
    defparam i7_4_lut_adj_906.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_907 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [12]), .I3(GND_net), .O(n25679));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_907.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_2_lut_adj_908 (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3688));
    defparam i5_2_lut_adj_908.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_909 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [11]), .I3(GND_net), .O(n7_adj_3689));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_909.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_4_lut_adj_910 (.I0(\FRAME_MATCHER.i [14]), .I1(n18_adj_3687), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n28207), .O(n20_adj_3690));
    defparam i9_4_lut_adj_910.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_911 (.I0(\FRAME_MATCHER.i [9]), .I1(n20_adj_3690), 
            .I2(n16_adj_3688), .I3(\FRAME_MATCHER.i [27]), .O(n13538));
    defparam i10_4_lut_adj_911.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_912 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [10]), .I3(GND_net), .O(n25677));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_912.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\FRAME_MATCHER.i [4]), .I1(n13538), .I2(GND_net), 
            .I3(GND_net), .O(n13372));
    defparam i1_2_lut_adj_913.LUT_INIT = 16'heeee;
    SB_CARRY add_43_10 (.CI(n21975), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n21976));
    SB_LUT4 i11364_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n15169));
    defparam i11364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14946_4_lut (.I0(n8_adj_3691), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n13372), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i14946_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_3_lut_adj_914 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [9]), .I3(GND_net), .O(n25675));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_914.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_915 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [8]), .I3(GND_net), .O(n25673));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_915.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_9_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n21974), .O(n2_adj_3692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3971_8 (.CI(n22004), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n22005));
    SB_LUT4 i1_2_lut_3_lut_adj_916 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [7]), .I3(GND_net), .O(n7_adj_3693));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_916.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_9 (.CI(n21974), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n21975));
    SB_LUT4 i11365_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n15170));
    defparam i11365_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut (.I0(n63), .I1(\FRAME_MATCHER.state_31__N_2380 [0]), 
            .I2(n3), .I3(n4_adj_3695), .O(n25725));
    defparam i1_4_lut.LUT_INIT = 16'hddd5;
    SB_LUT4 i1_2_lut_3_lut_adj_917 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [6]), .I3(GND_net), .O(n25663));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_917.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_918 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [5]), .I3(GND_net), .O(n7_adj_3696));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_918.LUT_INIT = 16'he0e0;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n14614), .D(n8825[1]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11366_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n15171));
    defparam i11366_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_919 (.I0(n2_adj_3663), .I1(n2_adj_3664), 
            .I2(\FRAME_MATCHER.state [4]), .I3(GND_net), .O(n25669));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_adj_919.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_920 (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [30]), .O(n25481));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_920.LUT_INIT = 16'hfe00;
    SB_LUT4 i11351_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n15156));
    defparam i11351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n22003), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11352_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n15157));
    defparam i11352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_921 (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [26]), .O(n19229));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_921.LUT_INIT = 16'hfe00;
    SB_LUT4 i11353_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n15158));
    defparam i11353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_922 (.I0(n26486), .I1(n26154), .I2(\data_in_frame[6] [6]), 
            .I3(n6_adj_3662), .O(n13826));   // verilog/coms.v(166[9:87])
    defparam i4_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n130));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_924 (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_3698));
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h8888;
    SB_LUT4 i18117_2_lut_4_lut (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [25]), .O(n23168));   // verilog/coms.v(115[11:12])
    defparam i18117_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i2_4_lut_adj_925 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[4]), .I3(n2_adj_3698), .O(n27344));
    defparam i2_4_lut_adj_925.LUT_INIT = 16'ha080;
    SB_LUT4 i25158_4_lut (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[7]), .I3(n27344), .O(tx_transmit_N_3233));
    defparam i25158_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n88));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_927 (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [24]), .O(n19227));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_927.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_4_lut_adj_928 (.I0(\FRAME_MATCHER.state [1]), .I1(n26051), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n88), .O(n26052));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_928.LUT_INIT = 16'hfcec;
    SB_LUT4 i41_4_lut (.I0(n13), .I1(n29270), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n2786[0]));   // verilog/coms.v(102[12:33])
    defparam i41_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i11354_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n15159));
    defparam i11354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15426_2_lut_4_lut (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [16]), .O(n19225));   // verilog/coms.v(115[11:12])
    defparam i15426_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_CARRY add_3971_7 (.CI(n22003), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n22004));
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n22002), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i134_2_lut_4_lut (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [7]), .O(n8_adj_3699));   // verilog/coms.v(115[11:12])
    defparam i134_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i11355_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n15160));
    defparam i11355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11356_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n15161));
    defparam i11356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i139_2_lut_4_lut (.I0(n101), .I1(n3_adj_3661), .I2(n112), 
            .I3(\FRAME_MATCHER.state [5]), .O(n8_adj_3700));   // verilog/coms.v(115[11:12])
    defparam i139_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i18119_2_lut_4_lut (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [22]), .O(n23172));   // verilog/coms.v(95[12:19])
    defparam i18119_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_929 (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [20]), .O(n8_adj_3701));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_4_lut_adj_929.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_930 (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [18]), .O(n8_adj_3702));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_4_lut_adj_930.LUT_INIT = 16'hfe00;
    SB_CARRY add_3971_6 (.CI(n22002), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n22003));
    SB_LUT4 add_43_8_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n21973), .O(n2_adj_3703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_931 (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [15]), .O(n8_adj_3704));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_4_lut_adj_931.LUT_INIT = 16'hfe00;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n22001), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_8 (.CI(n21973), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n21974));
    SB_LUT4 i15425_2_lut_4_lut (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [14]), .O(n19223));   // verilog/coms.v(95[12:19])
    defparam i15425_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_CARRY add_3971_5 (.CI(n22001), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n22002));
    SB_LUT4 i1_2_lut_4_lut_adj_932 (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [13]), .O(n25459));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_4_lut_adj_932.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_933 (.I0(n112), .I1(n101), .I2(n3_adj_3661), 
            .I3(\FRAME_MATCHER.state [11]), .O(n8_adj_3705));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_4_lut_adj_933.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_934 (.I0(n26334), .I1(n26544), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[16] [6]), .O(n26380));
    defparam i1_2_lut_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_935 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3706));
    defparam i5_4_lut_adj_935.LUT_INIT = 16'h0200;
    SB_LUT4 i11357_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n15162));
    defparam i11357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_936 (.I0(n26334), .I1(n26544), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[16] [5]), .O(n26362));
    defparam i1_2_lut_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_937 (.I0(n18732), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n26044));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_937.LUT_INIT = 16'hffdf;
    SB_LUT4 i17_3_lut_4_lut (.I0(n14289), .I1(n26500), .I2(n34), .I3(\data_in_frame[9] [6]), 
            .O(n39));   // verilog/coms.v(73[16:42])
    defparam i17_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_7_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n21972), .O(n2_adj_3707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n21972), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n21973));
    SB_LUT4 i11358_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n15163));
    defparam i11358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11343_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n15148));
    defparam i11343_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_938 (.I0(\FRAME_MATCHER.state [1]), .I1(n83), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n13503));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_938.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_939 (.I0(n14289), .I1(n26500), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n13604));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_939.LUT_INIT = 16'h9696;
    SB_LUT4 i11344_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n15149));
    defparam i11344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_940 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n26278), .I3(\data_in_frame[6] [7]), .O(Kp_23__N_650));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_940.LUT_INIT = 16'h6996;
    SB_LUT4 i11345_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n15150));
    defparam i11345_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_6_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n21971), .O(n2_adj_3709)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n22000), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11346_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n15151));
    defparam i11346_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_941 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[8] [7]), .I3(n14111), .O(n26209));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_942 (.I0(\data_in_frame[6] [5]), .I1(n14224), .I2(n26145), 
            .I3(n6_adj_3710), .O(Kp_23__N_915));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_943 (.I0(\data_in_frame[6] [2]), .I1(n26482), 
            .I2(\data_in_frame[8] [3]), .I3(n26244), .O(n6_adj_3711));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i11347_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n15152));
    defparam i11347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_944 (.I0(\data_in_frame[6] [2]), .I1(n26482), 
            .I2(\data_in_frame[8] [3]), .I3(\data_in_frame[3] [7]), .O(n6_adj_3712));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_945 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[6] [4]), .O(n26278));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i11348_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n15153));
    defparam i11348_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_946 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[8] [4]), .I3(n14273), .O(n14294));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i11349_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n15154));
    defparam i11349_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_947 (.I0(n12779), .I1(\data_in_frame[2] [7]), 
            .I2(n10_adj_3713), .I3(Kp_23__N_708), .O(n23701));
    defparam i5_3_lut_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_948 (.I0(n12779), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[5] [3]), .I3(GND_net), .O(n26457));
    defparam i1_2_lut_3_lut_adj_948.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_4 (.CI(n22000), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n22001));
    SB_LUT4 i2_3_lut_4_lut_adj_949 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[3] [0]), .I3(Kp_23__N_708), .O(n14403));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_950 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [2]), .O(n26106));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i23288_2_lut (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28350));
    defparam i23288_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_43_6 (.CI(n21971), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n21972));
    SB_LUT4 add_43_5_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n21970), .O(n2_adj_3714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[0] [5]), .I2(\data_in[2] [4]), 
            .I3(GND_net), .O(n8_adj_3715));
    defparam i3_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i11350_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n15155));
    defparam i11350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n17879), .I1(n92[1]), .I2(n8_adj_3715), 
            .I3(\data_in[3] [7]), .O(\FRAME_MATCHER.state_31__N_2380 [1]));   // verilog/coms.v(95[12:19])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'hccdc;
    SB_LUT4 i11335_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n15140));
    defparam i11335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26559));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_953 (.I0(n26581), .I1(n26343), .I2(\data_in_frame[10] [7]), 
            .I3(n26649), .O(n10_adj_3717));
    defparam i4_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_954 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[10] [6]), 
            .I2(n26559), .I3(Kp_23__N_915), .O(n14_adj_3718));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\data_in_frame[15] [4]), .I1(n26636), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3719));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_956 (.I0(n9_adj_3719), .I1(n14_adj_3718), .I2(n24641), 
            .I3(n14294), .O(n23804));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_956.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26405));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_958 (.I0(n82), .I1(\FRAME_MATCHER.state [2]), .I2(n63_c), 
            .I3(n63_adj_3681), .O(\FRAME_MATCHER.state_31__N_2380[2] ));   // verilog/coms.v(95[12:19])
    defparam i1_4_lut_adj_958.LUT_INIT = 16'h8a0a;
    SB_LUT4 equal_1120_i7_2_lut (.I0(Kp_23__N_915), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3720));   // verilog/coms.v(236[9:81])
    defparam equal_1120_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11336_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n15141));
    defparam i11336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_959 (.I0(\FRAME_MATCHER.state [1]), .I1(n17197), 
            .I2(n17173), .I3(GND_net), .O(n1656));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut_3_lut_adj_959.LUT_INIT = 16'hf4f4;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n21999), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(n26571), .I3(n26214), .O(n6_adj_3721));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_960 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(Kp_23__N_1026), .I3(n26214), .O(n26526));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_961 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(n26343), .I3(GND_net), .O(n26547));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_961.LUT_INIT = 16'h9696;
    SB_LUT4 i11337_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n15142));
    defparam i11337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_962 (.I0(n13826), .I1(n26500), .I2(\data_in_frame[9] [2]), 
            .I3(GND_net), .O(n26445));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_962.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_963 (.I0(n23804), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26645));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_964 (.I0(\data_in_frame[11] [4]), .I1(n13604), 
            .I2(GND_net), .I3(GND_net), .O(n14149));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(n14429), .I1(n23657), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_3722));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_965 (.I0(\data_in_frame[16] [3]), .I1(n14149), 
            .I2(n26445), .I3(\data_in_frame[14] [0]), .O(n14_adj_3723));
    defparam i6_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_966 (.I0(\data_in_frame[18] [4]), .I1(n14_adj_3723), 
            .I2(n10_adj_3722), .I3(n26596), .O(n26136));
    defparam i7_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_3 (.CI(n21999), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n22000));
    SB_LUT4 i2_3_lut_4_lut_adj_967 (.I0(n24179), .I1(n27569), .I2(\data_in_frame[9] [5]), 
            .I3(n23779), .O(n26649));
    defparam i2_3_lut_4_lut_adj_967.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26203));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_969 (.I0(n26214), .I1(\data_in_frame[11] [6]), 
            .I2(n26190), .I3(n24616), .O(n28_adj_3724));
    defparam i12_4_lut_adj_969.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_970 (.I0(\data_in_frame[6] [5]), .I1(n26259), 
            .I2(n26655), .I3(\data_in_frame[5] [0]), .O(n26_adj_3725));
    defparam i10_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_971 (.I0(n23828), .I1(n26609), .I2(n26689), 
            .I3(n26278), .O(n27_adj_3726));
    defparam i11_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_972 (.I0(\data_in_frame[14] [2]), .I1(n26203), 
            .I2(n26699), .I3(n26486), .O(n25_adj_3727));
    defparam i9_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_973 (.I0(n25_adj_3727), .I1(n27_adj_3726), .I2(n26_adj_3725), 
            .I3(n28_adj_3724), .O(n23657));
    defparam i15_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_974 (.I0(n23657), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26565));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_975 (.I0(n26380), .I1(n27426), .I2(\data_in_frame[19] [0]), 
            .I3(n26565), .O(n10_adj_3728));
    defparam i4_4_lut_adj_975.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_976 (.I0(\data_in_frame[18] [7]), .I1(n10_adj_3728), 
            .I2(n23841), .I3(GND_net), .O(n24618));
    defparam i5_3_lut_adj_976.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_15__7__I_0_3897_2_lut (.I0(\data_in_frame[15] [7]), 
            .I1(\data_in_frame[15] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1237));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_15__7__I_0_3897_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_977 (.I0(\data_in_frame[13] [6]), .I1(n26547), 
            .I2(\data_in_frame[11] [5]), .I3(\data_in_frame[11] [4]), .O(n24653));
    defparam i3_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[16] [0]), .I1(n24653), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n6_adj_3729));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_978 (.I0(Kp_23__N_1237), .I1(n24728), .I2(n26409), 
            .I3(n6_adj_3729), .O(n26337));
    defparam i4_4_lut_adj_978.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_979 (.I0(n24735), .I1(n24639), .I2(\data_in_frame[17] [1]), 
            .I3(GND_net), .O(n26421));
    defparam i2_3_lut_adj_979.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_980 (.I0(n13253), .I1(n26421), .I2(\data_in_frame[19] [3]), 
            .I3(\data_in_frame[19] [2]), .O(n26206));
    defparam i2_4_lut_adj_980.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_981 (.I0(n14315), .I1(\data_in_frame[19] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n26275));
    defparam i1_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_982 (.I0(n24179), .I1(n27569), .I2(\data_in_frame[12] [1]), 
            .I3(GND_net), .O(n26571));
    defparam i1_2_lut_3_lut_adj_982.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_983 (.I0(n26337), .I1(n26262), .I2(\data_in_frame[19] [7]), 
            .I3(n26395), .O(n10_adj_3730));
    defparam i4_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_984 (.I0(n26275), .I1(n10_adj_3730), .I2(n26206), 
            .I3(GND_net), .O(n24052));
    defparam i5_3_lut_adj_984.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_in_frame[9] [0]), .I1(n13670), .I2(GND_net), 
            .I3(GND_net), .O(n14309));
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_986 (.I0(\data_in_frame[9] [7]), .I1(n23701), .I2(\data_in_frame[11] [7]), 
            .I3(n6_adj_3721), .O(n26655));
    defparam i4_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_987 (.I0(\data_in_frame[12] [2]), .I1(n26655), 
            .I2(n14309), .I3(n24637), .O(n23621));
    defparam i3_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26418));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_989 (.I0(Kp_23__N_1026), .I1(n13882), .I2(n13890), 
            .I3(GND_net), .O(n23477));
    defparam i2_3_lut_adj_989.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_990 (.I0(n26529), .I1(Kp_23__N_915), .I2(\data_in_frame[8] [4]), 
            .I3(n26389), .O(n15_adj_3731));
    defparam i6_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_adj_3731), .I1(\data_in_frame[8] [2]), .I2(n14_adj_3732), 
            .I3(n23477), .O(n24616));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_991 (.I0(n27569), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[9] [6]), .I3(\data_in_frame[11] [7]), .O(n26689));
    defparam i2_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_992 (.I0(\data_in_frame[4] [1]), .I1(n24616), .I2(n14098), 
            .I3(n6_adj_3733), .O(n26340));
    defparam i4_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_993 (.I0(n23841), .I1(n26340), .I2(\data_in_frame[9] [1]), 
            .I3(n24599), .O(n10_adj_3734));
    defparam i4_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_994 (.I0(\data_in_frame[11] [5]), .I1(n4_adj_3735), 
            .I2(n10_adj_3734), .I3(\data_in_frame[13] [7]), .O(n26132));
    defparam i2_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26214));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i11328_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n15133));
    defparam i11328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_996 (.I0(n13826), .I1(n26190), .I2(GND_net), 
            .I3(GND_net), .O(n14503));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_997 (.I0(Kp_23__N_915), .I1(n13670), .I2(GND_net), 
            .I3(GND_net), .O(n26415));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_998 (.I0(n24179), .I1(n26526), .I2(n26259), .I3(n23681), 
            .O(n27569));
    defparam i3_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_CARRY add_43_5 (.CI(n21970), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n21971));
    SB_LUT4 i11329_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n15134));
    defparam i11329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11330_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n15135));
    defparam i11330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11331_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n15136));
    defparam i11331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_999 (.I0(n14111), .I1(Kp_23__N_656), .I2(n14273), 
            .I3(n26389), .O(n10_adj_3736));
    defparam i4_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i11332_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n15137));
    defparam i11332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11333_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n15138));
    defparam i11333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11334_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n15139));
    defparam i11334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1000 (.I0(n4_adj_3737), .I1(Kp_23__N_816), .I2(n10_adj_3736), 
            .I3(Kp_23__N_650), .O(n20_adj_3738));
    defparam i4_4_lut_adj_1000.LUT_INIT = 16'hebbe;
    SB_LUT4 i12_4_lut_adj_1001 (.I0(n23681), .I1(n7_adj_3720), .I2(n14294), 
            .I3(n13890), .O(n28_adj_3739));
    defparam i12_4_lut_adj_1001.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_4_lut_adj_1002 (.I0(n12779), .I1(n26184), .I2(\data_in_frame[7] [2]), 
            .I3(\data_in_frame[5] [1]), .O(n12_adj_3740));
    defparam i5_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1003 (.I0(n24659), .I1(n20_adj_3738), .I2(n26209), 
            .I3(\data_in_frame[7] [7]), .O(n26_adj_3741));
    defparam i10_4_lut_adj_1003.LUT_INIT = 16'hfefd;
    SB_LUT4 i6_4_lut_adj_1004 (.I0(n13685), .I1(n12_adj_3740), .I2(n26196), 
            .I3(n14403), .O(n14289));
    defparam i6_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1005 (.I0(n26500), .I1(n14140), .I2(n23701), 
            .I3(n13670), .O(n27_adj_3742));
    defparam i11_4_lut_adj_1005.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(n26180), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13882));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[8] [0]), .I1(n24006), 
            .I2(GND_net), .I3(GND_net), .O(n24719));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1008 (.I0(n24719), .I1(n13882), .I2(n14289), 
            .I3(n13826), .O(n25_adj_3743));
    defparam i9_4_lut_adj_1008.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut_adj_1009 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[6] [7]), .I3(GND_net), .O(n26699));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1009.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_1010 (.I0(n25_adj_3743), .I1(n27_adj_3742), .I2(n26_adj_3741), 
            .I3(n28_adj_3739), .O(n31));
    defparam i15_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1011 (.I0(\FRAME_MATCHER.state [1]), .I1(n31), 
            .I2(n11166), .I3(GND_net), .O(n3938));
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26492));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\FRAME_MATCHER.state [26]), .I1(\FRAME_MATCHER.state [20]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3744));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1014 (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(\FRAME_MATCHER.state [24]), .I3(n6_adj_3744), .O(n26033));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1014.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26154));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1016 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [17]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [23]), 
            .O(n18_adj_3745));
    defparam i7_4_lut_adj_1016.LUT_INIT = 16'hfffe;
    SB_LUT4 i11026_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n14831));
    defparam i11026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1017 (.I0(n27637), .I1(\data_out_frame[20] [2]), 
            .I2(n24635), .I3(GND_net), .O(n26556));
    defparam i1_2_lut_3_lut_adj_1017.LUT_INIT = 16'h9696;
    SB_LUT4 i5_2_lut_adj_1018 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3746));
    defparam i5_2_lut_adj_1018.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1019 (.I0(\FRAME_MATCHER.state [27]), .I1(n18_adj_3745), 
            .I2(\FRAME_MATCHER.state [22]), .I3(\FRAME_MATCHER.state [25]), 
            .O(n20_adj_3747));
    defparam i9_4_lut_adj_1019.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1020 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n18732), .O(n26057));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1020.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut_adj_1021 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n18732), .O(n26035));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1021.LUT_INIT = 16'hfeff;
    SB_LUT4 i10_4_lut_adj_1022 (.I0(\FRAME_MATCHER.state [28]), .I1(n20_adj_3747), 
            .I2(n16_adj_3746), .I3(\FRAME_MATCHER.state [19]), .O(n26079));
    defparam i10_4_lut_adj_1022.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1023 (.I0(n26529), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[1] [5]), .I3(n6_adj_3748), .O(n13670));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1024 (.I0(\data_in_frame[7] [3]), .I1(n26129), 
            .I2(\data_in_frame[0] [7]), .I3(n14432), .O(n10_adj_3713));   // verilog/coms.v(71[16:69])
    defparam i4_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1025 (.I0(\FRAME_MATCHER.state [7]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [5]), .I3(\FRAME_MATCHER.state [4]), 
            .O(n18866));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1026 (.I0(\FRAME_MATCHER.state [9]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(\FRAME_MATCHER.state [15]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n10_adj_3749));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1027 (.I0(\data_in_frame[6] [0]), .I1(Kp_23__N_656), 
            .I2(\data_in_frame[6] [1]), .I3(n26233), .O(n10_adj_3750));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [14]), 
            .I2(GND_net), .I3(GND_net), .O(n21564));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(\FRAME_MATCHER.state [11]), .I1(n21564), 
            .I2(n10_adj_3749), .I3(\FRAME_MATCHER.state [8]), .O(n6_adj_3751));   // verilog/coms.v(201[5:24])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(n26196), .I1(n26699), .I2(n14524), 
            .I3(GND_net), .O(n26500));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1031 (.I0(\FRAME_MATCHER.state [1]), .I1(n17197), 
            .I2(n3303), .I3(n2_adj_3752), .O(n4_adj_3695));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1031.LUT_INIT = 16'hff04;
    SB_LUT4 i7_4_lut_adj_1032 (.I0(\data_in_frame[0] [2]), .I1(n14_adj_3753), 
            .I2(n28350), .I3(\data_in_frame[0] [4]), .O(n11166));
    defparam i7_4_lut_adj_1032.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_1033 (.I0(n14524), .I1(\data_in_frame[6] [0]), 
            .I2(Kp_23__N_650), .I3(GND_net), .O(n14098));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1034 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n11166), .I3(n26051), .O(n10_adj_3754));
    defparam i4_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1035 (.I0(\data_in_frame[5] [5]), .I1(n13915), 
            .I2(n26250), .I3(n13804), .O(n26272));
    defparam i3_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i25084_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n10_adj_3754), 
            .I2(n10649), .I3(GND_net), .O(n14593));
    defparam i25084_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i3_2_lut_4_lut_4_lut (.I0(n23661), .I1(n16570), .I2(n24622), 
            .I3(n26303), .O(n11));
    defparam i3_2_lut_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1036 (.I0(n13685), .I1(n14196), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n14524));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_LUT4 i11338_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n15143));
    defparam i11338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1037 (.I0(n13685), .I1(n14196), .I2(n14192), 
            .I3(GND_net), .O(n6_adj_3656));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1037.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1038 (.I0(n13503), .I1(n25968), .I2(n31_adj_3653), 
            .I3(GND_net), .O(n4137));
    defparam i2_3_lut_adj_1038.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut_adj_1039 (.I0(n26079), .I1(n26033), .I2(n6_adj_3751), 
            .I3(n18866), .O(n9_adj_3755));
    defparam i2_3_lut_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1040 (.I0(n26079), .I1(n26033), .I2(n18866), 
            .I3(n6_adj_3751), .O(n26051));
    defparam i2_3_lut_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1041 (.I0(n26415), .I1(n26581), .I2(n24006), 
            .I3(n14503), .O(n12_adj_3756));
    defparam i5_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_4_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n21969), .O(n2_adj_3757)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_3_lut_adj_1042 (.I0(n26170), .I1(n26492), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n10_adj_3758));
    defparam i2_2_lut_3_lut_adj_1042.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1043 (.I0(Kp_23__N_1002), .I1(n12_adj_3756), .I2(n26630), 
            .I3(n14294), .O(n24179));
    defparam i6_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(n23681), .I1(n13890), .I2(GND_net), 
            .I3(GND_net), .O(n23779));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(n23701), .I1(n13890), .I2(GND_net), 
            .I3(GND_net), .O(n23794));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1026));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(n23701), .I1(n14289), .I2(GND_net), 
            .I3(GND_net), .O(n24599));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_in_frame[8] [6]), .I1(n26209), 
            .I2(GND_net), .I3(GND_net), .O(n13867));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1048 (.I0(Kp_23__N_915), .I1(n13867), .I2(\data_in_frame[9] [0]), 
            .I3(\data_in_frame[11] [2]), .O(n26089));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26140));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1050 (.I0(n26140), .I1(n26547), .I2(n13604), 
            .I3(n26089), .O(n12_adj_3759));
    defparam i5_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1051 (.I0(Kp_23__N_1026), .I1(n12_adj_3759), .I2(n26649), 
            .I3(n23794), .O(n24641));
    defparam i6_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1052 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[13] [3]), 
            .I2(n26409), .I3(n24641), .O(n23664));
    defparam i1_4_lut_adj_1052.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1053 (.I0(n26170), .I1(n26492), .I2(n10_adj_3750), 
            .I3(\data_in_frame[3] [6]), .O(n14140));
    defparam i5_3_lut_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26587));
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1256));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1055 (.I0(\data_in_frame[9] [4]), .I1(n26596), 
            .I2(n13604), .I3(GND_net), .O(n26671));
    defparam i2_3_lut_adj_1055.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1056 (.I0(Kp_23__N_1256), .I1(n26089), .I2(n26575), 
            .I3(n14429), .O(n14_adj_3760));   // verilog/coms.v(72[16:41])
    defparam i6_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1057 (.I0(\data_in_frame[18] [2]), .I1(n14_adj_3760), 
            .I2(n10_adj_3761), .I3(n26658), .O(n26624));   // verilog/coms.v(72[16:41])
    defparam i7_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1058 (.I0(\data_in_frame[16] [1]), .I1(n26340), 
            .I2(n26590), .I3(\data_in_frame[15] [7]), .O(n14_adj_3762));
    defparam i6_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1059 (.I0(\data_in_frame[18] [3]), .I1(n14_adj_3762), 
            .I2(n10_adj_3763), .I3(n26671), .O(n26476));
    defparam i7_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\data_in_frame[16] [0]), .I1(n23664), 
            .I2(GND_net), .I3(GND_net), .O(n23708));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1061 (.I0(n26132), .I1(n26362), .I2(n26136), 
            .I3(GND_net), .O(n42));
    defparam i5_3_lut_adj_1061.LUT_INIT = 16'h9696;
    SB_LUT4 i20_4_lut (.I0(n26308), .I1(n26421), .I2(n23664), .I3(n24689), 
            .O(n57));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1062 (.I0(\data_in_frame[14] [2]), .I1(n26571), 
            .I2(n23779), .I3(\data_in_frame[10] [3]), .O(n34));
    defparam i12_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[10] [1]), .I3(\data_in_frame[11] [4]), .O(n36));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n26328), .I1(n36), .I2(n26_adj_3764), .I3(\data_in_frame[10] [5]), 
            .O(n40));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\data_in_frame[9] [1]), .I1(n13882), .I2(\data_in_frame[10] [6]), 
            .I3(\data_in_frame[11] [3]), .O(n38));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(n28350), .I3(n13_adj_3706), .O(n25968));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3753));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i11339_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n15144));
    defparam i11339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1063 (.I0(n26652), .I1(n26334), .I2(n26423), 
            .I3(n26140), .O(n37));
    defparam i15_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n27143));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n57), .I1(\data_in_frame[18] [1]), .I2(n42), 
            .I3(n26645), .O(n66));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[11] [5]), 
            .I2(\data_in_frame[14] [4]), .I3(Kp_23__N_1237), .O(n64));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n24599), .I1(\data_in_frame[15] [0]), .I2(\data_in_frame[15] [4]), 
            .I3(n38_adj_3765), .O(n65));
    defparam i28_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n26658), .I1(n26418), .I2(n26520), .I3(\data_in_frame[16] [6]), 
            .O(n63_adj_3766));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(\data_in_frame[16] [5]), .I1(n26587), .I2(n27143), 
            .I3(\data_in_frame[13] [5]), .O(n60));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(n26476), .I1(\data_in_frame[16] [4]), .I2(n26624), 
            .I3(GND_net), .O(n43));
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[15] [2]), 
            .I2(n14485), .I3(n23708), .O(n62));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(\data_in_frame[15] [5]), .I1(n26517), .I2(n26671), 
            .I3(\data_in_frame[13] [3]), .O(n61));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(n63_adj_3766), .I1(n65), .I2(n64), .I3(n66), 
            .O(n72));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n43), .I1(n60), .I2(\data_in_frame[17] [7]), 
            .I3(n24414), .O(n67));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i36_4_lut (.I0(n67), .I1(n72), .I2(n61), .I3(n62), .O(n24728));
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1064 (.I0(n26203), .I1(n26233), .I2(n26492), 
            .I3(n6_adj_3711), .O(Kp_23__N_1002));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1065 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[12] [4]), .O(n26328));
    defparam i3_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1066 (.I0(n24719), .I1(n26630), .I2(n24659), 
            .I3(\data_in_frame[7] [7]), .O(n24206));
    defparam i3_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1067 (.I0(n26353), .I1(\data_in_frame[8] [0]), 
            .I2(n13719), .I3(n23681), .O(n14_adj_3767));
    defparam i6_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1068 (.I0(\data_in_frame[10] [1]), .I1(n14_adj_3767), 
            .I2(n10_adj_3758), .I3(n13813), .O(n24637));
    defparam i7_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1069 (.I0(\data_in_frame[12] [3]), .I1(n24637), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n26292));
    defparam i2_3_lut_adj_1069.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1070 (.I0(n26292), .I1(\data_in_frame[14] [5]), 
            .I2(n13904), .I3(GND_net), .O(n27426));
    defparam i2_3_lut_adj_1070.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1071 (.I0(\data_in_frame[14] [3]), .I1(n23621), 
            .I2(n26553), .I3(GND_net), .O(n8_adj_3768));
    defparam i3_3_lut_adj_1071.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(\data_in_frame[18] [7]), .I1(n27426), 
            .I2(n8_adj_3768), .I3(n26362), .O(n24689));
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 i126_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n17197), 
            .I2(n3303), .I3(n8604), .O(n112));   // verilog/coms.v(127[12] 300[6])
    defparam i126_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i4_4_lut_adj_1073 (.I0(\data_in_frame[14] [7]), .I1(n26292), 
            .I2(n26436), .I3(n6_adj_3769), .O(n24639));
    defparam i4_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1074 (.I0(\data_in_frame[14] [6]), .I1(n24206), 
            .I2(n26328), .I3(Kp_23__N_1002), .O(n27074));
    defparam i3_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1075 (.I0(\data_in_frame[17] [0]), .I1(n27074), 
            .I2(\data_in_frame[16] [7]), .I3(GND_net), .O(n26553));
    defparam i2_3_lut_adj_1075.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1076 (.I0(\data_in_frame[17] [1]), .I1(n26553), 
            .I2(n26380), .I3(n24639), .O(n13253));
    defparam i3_4_lut_adj_1076.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\data_in_frame[19] [1]), .I1(n24689), 
            .I2(GND_net), .I3(GND_net), .O(n26262));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1078 (.I0(\data_in_frame[7] [7]), .I1(n26272), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n13719));
    defparam i2_3_lut_adj_1078.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1079 (.I0(\data_in_frame[8] [1]), .I1(n26227), 
            .I2(\data_in_frame[6] [0]), .I3(n13719), .O(n13921));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1080 (.I0(n13921), .I1(n14140), .I2(\data_in_frame[10] [3]), 
            .I3(GND_net), .O(n13904));
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26517));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1082 (.I0(n26436), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3770));
    defparam i2_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1083 (.I0(n26544), .I1(\data_in_frame[12] [4]), 
            .I2(n26086), .I3(\data_in_frame[15] [1]), .O(n14_adj_3771));
    defparam i6_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1084 (.I0(\data_in_frame[17] [2]), .I1(n14_adj_3771), 
            .I2(n10_adj_3770), .I3(\data_in_frame[14] [6]), .O(n24735));
    defparam i7_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1085 (.I0(n26247), .I1(n26520), .I2(\data_in_frame[17] [4]), 
            .I3(n4_adj_3737), .O(n12_adj_3772));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1086 (.I0(\data_in_frame[11] [3]), .I1(n26445), 
            .I2(n26089), .I3(GND_net), .O(Kp_23__N_1283));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1086.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1087 (.I0(\data_in_frame[11] [3]), .I1(n26445), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n10_adj_3763));   // verilog/coms.v(73[16:42])
    defparam i2_2_lut_3_lut_adj_1087.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1088 (.I0(n14140), .I1(n12_adj_3772), .I2(n26636), 
            .I3(\data_in_frame[10] [4]), .O(n14152));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1089 (.I0(\data_in_frame[13] [1]), .I1(n26247), 
            .I2(\data_in_frame[17] [3]), .I3(\data_in_frame[10] [7]), .O(n12_adj_3773));
    defparam i5_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1090 (.I0(\data_in_frame[12] [5]), .I1(n12_adj_3773), 
            .I2(n26517), .I3(n13904), .O(n14315));
    defparam i6_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(n14315), .I1(n14152), .I2(GND_net), 
            .I3(GND_net), .O(n26308));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1092 (.I0(\data_in_frame[19] [4]), .I1(n24735), 
            .I2(n14315), .I3(GND_net), .O(n26395));
    defparam i1_3_lut_adj_1092.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n14485));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(n26337), .I1(\data_in_frame[19] [7]), 
            .I2(n24414), .I3(GND_net), .O(n26541));
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1095 (.I0(n26433), .I1(\data_in_frame[15] [3]), 
            .I2(n12002), .I3(n23804), .O(n14_adj_3774));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1096 (.I0(\data_in_frame[17] [5]), .I1(n14_adj_3774), 
            .I2(n10_adj_3775), .I3(n14485), .O(n24414));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1097 (.I0(Kp_23__N_1283), .I1(n26661), .I2(n26645), 
            .I3(n26405), .O(n26693));
    defparam i3_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1098 (.I0(\data_in_frame[20] [2]), .I1(n26693), 
            .I2(n26538), .I3(\data_in_frame[18] [0]), .O(n27162));
    defparam i3_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1099 (.I0(\data_in_frame[20] [1]), .I1(n24653), 
            .I2(n26541), .I3(GND_net), .O(n8_adj_3776));
    defparam i3_3_lut_adj_1099.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_adj_1100 (.I0(\data_in_frame[20] [6]), .I1(n26132), 
            .I2(n26136), .I3(GND_net), .O(n26480));
    defparam i1_3_lut_adj_1100.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1101 (.I0(\data_in_frame[21] [5]), .I1(n26395), 
            .I2(n26421), .I3(\data_in_frame[19] [3]), .O(n28168));
    defparam i3_4_lut_adj_1101.LUT_INIT = 16'h9669;
    SB_LUT4 i23296_4_lut (.I0(n24728), .I1(n26480), .I2(n8_adj_3776), 
            .I3(n26331), .O(n28358));
    defparam i23296_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i3_4_lut_adj_1102 (.I0(\data_in_frame[20] [3]), .I1(n26624), 
            .I2(n26538), .I3(n26331), .O(n28018));
    defparam i3_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1103 (.I0(n24653), .I1(n14152), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n10_adj_3777));
    defparam i3_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(n26693), .I1(\data_in_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3778));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1105 (.I0(n24414), .I1(n10_adj_3777), .I2(\data_in_frame[19] [6]), 
            .I3(n26541), .O(n12_adj_3779));
    defparam i5_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1106 (.I0(\data_in_frame[19] [2]), .I1(n26262), 
            .I2(\data_in_frame[21] [3]), .I3(n13253), .O(n27630));
    defparam i3_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1107 (.I0(\data_in_frame[19] [5]), .I1(n26395), 
            .I2(n26308), .I3(\data_in_frame[21] [6]), .O(n26964));
    defparam i3_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i23292_4_lut (.I0(n24728), .I1(n27630), .I2(n12_adj_3779), 
            .I3(n8_adj_3778), .O(n28354));
    defparam i23292_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [0]), 
            .I2(n26689), .I3(GND_net), .O(n26_adj_3764));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n12_adj_3780));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1108 (.I0(n24414), .I1(n12_adj_3780), .I2(\data_in_frame[19] [1]), 
            .I3(n26541), .O(n14_adj_3781));
    defparam i6_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1109 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[19] [2]), .I3(GND_net), .O(n9_adj_3782));
    defparam i1_3_lut_adj_1109.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1110 (.I0(n9_adj_3782), .I1(n14_adj_3781), .I2(n26132), 
            .I3(\data_in_frame[19] [0]), .O(n27416));
    defparam i7_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(n23683), .I1(n14098), .I2(GND_net), 
            .I3(GND_net), .O(n23699));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30565));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30565_bdd_4_lut (.I0(n30565), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30568));
    defparam n30565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n29799), .I2(n29274), .I3(byte_transmit_counter[4]), .O(n30559));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30559_bdd_4_lut (.I0(n30559), .I1(n14_adj_3648), .I2(n7_adj_3647), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n30559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25446 (.I0(byte_transmit_counter[3]), 
            .I1(n30304), .I2(n29238), .I3(byte_transmit_counter[4]), .O(n30553));
    defparam byte_transmit_counter_3__bdd_4_lut_25446.LUT_INIT = 16'he4aa;
    SB_LUT4 n30553_bdd_4_lut (.I0(n30553), .I1(n14_adj_3645), .I2(n7_adj_3644), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n30553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25451 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30547));
    defparam byte_transmit_counter_0__bdd_4_lut_25451.LUT_INIT = 16'he4aa;
    SB_LUT4 n30547_bdd_4_lut (.I0(n30547), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30550));
    defparam n30547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25441 (.I0(byte_transmit_counter[3]), 
            .I1(n30310), .I2(n29231), .I3(byte_transmit_counter[4]), .O(n30541));
    defparam byte_transmit_counter_3__bdd_4_lut_25441.LUT_INIT = 16'he4aa;
    SB_LUT4 n30541_bdd_4_lut (.I0(n30541), .I1(n14_adj_3642), .I2(n7_adj_3641), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n30541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n13804));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25431 (.I0(byte_transmit_counter[3]), 
            .I1(n30316), .I2(n29228), .I3(byte_transmit_counter[4]), .O(n30535));
    defparam byte_transmit_counter_3__bdd_4_lut_25431.LUT_INIT = 16'he4aa;
    SB_LUT4 n30535_bdd_4_lut (.I0(n30535), .I1(n14_adj_3638), .I2(n7_adj_3637), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n30535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25426 (.I0(byte_transmit_counter[3]), 
            .I1(n30526), .I2(n29225), .I3(byte_transmit_counter[4]), .O(n30529));
    defparam byte_transmit_counter_3__bdd_4_lut_25426.LUT_INIT = 16'he4aa;
    SB_LUT4 n30529_bdd_4_lut (.I0(n30529), .I1(n14_adj_3635), .I2(n7_adj_3634), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n30529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1113 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_708), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n12779));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n29226), .I2(n29227), .I3(byte_transmit_counter[2]), .O(n30523));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30523_bdd_4_lut (.I0(n30523), .I1(n17_adj_3632), .I2(n16_adj_3631), 
            .I3(byte_transmit_counter[2]), .O(n30526));
    defparam n30523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'hbbbb;
    SB_LUT4 i25170_4_lut (.I0(n133), .I1(\FRAME_MATCHER.state [0]), .I2(n9_adj_3755), 
            .I3(\FRAME_MATCHER.state [2]), .O(n27310));
    defparam i25170_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i5_3_lut_4_lut_adj_1115 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [0]), 
            .I2(n13719), .I3(\data_in_frame[8] [3]), .O(n14_adj_3732));
    defparam i5_3_lut_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25421 (.I0(byte_transmit_counter[3]), 
            .I1(n30328), .I2(n29222), .I3(byte_transmit_counter[4]), .O(n30517));
    defparam byte_transmit_counter_3__bdd_4_lut_25421.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut_adj_1116 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n11166), .I3(n10649), .O(n27889));
    defparam i2_4_lut_adj_1116.LUT_INIT = 16'h4440;
    SB_LUT4 i1_4_lut_adj_1117 (.I0(n27889), .I1(n4_c), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state_31__N_2444 [3]), .O(n14_adj_3783));
    defparam i1_4_lut_adj_1117.LUT_INIT = 16'haaab;
    SB_LUT4 n30517_bdd_4_lut (.I0(n30517), .I1(n14_adj_3629), .I2(n7_adj_3628), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n30517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i25173_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n4_adj_3784), 
            .I2(n14_adj_3783), .I3(n13), .O(n26987));
    defparam i25173_4_lut.LUT_INIT = 16'h0313;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26170));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25411 (.I0(byte_transmit_counter[3]), 
            .I1(n30334), .I2(n29219), .I3(byte_transmit_counter[4]), .O(n30511));
    defparam byte_transmit_counter_3__bdd_4_lut_25411.LUT_INIT = 16'he4aa;
    SB_LUT4 n30511_bdd_4_lut (.I0(n30511), .I1(n14_adj_3625), .I2(n7_adj_3624), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n30511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25436 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30505));
    defparam byte_transmit_counter_0__bdd_4_lut_25436.LUT_INIT = 16'he4aa;
    SB_LUT4 n30505_bdd_4_lut (.I0(n30505), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30508));
    defparam n30505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25401 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30499));
    defparam byte_transmit_counter_0__bdd_4_lut_25401.LUT_INIT = 16'he4aa;
    SB_LUT4 n30499_bdd_4_lut (.I0(n30499), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30502));
    defparam n30499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(n14403), .I1(n26457), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3785));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25396 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30493));
    defparam byte_transmit_counter_0__bdd_4_lut_25396.LUT_INIT = 16'he4aa;
    SB_LUT4 n30493_bdd_4_lut (.I0(n30493), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30496));
    defparam n30493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1120 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[7] [4]), 
            .I2(n26106), .I3(n6_adj_3785), .O(n26609));
    defparam i4_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25391 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30487));
    defparam byte_transmit_counter_0__bdd_4_lut_25391.LUT_INIT = 16'he4aa;
    SB_LUT4 n30487_bdd_4_lut (.I0(n30487), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30490));
    defparam n30487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25386 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30475));
    defparam byte_transmit_counter_0__bdd_4_lut_25386.LUT_INIT = 16'he4aa;
    SB_LUT4 n30475_bdd_4_lut (.I0(n30475), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30478));
    defparam n30475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1121 (.I0(n26457), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[7] [5]), .I3(n26495), .O(n10_adj_3786));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25376 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30469));
    defparam byte_transmit_counter_0__bdd_4_lut_25376.LUT_INIT = 16'he4aa;
    SB_LUT4 n30469_bdd_4_lut (.I0(n30469), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30472));
    defparam n30469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1122 (.I0(\data_in_frame[3] [1]), .I1(n10_adj_3786), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n23681));   // verilog/coms.v(85[17:63])
    defparam i5_3_lut_adj_1122.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25371 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30463));
    defparam byte_transmit_counter_0__bdd_4_lut_25371.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[14] [3]), 
            .I2(n23621), .I3(GND_net), .O(n23841));
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'h9696;
    SB_LUT4 n30463_bdd_4_lut (.I0(n30463), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30466));
    defparam n30463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25366 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30451));
    defparam byte_transmit_counter_0__bdd_4_lut_25366.LUT_INIT = 16'he4aa;
    SB_LUT4 n30451_bdd_4_lut (.I0(n30451), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30454));
    defparam n30451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(\data_out_frame[19] [4]), .I1(n16570), 
            .I2(n24622), .I3(GND_net), .O(n24756));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25356 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30445));
    defparam byte_transmit_counter_0__bdd_4_lut_25356.LUT_INIT = 16'he4aa;
    SB_LUT4 n30445_bdd_4_lut (.I0(n30445), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30448));
    defparam n30445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1125 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(n13178), .I3(GND_net), .O(n4_adj_3787));
    defparam i1_2_lut_3_lut_adj_1125.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25351 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30439));
    defparam byte_transmit_counter_0__bdd_4_lut_25351.LUT_INIT = 16'he4aa;
    SB_LUT4 n30439_bdd_4_lut (.I0(n30439), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30442));
    defparam n30439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1126 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[5] [6]), .O(n14_adj_3788));   // verilog/coms.v(85[17:63])
    defparam i5_3_lut_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25346 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30433));
    defparam byte_transmit_counter_0__bdd_4_lut_25346.LUT_INIT = 16'he4aa;
    SB_LUT4 n30433_bdd_4_lut (.I0(n30433), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30436));
    defparam n30433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1127 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n26677));
    defparam i1_2_lut_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25341 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30427));
    defparam byte_transmit_counter_0__bdd_4_lut_25341.LUT_INIT = 16'he4aa;
    SB_LUT4 n30427_bdd_4_lut (.I0(n30427), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30430));
    defparam n30427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[14] [2]), .I3(GND_net), .O(n26454));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25336 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30421));
    defparam byte_transmit_counter_0__bdd_4_lut_25336.LUT_INIT = 16'he4aa;
    SB_LUT4 n30421_bdd_4_lut (.I0(n30421), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30424));
    defparam n30421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1129 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[4] [1]), 
            .I2(n26227), .I3(n6_adj_3712), .O(n4_adj_3737));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25331 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30415));
    defparam byte_transmit_counter_0__bdd_4_lut_25331.LUT_INIT = 16'he4aa;
    SB_LUT4 n30415_bdd_4_lut (.I0(n30415), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30418));
    defparam n30415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n14224));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(n13826), .I1(n26209), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n26590));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'h9696;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3233), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut_4_lut_adj_1132 (.I0(n13826), .I1(n26209), .I2(n10_adj_3717), 
            .I3(n26526), .O(n12002));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(n26033), .I1(n26079), .I2(n18866), 
            .I3(n6_adj_3751), .O(n17125));   // verilog/coms.v(201[5:24])
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25326 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30409));
    defparam byte_transmit_counter_0__bdd_4_lut_25326.LUT_INIT = 16'he4aa;
    SB_LUT4 n30409_bdd_4_lut (.I0(n30409), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30412));
    defparam n30409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26151));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1135 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n26164));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26353));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25321 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30391));
    defparam byte_transmit_counter_0__bdd_4_lut_25321.LUT_INIT = 16'he4aa;
    SB_LUT4 n30391_bdd_4_lut (.I0(n30391), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30394));
    defparam n30391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1137 (.I0(n14446), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n26461));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25306 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30379));
    defparam byte_transmit_counter_0__bdd_4_lut_25306.LUT_INIT = 16'he4aa;
    SB_LUT4 n30379_bdd_4_lut (.I0(n30379), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30382));
    defparam n30379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3789));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1139 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[5] [2]), 
            .I2(\data_in_frame[5] [1]), .I3(n6_adj_3789), .O(n26129));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1140 (.I0(n13915), .I1(\data_in_frame[5] [5]), 
            .I2(n26106), .I3(\data_in_frame[5] [4]), .O(n26180));
    defparam i3_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25406 (.I0(byte_transmit_counter[3]), 
            .I1(n30352), .I2(n29216), .I3(byte_transmit_counter[4]), .O(n30361));
    defparam byte_transmit_counter_3__bdd_4_lut_25406.LUT_INIT = 16'he4aa;
    SB_LUT4 n30361_bdd_4_lut (.I0(n30361), .I1(n14), .I2(n7_adj_3621), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n30361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26250));
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_CARRY add_43_4 (.CI(n21969), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n21970));
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3233), 
            .CO(n21999));
    SB_LUT4 add_43_33_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n21998), .O(n2_adj_3790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26184));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25416 (.I0(byte_transmit_counter[1]), 
            .I1(n29217), .I2(n29218), .I3(byte_transmit_counter[2]), .O(n30349));
    defparam byte_transmit_counter_1__bdd_4_lut_25416.LUT_INIT = 16'he4aa;
    SB_LUT4 n30349_bdd_4_lut (.I0(n30349), .I1(n17_adj_3619), .I2(n16_adj_3618), 
            .I3(byte_transmit_counter[2]), .O(n30352));
    defparam n30349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26256));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25296 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30343));
    defparam byte_transmit_counter_0__bdd_4_lut_25296.LUT_INIT = 16'he4aa;
    SB_LUT4 n30343_bdd_4_lut (.I0(n30343), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30346));
    defparam n30343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11_4_lut_adj_1144 (.I0(n26256), .I1(\data_in_frame[4] [1]), 
            .I2(n26113), .I3(n26184), .O(n30));   // verilog/coms.v(85[17:63])
    defparam i11_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25270 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27][0] ), 
            .I3(byte_transmit_counter[1]), .O(n30337));
    defparam byte_transmit_counter_0__bdd_4_lut_25270.LUT_INIT = 16'he4aa;
    SB_LUT4 n30337_bdd_4_lut (.I0(n30337), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30340));
    defparam n30337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15_4_lut_adj_1145 (.I0(\data_in_frame[3] [0]), .I1(n30), .I2(\data_in_frame[1] [5]), 
            .I3(n26164), .O(n34_adj_3791));   // verilog/coms.v(85[17:63])
    defparam i15_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25275 (.I0(byte_transmit_counter[1]), 
            .I1(n29220), .I2(n29221), .I3(byte_transmit_counter[2]), .O(n30331));
    defparam byte_transmit_counter_1__bdd_4_lut_25275.LUT_INIT = 16'he4aa;
    SB_LUT4 n30331_bdd_4_lut (.I0(n30331), .I1(n17_adj_3617), .I2(n16_adj_3616), 
            .I3(byte_transmit_counter[2]), .O(n30334));
    defparam n30331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13_4_lut_adj_1146 (.I0(n26250), .I1(n26157), .I2(n26180), 
            .I3(n26129), .O(n32));   // verilog/coms.v(85[17:63])
    defparam i13_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25260 (.I0(byte_transmit_counter[1]), 
            .I1(n29223), .I2(n29224), .I3(byte_transmit_counter[2]), .O(n30325));
    defparam byte_transmit_counter_1__bdd_4_lut_25260.LUT_INIT = 16'he4aa;
    SB_LUT4 n30325_bdd_4_lut (.I0(n30325), .I1(n17_adj_3615), .I2(n16_adj_3614), 
            .I3(byte_transmit_counter[2]), .O(n30328));
    defparam n30325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14_4_lut_adj_1147 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[2] [5]), .I3(n14224), .O(n33));   // verilog/coms.v(85[17:63])
    defparam i14_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25265 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30319));
    defparam byte_transmit_counter_0__bdd_4_lut_25265.LUT_INIT = 16'he4aa;
    SB_LUT4 n30319_bdd_4_lut (.I0(n30319), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30322));
    defparam n30319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1148 (.I0(n26151), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[5] [3]), .O(n31_adj_3792));   // verilog/coms.v(85[17:63])
    defparam i12_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25255 (.I0(byte_transmit_counter[1]), 
            .I1(n29229), .I2(n29230), .I3(byte_transmit_counter[2]), .O(n30313));
    defparam byte_transmit_counter_1__bdd_4_lut_25255.LUT_INIT = 16'he4aa;
    SB_LUT4 n30313_bdd_4_lut (.I0(n30313), .I1(n17_adj_3613), .I2(n16_adj_3612), 
            .I3(byte_transmit_counter[2]), .O(n30316));
    defparam n30313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i18_4_lut_adj_1149 (.I0(n31_adj_3792), .I1(n33), .I2(n32), 
            .I3(n34_adj_3791), .O(n23683));   // verilog/coms.v(85[17:63])
    defparam i18_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25245 (.I0(byte_transmit_counter[1]), 
            .I1(n29236), .I2(n29237), .I3(byte_transmit_counter[2]), .O(n30307));
    defparam byte_transmit_counter_1__bdd_4_lut_25245.LUT_INIT = 16'he4aa;
    SB_LUT4 n30307_bdd_4_lut (.I0(n30307), .I1(n17), .I2(n16), .I3(byte_transmit_counter[2]), 
            .O(n30310));
    defparam n30307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1150 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n13685));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1150.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25240 (.I0(byte_transmit_counter[1]), 
            .I1(n29239), .I2(n29240), .I3(byte_transmit_counter[2]), .O(n30301));
    defparam byte_transmit_counter_1__bdd_4_lut_25240.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_984_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n3938), .I3(GND_net), .O(n3939));
    defparam mux_984_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n14593), .D(n3940));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11495_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n15300));
    defparam i11495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11496_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n15301));
    defparam i11496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n14593), .D(n3941));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n14593), .D(n3942));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n14593), .D(n3943));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n14593), .D(n3944));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n14593), .D(n3945));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n14593), .D(n3946));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n14593), .D(n3947));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n14593), .D(n3948));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n14593), 
            .D(n3949));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n14593), 
            .D(n3950));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n14593), 
            .D(n3951));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n14593), 
            .D(n3952));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n14593), 
            .D(n3953));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n14593), 
            .D(n3954));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n14593), 
            .D(n3955));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n14593), 
            .D(n3956));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n14593), 
            .D(n3957));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n14593), 
            .D(n3958));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n14593), 
            .D(n3959));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n14593), 
            .D(n3960));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n14593), 
            .D(n3961));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n14593), 
            .D(n3962));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3793), .S(n3_adj_3611));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_32_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n21997), .O(n2_adj_3794)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11497_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n15302));
    defparam i11497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11498_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n15303));
    defparam i11498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1151 (.I0(\FRAME_MATCHER.state [1]), .I1(n17197), 
            .I2(\FRAME_MATCHER.state_31__N_2380 [1]), .I3(n3303), .O(n4));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1151.LUT_INIT = 16'h4440;
    SB_LUT4 i11499_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n15304));
    defparam i11499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11500_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n15305));
    defparam i11500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11501_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n15306));
    defparam i11501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11502_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26044), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n15307));
    defparam i11502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3757), .S(n3_adj_3610));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_75_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3650));   // verilog/coms.v(154[7:23])
    defparam equal_75_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_76_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3666));   // verilog/coms.v(154[7:23])
    defparam equal_76_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1152 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[9] [5]), .I3(GND_net), .O(n26464));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_LUT4 i11340_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n15145));
    defparam i11340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1153 (.I0(\FRAME_MATCHER.state [0]), .I1(n9_adj_3755), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n13));
    defparam i1_2_lut_3_lut_adj_1153.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1154 (.I0(\FRAME_MATCHER.state [0]), .I1(n9_adj_3755), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n4_adj_3784));
    defparam i1_2_lut_3_lut_adj_1154.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1155 (.I0(\data_out_frame[16] [5]), .I1(n13998), 
            .I2(n14360), .I3(GND_net), .O(n23654));
    defparam i1_2_lut_3_lut_adj_1155.LUT_INIT = 16'h9696;
    SB_LUT4 i24369_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3336[0]), 
            .I2(n130), .I3(tx_transmit_N_3233), .O(n29270));
    defparam i24369_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_adj_1156 (.I0(tx_active), .I1(r_SM_Main_2__N_3336[0]), 
            .I2(tx_transmit_N_3233), .I3(GND_net), .O(n807));
    defparam i1_2_lut_3_lut_adj_1156.LUT_INIT = 16'hfefe;
    SB_LUT4 i25081_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3336[0]), 
            .I2(n1_c), .I3(n63), .O(n14614));
    defparam i25081_3_lut_4_lut.LUT_INIT = 16'h10ff;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3714), .S(n3_adj_3609));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3709), .S(n3_adj_3608));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3707), .S(n3_adj_3607));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3703), .S(n3_adj_3606));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3692), .S(n3_adj_3605));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3679), .S(n3_adj_3604));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3669), .S(n3_adj_3603));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3660), .S(n3_adj_3602));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3659), .S(n3_adj_3601));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3658), .S(n3_adj_3600));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3654), .S(n3_adj_3599));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3630), .S(n3_adj_3598));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3796), .S(n3_adj_3597));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3797), .S(n3_adj_3596));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3798), .S(n3_adj_3595));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3799), .S(n3_adj_3594));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3800), .S(n3_adj_3593));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3801), .S(n3_adj_3592));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3802), .S(n3_adj_3591));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3803), .S(n3_adj_3590));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3804), .S(n3_adj_3589));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3805), .S(n3_adj_3588));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3806), .S(n3_adj_3587));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3807), .S(n3_adj_3585));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3808), .S(n3_adj_3584));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3809), .S(n3_adj_3583));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3810), .S(n3_adj_3582));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3794), .S(n3_adj_3581));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3790), .S(n3_c));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n14641), .D(n27865));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_3_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n21968), .O(n2_adj_3793)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n30301_bdd_4_lut (.I0(n30301), .I1(n17_adj_3811), .I2(n16_adj_3812), 
            .I3(byte_transmit_counter[2]), .O(n30304));
    defparam n30301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1157 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[16] [6]), .I3(\data_out_frame[14] [6]), 
            .O(n4_adj_3813));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i11487_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n15292));
    defparam i11487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11341_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n15146));
    defparam i11341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n14641), .D(n28031));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n14641), .D(n27106));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n14641), .D(n27586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n14641), .D(n27731));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n14641), .D(n27602));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n14641), .D(n26125));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n14641), .D(n27190));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n14641), .D(n24343));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n14641), .D(n26401));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n14641), .D(n27494));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n14641), .D(n26427));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n14641), .D(n26524));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n14641), .D(n26255));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n14641), .D(n27842));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_32 (.CI(n21997), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n21998));
    SB_LUT4 i11488_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n15293));
    defparam i11488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11342_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26035), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n15147));
    defparam i11342_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11489_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n15294));
    defparam i11489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1158 (.I0(n16570), .I1(n24622), .I2(n26347), 
            .I3(n13872), .O(n23877));
    defparam i2_3_lut_4_lut_adj_1158.LUT_INIT = 16'h9669;
    SB_LUT4 i11490_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n15295));
    defparam i11490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11491_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n15296));
    defparam i11491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n25515), .S(n25667));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n25669), .S(n25521));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n7_adj_3696), .S(n8_adj_3700));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n25663), .S(n25643));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n7_adj_3693), .S(n8_adj_3699));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n25673), .S(n25631));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n25675), .S(n25609));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n25677), .S(n25603));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n7_adj_3689), .S(n8_adj_3705));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n25679), .S(n25597));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n7_adj_3684), .S(n25459));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n18713), .S(n19223));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n7_adj_3683), .S(n8_adj_3704));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n18717), .S(n19225));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n25681), .S(n25591));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_3677), .S(n8_adj_3702));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n25683), .S(n25585));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n7_adj_3674), .S(n8_adj_3701));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n25685), .S(n25579));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n23166), .S(n23172));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n25687), .S(n25573));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n18719), .S(n19227));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n18721), .S(n23168));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n18723), .S(n19229));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n25689), .S(n25567));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n25691), .S(n25561));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n25693), .S(n25555));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n25671), .S(n25481));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n25695), .S(n25549));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n14614), .D(n8825[0]), .R(n14738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11492_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n15297));
    defparam i11492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11493_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n15298));
    defparam i11493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11494_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26044), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n15299));
    defparam i11494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_63_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3716));   // verilog/coms.v(154[7:23])
    defparam equal_63_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_64_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3691));   // verilog/coms.v(154[7:23])
    defparam equal_64_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1159 (.I0(\FRAME_MATCHER.state [1]), .I1(n17173), 
            .I2(n771), .I3(GND_net), .O(n3));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1159.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n133));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'heeee;
    SB_LUT4 select_320_Select_1_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n17173), .I2(\FRAME_MATCHER.state_31__N_2380 [1]), .I3(n771), 
            .O(n1));   // verilog/coms.v(127[12] 300[6])
    defparam select_320_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'h4440;
    SB_LUT4 i1_3_lut_4_lut_adj_1161 (.I0(\FRAME_MATCHER.state [1]), .I1(n17173), 
            .I2(n8604), .I3(n771), .O(n101));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1161.LUT_INIT = 16'h0040;
    SB_LUT4 i25164_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_3815));
    defparam i25164_2_lut.LUT_INIT = 16'h1111;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(n27319), 
            .D(n62_adj_3815), .R(n135));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1162 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[19] [4]), 
            .I2(n24770), .I3(n26359), .O(n6_adj_3816));
    defparam i1_2_lut_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1163 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[13] [2]), 
            .I2(n14002), .I3(GND_net), .O(n10_adj_3817));   // verilog/coms.v(85[17:63])
    defparam i2_2_lut_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1164 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26658));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h6666;
    SB_LUT4 i15383_2_lut_3_lut (.I0(n63_adj_3681), .I1(n63_c), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n92[1]));
    defparam i15383_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1165 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[10] [6]), .O(n6_adj_3818));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [3]), 
            .I2(n23828), .I3(GND_net), .O(n26334));
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1167 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n26467));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1168 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(n10_adj_3819), .I3(\data_out_frame[7] [0]), .O(n26167));   // verilog/coms.v(85[17:63])
    defparam i5_3_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1169 (.I0(\data_in_frame[12] [6]), .I1(n14294), 
            .I2(\data_in_frame[15] [0]), .I3(\data_in_frame[12] [5]), .O(n26436));
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_in_frame[10] [2]), .I1(n24206), 
            .I2(GND_net), .I3(GND_net), .O(n26544));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26520));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26652));
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1173 (.I0(\data_in_frame[15] [2]), .I1(n26652), 
            .I2(n26559), .I3(n26415), .O(n26247));
    defparam i3_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1174 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(n13670), .I3(GND_net), .O(n26086));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_31_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n21996), .O(n2_adj_3810)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_in_frame[10] [5]), .I1(n4_adj_3737), 
            .I2(GND_net), .I3(GND_net), .O(n26433));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1176 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n26126));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1177 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[11] [0]), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[8] [6]), .O(n26120));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_CARRY add_43_3 (.CI(n21968), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n21969));
    SB_CARRY add_43_31 (.CI(n21996), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n21997));
    SB_LUT4 i1_2_lut_4_lut_adj_1178 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[6] [5]), .I3(\data_out_frame[8] [6]), .O(n6_adj_3820));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1179 (.I0(\data_out_frame[24] [0]), .I1(n23661), 
            .I2(n26373), .I3(\data_out_frame[19] [6]), .O(n6_adj_3821));
    defparam i1_2_lut_4_lut_adj_1179.LUT_INIT = 16'h9669;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[20]_c [1]), .I1(n26287), 
            .I2(n26323), .I3(GND_net), .O(n11_adj_3822));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1180 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[11] [3]), 
            .I2(n26575), .I3(n6_adj_3823), .O(n26331));
    defparam i4_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_in_frame[18] [1]), .I1(n24653), 
            .I2(GND_net), .I3(GND_net), .O(n26538));
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1182 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[16] [2]), .I3(\data_out_frame[13] [7]), 
            .O(n26448));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1183 (.I0(n63_adj_3681), .I1(n63_c), .I2(n82), 
            .I3(GND_net), .O(n8604));
    defparam i1_2_lut_3_lut_adj_1183.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n13813));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1185 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[9] [3]), .I3(\data_out_frame[5] [1]), .O(n26223));
    defparam i2_3_lut_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1186 (.I0(\data_in[2] [2]), .I1(n10_adj_3668), 
            .I2(\data_in[1] [5]), .I3(\data_in[2] [6]), .O(n12));
    defparam i1_2_lut_4_lut_adj_1186.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut_4_lut_adj_1187 (.I0(n13178), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[16] [5]), .I3(n13990), .O(n26287));
    defparam i2_3_lut_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1188 (.I0(\data_in[2] [2]), .I1(n10_adj_3668), 
            .I2(\data_in[1] [5]), .I3(n97), .O(n12_adj_3680));
    defparam i1_2_lut_4_lut_adj_1188.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1189 (.I0(\FRAME_MATCHER.state [0]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n17125), .I3(\FRAME_MATCHER.state [2]), 
            .O(n17173));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1189.LUT_INIT = 16'h0002;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[18] [2]), .I1(n23458), .I2(n27637), 
            .I3(n26367), .O(n7_adj_3824));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_2_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1190 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [2]), 
            .I2(n27708), .I3(n14506), .O(n27647));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1190.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1191 (.I0(n2252), .I1(n26748), .I2(n2_adj_3752), 
            .I3(\FRAME_MATCHER.state_31__N_2380 [1]), .O(n7));
    defparam i1_3_lut_4_lut_adj_1191.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1192 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(n26323), .I3(GND_net), .O(n23796));
    defparam i1_2_lut_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1193 (.I0(\FRAME_MATCHER.state [0]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n17125), .I3(\FRAME_MATCHER.state [2]), 
            .O(n17197));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1193.LUT_INIT = 16'h0200;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[23] [0]), .I1(\data_out_frame[20] [6]), 
            .I2(n23796), .I3(n26535), .O(n8_adj_3826));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n21968));
    SB_LUT4 i11479_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n15284));
    defparam i11479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11480_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n15285));
    defparam i11480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11481_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n15286));
    defparam i11481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11482_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n15287));
    defparam i11482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1194 (.I0(n24605), .I1(n10_adj_3827), .I2(n27710), 
            .I3(n26426), .O(n26427));
    defparam i1_2_lut_4_lut_adj_1194.LUT_INIT = 16'h9669;
    SB_LUT4 i11483_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n15288));
    defparam i11483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1195 (.I0(n24055), .I1(\data_out_frame[25] [5]), 
            .I2(n27908), .I3(n26253), .O(n26255));
    defparam i1_2_lut_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1196 (.I0(\FRAME_MATCHER.state [3]), .I1(n8604), 
            .I2(n2252), .I3(n2_adj_3664), .O(n25515));
    defparam i1_3_lut_4_lut_adj_1196.LUT_INIT = 16'haa80;
    SB_LUT4 i11484_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n15289));
    defparam i11484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1197 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[8] [2]), .O(n26233));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1198 (.I0(\data_out_frame[19] [4]), .I1(n16570), 
            .I2(n24622), .I3(n26359), .O(n24632));
    defparam i1_2_lut_3_lut_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i11485_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n15290));
    defparam i11485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1199 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n17125), .I3(\FRAME_MATCHER.state [0]), 
            .O(n15));
    defparam i1_2_lut_3_lut_4_lut_adj_1199.LUT_INIT = 16'hfffd;
    SB_LUT4 i11486_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26044), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n15291));
    defparam i11486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_69_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3697));   // verilog/coms.v(154[7:23])
    defparam equal_69_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 equal_78_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3708));   // verilog/coms.v(154[7:23])
    defparam equal_78_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1200 (.I0(n2252), .I1(n26748), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n8604), .O(n25509));
    defparam i1_2_lut_3_lut_4_lut_adj_1200.LUT_INIT = 16'he0ee;
    SB_LUT4 i1_2_lut_3_lut_adj_1201 (.I0(\data_in_frame[11] [4]), .I1(n13604), 
            .I2(n26661), .I3(GND_net), .O(n6_adj_3823));
    defparam i1_2_lut_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1202 (.I0(\data_in_frame[9] [1]), .I1(n13826), 
            .I2(n26209), .I3(\data_in_frame[13] [5]), .O(n26575));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i25147_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n9_adj_3755), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [3]), 
            .O(n27319));
    defparam i25147_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 reduce_nor_260_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n17197), .I2(n63), .I3(GND_net), .O(n1_c));   // verilog/coms.v(127[12] 300[6])
    defparam reduce_nor_260_i1_2_lut_3_lut.LUT_INIT = 16'h8f8f;
    SB_LUT4 i25144_2_lut_3_lut (.I0(n13), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n135));
    defparam i25144_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_3_lut_adj_1203 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n13915));
    defparam i1_2_lut_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1204 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[14] [3]), 
            .I2(n23657), .I3(\data_in_frame[18] [6]), .O(n38_adj_3765));
    defparam i1_2_lut_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1205 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[1] [3]), .O(n26227));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i25160_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n60_adj_3828));
    defparam i25160_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i21694_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n17197), 
            .I2(n807), .I3(GND_net), .O(n26748));   // verilog/coms.v(127[12] 300[6])
    defparam i21694_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_4_lut_adj_1206 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(n26609), .O(n13890));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_30_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n21995), .O(n2_adj_3809)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1207 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(n26495), .I3(GND_net), .O(Kp_23__N_708));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1207.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1208 (.I0(n23683), .I1(n14098), .I2(n26272), 
            .I3(GND_net), .O(n24659));
    defparam i1_2_lut_3_lut_adj_1208.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1209 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(n13670), .I3(\data_in_frame[11] [1]), .O(n10_adj_3775));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_CARRY add_43_30 (.CI(n21995), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n21996));
    SB_LUT4 i1_3_lut_4_lut_adj_1210 (.I0(\FRAME_MATCHER.state [1]), .I1(n17197), 
            .I2(n8604), .I3(n807), .O(n2_adj_3663));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1210.LUT_INIT = 16'h8000;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25250 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30295));
    defparam byte_transmit_counter_0__bdd_4_lut_25250.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1211 (.I0(\data_in_frame[10] [5]), .I1(n4_adj_3737), 
            .I2(\data_in_frame[16] [7]), .I3(\data_in_frame[14] [5]), .O(n6_adj_3769));
    defparam i1_2_lut_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 n30295_bdd_4_lut (.I0(n30295), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30298));
    defparam n30295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10933_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n17129), 
            .I2(n130), .I3(n14614), .O(n14738));
    defparam i10933_3_lut_4_lut.LUT_INIT = 16'hdf00;
    SB_LUT4 select_320_Select_2_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n17173), .I2(n4452), .I3(\FRAME_MATCHER.state_31__N_2380[2] ), 
            .O(n7_adj_3));   // verilog/coms.v(127[12] 300[6])
    defparam select_320_Select_2_i7_3_lut_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 add_43_29_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n21994), .O(n2_adj_3808)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1212 (.I0(\FRAME_MATCHER.state [1]), .I1(n17173), 
            .I2(n4452), .I3(GND_net), .O(n2_adj_3752));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1212.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_1213 (.I0(n26180), .I1(\data_in_frame[7] [6]), 
            .I2(n13921), .I3(GND_net), .O(n26630));
    defparam i1_2_lut_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1214 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n10_adj_3761));   // verilog/coms.v(72[16:41])
    defparam i2_2_lut_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1215 (.I0(\FRAME_MATCHER.state [1]), .I1(n17173), 
            .I2(n8604), .I3(n4452), .O(n2_adj_3664));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1215.LUT_INIT = 16'h0080;
    SB_LUT4 equal_66_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));
    defparam equal_66_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1216 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[16] [2]), .I3(GND_net), .O(n26596));
    defparam i1_2_lut_3_lut_adj_1216.LUT_INIT = 16'h9696;
    SB_LUT4 i15450_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n19251));
    defparam i15450_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1360_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_3665));
    defparam i1360_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_4_lut_adj_1217 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[11] [3]), 
            .I2(n26445), .I3(n26089), .O(n26409));
    defparam i1_2_lut_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i11471_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n15276));
    defparam i11471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14939_2_lut_3_lut (.I0(n1656), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n18732));
    defparam i14939_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i3_3_lut_4_lut_adj_1218 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(n23654), .I3(n24657), .O(n8_adj_3830));   // verilog/coms.v(85[17:63])
    defparam i3_3_lut_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i11472_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n15277));
    defparam i11472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1219 (.I0(\data_in_frame[6] [3]), .I1(n26164), 
            .I2(n26489), .I3(GND_net), .O(n26529));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1219.LUT_INIT = 16'h9696;
    SB_LUT4 i11473_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n15278));
    defparam i11473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_29 (.CI(n21994), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n21995));
    SB_LUT4 i11474_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n15279));
    defparam i11474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11475_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n15280));
    defparam i11475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i47_2_lut (.I0(n8604), .I1(n2252), .I2(GND_net), .I3(GND_net), 
            .O(n3_adj_3661));   // verilog/coms.v(95[12:19])
    defparam i47_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1220 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n14432));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i11476_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n15281));
    defparam i11476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(n112), .I1(n101), .I2(GND_net), .I3(GND_net), 
            .O(n26074));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1222 (.I0(\data_in_frame[0] [5]), .I1(n26154), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[5] [0]), .O(n26196));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i23270_2_lut (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28332));
    defparam i23270_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1223 (.I0(n28332), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[2] [5]), .O(n30_adj_3831));
    defparam i13_4_lut_adj_1223.LUT_INIT = 16'h0010;
    SB_LUT4 i11_4_lut_adj_1224 (.I0(n25968), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[1] [1]), .O(n28_adj_3832));
    defparam i11_4_lut_adj_1224.LUT_INIT = 16'h8000;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n26987), .D(n60_adj_3828), 
            .R(n27310));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1225 (.I0(\data_in_frame[1] [3]), .I1(n13685), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[2] [6]), .O(n29_adj_3833));
    defparam i12_4_lut_adj_1225.LUT_INIT = 16'h0002;
    SB_LUT4 i10_4_lut_adj_1226 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[1] [4]), .O(n27_adj_3834));
    defparam i10_4_lut_adj_1226.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_1227 (.I0(n27_adj_3834), .I1(n29_adj_3833), .I2(n28_adj_3832), 
            .I3(n30_adj_3831), .O(\FRAME_MATCHER.state_31__N_2444 [3]));
    defparam i16_4_lut_adj_1227.LUT_INIT = 16'h8000;
    SB_LUT4 select_320_Select_2_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n17197), .I2(\FRAME_MATCHER.state_31__N_2380[2] ), .I3(n3303), 
            .O(n5));   // verilog/coms.v(127[12] 300[6])
    defparam select_320_Select_2_i5_3_lut_4_lut.LUT_INIT = 16'h4440;
    SB_LUT4 i11477_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n15282));
    defparam i11477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1228 (.I0(\FRAME_MATCHER.state_31__N_2444 [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n83), .I3(\FRAME_MATCHER.state [1]), .O(n28244));
    defparam i3_4_lut_adj_1228.LUT_INIT = 16'h0200;
    SB_LUT4 i11478_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26044), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n15283));
    defparam i11478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1229 (.I0(n28244), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n2_adj_3663), .I3(n26074), .O(n25667));
    defparam i1_4_lut_adj_1229.LUT_INIT = 16'heeea;
    SB_LUT4 add_43_28_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n21993), .O(n2_adj_3807)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11463_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n15268));
    defparam i11463_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11464_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n15269));
    defparam i11464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1230 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n14196));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_LUT4 i11465_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n15270));
    defparam i11465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11466_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n15271));
    defparam i11466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11467_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n15272));
    defparam i11467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11468_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n15273));
    defparam i11468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11469_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n15274));
    defparam i11469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_28 (.CI(n21993), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n21994));
    SB_LUT4 i11470_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26044), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n15275));
    defparam i11470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1231 (.I0(n23800), .I1(n26377), .I2(n23771), 
            .I3(GND_net), .O(n27842));
    defparam i2_3_lut_adj_1231.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1232 (.I0(n24055), .I1(\data_out_frame[25] [5]), 
            .I2(n27908), .I3(GND_net), .O(n23771));
    defparam i2_3_lut_adj_1232.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1233 (.I0(\data_out_frame[25] [4]), .I1(n14506), 
            .I2(n24055), .I3(\data_out_frame[23] [2]), .O(n26253));
    defparam i1_4_lut_adj_1233.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1234 (.I0(n26253), .I1(n26523), .I2(GND_net), 
            .I3(GND_net), .O(n26524));
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h9999;
    SB_LUT4 i11455_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n15260));
    defparam i11455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1235 (.I0(n26350), .I1(\data_out_frame[18] [4]), 
            .I2(n24657), .I3(n26508), .O(n10_adj_3827));
    defparam i4_4_lut_adj_1235.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1236 (.I0(n24605), .I1(n10_adj_3827), .I2(n27710), 
            .I3(GND_net), .O(n24645));
    defparam i5_3_lut_adj_1236.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1237 (.I0(n24645), .I1(n26281), .I2(\data_out_frame[25] [2]), 
            .I3(GND_net), .O(n27494));
    defparam i2_3_lut_adj_1237.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1238 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[24] [7]), 
            .I2(n8_adj_3826), .I3(n26284), .O(n26281));
    defparam i1_4_lut_adj_1238.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(n26281), .I1(n26399), .I2(GND_net), 
            .I3(GND_net), .O(n26401));
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1240 (.I0(n26217), .I1(\data_out_frame[19] [1]), 
            .I2(\data_out_frame[23] [3]), .I3(n26230), .O(n10_adj_3836));
    defparam i4_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1241 (.I0(n26303), .I1(n10_adj_3836), .I2(n24605), 
            .I3(GND_net), .O(n24055));
    defparam i5_3_lut_adj_1241.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1242 (.I0(n23796), .I1(n26386), .I2(n26174), 
            .I3(n13291), .O(n13_adj_3837));
    defparam i5_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1243 (.I0(n13_adj_3837), .I1(n11), .I2(n24622), 
            .I3(n26175), .O(n14506));
    defparam i7_4_lut_adj_1243.LUT_INIT = 16'h9669;
    SB_LUT4 i11456_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n15261));
    defparam i11456_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1244 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(n26297), .I3(n13221), .O(n27708));
    defparam i3_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_out_frame[20] [3]), .I1(n27708), 
            .I2(GND_net), .I3(GND_net), .O(n26535));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [0]), 
            .I2(n13670), .I3(GND_net), .O(n26259));
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i11457_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n15262));
    defparam i11457_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_1247 (.I0(\data_out_frame[20] [7]), .I1(n26110), 
            .I2(\data_out_frame[15] [7]), .I3(n26593), .O(n52));
    defparam i18_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1248 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(n13990), .O(n59));
    defparam i25_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1249 (.I0(\data_out_frame[15] [5]), .I1(n26696), 
            .I2(n24630), .I3(n26642), .O(n56));
    defparam i22_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1250 (.I0(\data_out_frame[14] [1]), .I1(n26633), 
            .I2(n26702), .I3(n26502), .O(n54));
    defparam i20_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1251 (.I0(n26241), .I1(n14240), .I2(n23824), 
            .I3(\data_out_frame[11] [5]), .O(n55));
    defparam i21_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i11458_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n15263));
    defparam i11458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[7] [1]), .I1(n26356), .I2(n26683), 
            .I3(\data_out_frame[16] [3]), .O(n53));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1252 (.I0(n26236), .I1(\data_out_frame[9] [3]), 
            .I2(n26093), .I3(\data_out_frame[10] [4]), .O(n58));
    defparam i24_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut_adj_1253 (.I0(n59), .I1(\data_out_frame[15] [0]), 
            .I2(n52), .I3(n24620), .O(n64_adj_3838));
    defparam i30_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1254 (.I0(n14446), .I1(n26467), .I2(n26568), 
            .I3(n26287), .O(n57_adj_3839));
    defparam i23_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n65_adj_3840));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n65_adj_3840), .I1(n57_adj_3839), .I2(n64_adj_3838), 
            .I3(n58), .O(n26174));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_out_frame[20] [6]), .I1(n26174), 
            .I2(GND_net), .I3(GND_net), .O(n26175));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1256 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n4_adj_3735));
    defparam i1_2_lut_3_lut_adj_1256.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26230));
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n13726));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_out_frame[20] [6]), .I1(n23796), 
            .I2(GND_net), .I3(GND_net), .O(n24657));
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i11459_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n15264));
    defparam i11459_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1260 (.I0(\data_out_frame[23] [1]), .I1(n13726), 
            .I2(n8_adj_3830), .I3(n26187), .O(n26508));
    defparam i1_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(n26508), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3841));
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1262 (.I0(\data_out_frame[20] [6]), .I1(n26230), 
            .I2(n13221), .I3(n23715), .O(n12_adj_3842));
    defparam i5_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1263 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[23] [2]), 
            .I2(n12_adj_3842), .I3(n8_adj_3841), .O(n26523));
    defparam i1_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[25] [2]), .I1(n26523), 
            .I2(GND_net), .I3(GND_net), .O(n26426));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3843));   // verilog/coms.v(97[12:26])
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[18] [3]), .I1(n24375), 
            .I2(GND_net), .I3(GND_net), .O(n26297));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1267 (.I0(n23761), .I1(n26297), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n27710));
    defparam i2_3_lut_adj_1267.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(n27708), .I1(n14506), .I2(GND_net), 
            .I3(GND_net), .O(n26187));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h9999;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n14833));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n14832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n14831));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11460_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n15265));
    defparam i11460_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1269 (.I0(\data_out_frame[24] [6]), .I1(n26535), 
            .I2(n26367), .I3(n23761), .O(n12_adj_3844));
    defparam i5_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1270 (.I0(\data_out_frame[24] [7]), .I1(n12_adj_3844), 
            .I2(n27710), .I3(\data_out_frame[25] [0]), .O(n26399));
    defparam i6_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_LUT4 i11461_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n15266));
    defparam i11461_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20_4_lut_adj_1271 (.I0(n13872), .I1(n26_adj_3843), .I2(\data_out_frame[18] [5]), 
            .I3(\data_out_frame[24] [5]), .O(n48));   // verilog/coms.v(71[16:27])
    defparam i20_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1272 (.I0(n13816), .I1(n26562), .I2(\data_out_frame[25] [1]), 
            .I3(n26426), .O(n46));   // verilog/coms.v(71[16:27])
    defparam i18_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1273 (.I0(n26350), .I1(\data_out_frame[19] [1]), 
            .I2(n26300), .I3(n26175), .O(n47));   // verilog/coms.v(71[16:27])
    defparam i19_4_lut_adj_1273.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut (.I0(n26314), .I1(\data_out_frame[20] [4]), .I2(n27647), 
            .I3(\data_out_frame[23] [4]), .O(n45));   // verilog/coms.v(71[16:27])
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11462_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26044), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n15267));
    defparam i11462_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1274 (.I0(n26289), .I1(\data_out_frame[25] [4]), 
            .I2(n16570), .I3(n26556), .O(n44));   // verilog/coms.v(71[16:27])
    defparam i16_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1275 (.I0(n23765), .I1(\data_out_frame[24] [6]), 
            .I2(n24632), .I3(\data_out_frame[25] [5]), .O(n43_adj_3845));   // verilog/coms.v(71[16:27])
    defparam i15_4_lut_adj_1275.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_27_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n21992), .O(n2_adj_3806)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11447_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n15252));
    defparam i11447_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11448_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n15253));
    defparam i11448_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11449_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n15254));
    defparam i11449_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i26_4_lut_adj_1276 (.I0(n45), .I1(n47), .I2(n46), .I3(n48), 
            .O(n54_adj_3846));   // verilog/coms.v(71[16:27])
    defparam i26_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_CARRY add_43_27 (.CI(n21992), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n21993));
    SB_LUT4 i21_4_lut_adj_1277 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[23] [7]), 
            .I2(n24055), .I3(\data_out_frame[23] [6]), .O(n49));   // verilog/coms.v(71[16:27])
    defparam i21_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i11450_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n15255));
    defparam i11450_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_43_26_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n21991), .O(n2_adj_3805)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i27_4_lut_adj_1278 (.I0(n49), .I1(n54_adj_3846), .I2(n43_adj_3845), 
            .I3(n44), .O(n24343));   // verilog/coms.v(71[16:27])
    defparam i27_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i11451_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n15256));
    defparam i11451_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(n24343), .I1(n26399), .I2(GND_net), 
            .I3(GND_net), .O(n14501));
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1280 (.I0(\data_out_frame[18] [3]), .I1(n24674), 
            .I2(\data_out_frame[20] [4]), .I3(\data_out_frame[18] [1]), 
            .O(n26284));
    defparam i3_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_CARRY add_43_26 (.CI(n21991), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n21992));
    SB_LUT4 i2_3_lut_adj_1281 (.I0(n14196), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n26145));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1281.LUT_INIT = 16'h9696;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n28285));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1282 (.I0(\data_out_frame[20] [2]), .I1(n26284), 
            .I2(n24635), .I3(n23761), .O(n27564));
    defparam i3_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n30820));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1283 (.I0(\data_out_frame[24] [6]), .I1(n26123), 
            .I2(n27564), .I3(n14501), .O(n27190));
    defparam i3_4_lut_adj_1283.LUT_INIT = 16'h9669;
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n15337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n15336));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11452_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n15257));
    defparam i11452_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n15335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n15334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n15333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n15332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n15331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n15330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n15329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n15328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n15327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n15326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n15325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n15324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n15323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n15322));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n15321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n15320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n15319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n15318));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n15317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n15316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n15315));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n15314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n15313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n15312));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11453_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n15258));
    defparam i11453_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1284 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n26356));
    defparam i2_3_lut_adj_1284.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1285 (.I0(n24601), .I1(n26550), .I2(n26356), 
            .I3(n13970), .O(n24635));
    defparam i3_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n15311));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11454_3_lut_4_lut (.I0(n19251), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n15259));
    defparam i11454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26244));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n15310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n15309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n15308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n15307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n15306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n15305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n15304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n15303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n15302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n15301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n15300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n15299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n15298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n15297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n15296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n15295));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11439_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n15244));
    defparam i11439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n15294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n15293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n15292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n15291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n15290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n15289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n15288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n15287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n15286));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n15285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n15284));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_out_frame[20] [2]), .I1(n24635), 
            .I2(GND_net), .I3(GND_net), .O(n26367));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h9999;
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n15283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n15282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n15281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n15280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n15279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n15278));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_out_frame[18] [2]), .I1(n23458), 
            .I2(GND_net), .I3(GND_net), .O(n23761));
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n15277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n15276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n15275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n15274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n15273));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n15272));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n15271));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n15270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n15269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n15268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n15267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n15266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n15265));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1289 (.I0(n7_adj_3824), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[24] [5]), .I3(n24607), .O(n26123));
    defparam i4_4_lut_adj_1289.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n15264));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_25_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n21990), .O(n2_adj_3804)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n15263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n15262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n15261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n15260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n15259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n15258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n15257));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1290 (.I0(n23765), .I1(n26123), .I2(GND_net), 
            .I3(GND_net), .O(n26125));
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n15256));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11440_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n15245));
    defparam i11440_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n15255));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_out_frame[18] [0]), .I1(n24722), 
            .I2(GND_net), .I3(GND_net), .O(n26550));
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h9999;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n15254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n15253));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n15252));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n15251));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n15250));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_25 (.CI(n21990), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n21991));
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n15249));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_out_frame[20] [2]), .I1(n26550), 
            .I2(n26317), .I3(\data_out_frame[18] [1]), .O(n10_adj_3657));
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i11441_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n15246));
    defparam i11441_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1293 (.I0(n13826), .I1(n26190), .I2(n26689), 
            .I3(GND_net), .O(n6_adj_3733));
    defparam i1_2_lut_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1294 (.I0(\data_out_frame[24] [4]), .I1(n24607), 
            .I2(n27637), .I3(n27795), .O(n23765));
    defparam i1_4_lut_adj_1294.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(n26209), .I3(GND_net), .O(n26190));
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1296 (.I0(Kp_23__N_1026), .I1(n13882), .I2(n13890), 
            .I3(\data_in_frame[10] [0]), .O(n23828));
    defparam i1_2_lut_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(n14336), .I1(n26099), .I2(GND_net), 
            .I3(GND_net), .O(n24601));
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1298 (.I0(n26505), .I1(n14336), .I2(\data_out_frame[16] [0]), 
            .I3(GND_net), .O(n8_adj_3847));
    defparam i3_3_lut_adj_1298.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1299 (.I0(n13788), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3848));
    defparam i2_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1300 (.I0(n24614), .I1(\data_out_frame[15] [7]), 
            .I2(n7_adj_3848), .I3(n8_adj_3847), .O(n26317));
    defparam i2_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1301 (.I0(n13826), .I1(n26500), .I2(n23701), 
            .I3(n14289), .O(n26343));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n15248));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n15247));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n15246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n15245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n15244));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n15243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n15242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n15241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n15240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n15239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n15238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n15237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n15236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n15235));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n15234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n15233));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n15232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n15231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n15230));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n15229));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n15228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n15227));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n15226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n15225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n15224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n15223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n15222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n15221));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n15220));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n15219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n15218));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n15217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n15216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n15215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n15214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n15213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n15212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n15211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n15210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n15209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n15208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n15207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n15206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n15205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n15204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n15203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n15202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n15201));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n15200));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n15199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n15198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n15197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n15196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n15195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n15194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n15193));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n15192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n15191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n15190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n15189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n15188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n15187));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n15186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n15185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n15184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n15183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n15182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n15181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n15180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n15179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n15178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n15177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n15176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n15175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n15174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n15173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n15172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n15171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n15170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n15169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n15168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n15167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n15166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n15165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n15164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n15163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n15162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n15161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n15160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n15159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n15158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n15157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n15156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n15155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n15154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n15153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n15152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n15151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n15150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n15149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n15148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n15147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n15146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n15145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n15144));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n15143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n15142));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n15141));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11442_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n15247));
    defparam i11442_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(n26680), .I1(\data_out_frame[16] [1]), 
            .I2(n26099), .I3(n26615), .O(n15_adj_3849));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1303 (.I0(n15_adj_3849), .I1(n26448), .I2(n14_adj_3655), 
            .I3(\data_out_frame[9] [6]), .O(n24375));   // verilog/coms.v(76[16:43])
    defparam i8_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i11443_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n15248));
    defparam i11443_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1304 (.I0(n24375), .I1(n26317), .I2(n24601), 
            .I3(\data_out_frame[17] [7]), .O(n24674));
    defparam i3_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1305 (.I0(n13974), .I1(n26223), .I2(\data_out_frame[11] [5]), 
            .I3(GND_net), .O(n26505));
    defparam i2_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26683));
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26615));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1308 (.I0(\data_out_frame[13] [7]), .I1(n26683), 
            .I2(n26461), .I3(n26505), .O(n12_adj_3850));
    defparam i5_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1309 (.I0(n26454), .I1(n12_adj_3850), .I2(\data_out_frame[16] [3]), 
            .I3(n26615), .O(n26217));
    defparam i6_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i11444_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n15249));
    defparam i11444_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11445_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n15250));
    defparam i11445_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1310 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[13] [7]), .I3(GND_net), .O(n26702));   // verilog/coms.v(97[12:26])
    defparam i2_3_lut_adj_1310.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26502));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3851));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1313 (.I0(n26502), .I1(\data_out_frame[6] [6]), 
            .I2(n26223), .I3(n4_adj_3851), .O(n14336));
    defparam i2_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1314 (.I0(n26448), .I1(n26600), .I2(n14336), 
            .I3(\data_out_frame[14] [0]), .O(n12_adj_3852));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1315 (.I0(\data_out_frame[16] [3]), .I1(n12_adj_3852), 
            .I2(n26674), .I3(n14446), .O(n13221));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1316 (.I0(n23701), .I1(n13890), .I2(n26423), 
            .I3(\data_in_frame[9] [4]), .O(n14429));
    defparam i2_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i11446_3_lut_4_lut (.I0(n8), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n15251));
    defparam i11446_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1317 (.I0(\data_in_frame[11] [6]), .I1(n23701), 
            .I2(n14289), .I3(\data_in_frame[9] [5]), .O(n26423));
    defparam i2_3_lut_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_out_frame[20]_c [1]), .I1(n26287), 
            .I2(GND_net), .I3(GND_net), .O(n26562));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1319 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[14] [0]), .I3(\data_out_frame[13] [5]), 
            .O(n26593));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1320 (.I0(n26442), .I1(n26593), .I2(\data_out_frame[11] [6]), 
            .I3(\data_out_frame[13] [6]), .O(n12_adj_3853));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1321 (.I0(\data_out_frame[13] [7]), .I1(n12_adj_3853), 
            .I2(n26668), .I3(\data_out_frame[15] [6]), .O(n23458));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1322 (.I0(n23654), .I1(n26373), .I2(\data_out_frame[18] [0]), 
            .I3(n23458), .O(n13_adj_3854));
    defparam i5_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25231 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30289));
    defparam byte_transmit_counter_0__bdd_4_lut_25231.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1323 (.I0(n13_adj_3854), .I1(n11_adj_3822), .I2(n24674), 
            .I3(\data_out_frame[19] [7]), .O(n24607));
    defparam i7_4_lut_adj_1323.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1324 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[20] [0]), 
            .I2(n26413), .I3(n23661), .O(n26300));
    defparam i3_4_lut_adj_1324.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1325 (.I0(\data_out_frame[19] [6]), .I1(n26300), 
            .I2(n24607), .I3(GND_net), .O(n27795));
    defparam i2_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1326 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n13816));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1326.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1327 (.I0(\data_in_frame[16] [0]), .I1(n23664), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n26661));
    defparam i1_2_lut_3_lut_adj_1327.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1328 (.I0(\data_in_frame[13] [2]), .I1(n12002), 
            .I2(\data_in_frame[11] [1]), .I3(\data_in_frame[10] [7]), .O(n26636));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(\data_out_frame[24] [1]), .I1(n23877), 
            .I2(GND_net), .I3(GND_net), .O(n26289));
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1330 (.I0(n28172), .I1(n26289), .I2(\data_out_frame[24] [2]), 
            .I3(GND_net), .O(n27586));
    defparam i2_3_lut_adj_1330.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1331 (.I0(\data_out_frame[24] [1]), .I1(n23824), 
            .I2(n26311), .I3(n6_adj_3821), .O(n27106));
    defparam i4_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n13872));
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1333 (.I0(\data_out_frame[19] [3]), .I1(n24622), 
            .I2(n23824), .I3(GND_net), .O(n26359));
    defparam i2_3_lut_adj_1333.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1334 (.I0(\data_out_frame[23] [5]), .I1(\data_out_frame[19] [1]), 
            .I2(n26359), .I3(n13236), .O(n23800));
    defparam i1_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1335 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n13974));
    defparam i2_3_lut_adj_1335.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1336 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n26093));
    defparam i2_3_lut_adj_1336.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1337 (.I0(n26621), .I1(n26320), .I2(\data_out_frame[7] [0]), 
            .I3(n6_adj_3820), .O(n26442));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n15140));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n15139));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n15138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n15137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n15136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n15135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n15134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n15133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n15132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n15131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n15130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n15129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n15128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n15127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n15126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n15125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n15124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n15123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n15122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n15121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n15120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n15119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n15118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n15117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n15116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n15115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n15114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n15113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n15112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n15111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n15110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i217 (.Q(\data_out_frame[27][0] ), .C(clk32MHz), 
           .D(n15109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n15108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n15107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n15106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n15105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n15104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n15103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n15102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n15101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n15100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n15099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n15098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n15097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n15096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n15095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n15094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n15093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n15092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n15091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n15090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n15089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n15088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n15087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n15086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n15085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n15084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n15083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n15082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n15081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n15080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n15079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20]_c [1]), .C(clk32MHz), 
           .D(n15078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n15077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n15076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n15075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n15074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n15073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n15072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n15071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n15070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n15069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n15068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n15067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n15066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n15065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n15064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n15063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n15062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n15061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n15060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n15059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n15058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n15057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n15056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n15055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n15054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n15053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n15052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n15051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n15050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n15049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n15048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n15047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n15046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n15045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n15044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n15043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n15042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n15041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n15040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n15039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n15038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n15037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n15036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n15035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n15034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n15033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n15032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n15031));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n15030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n15029));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n15028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n15027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n15026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n15025));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1338 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[9] [1]), .I3(n13974), .O(n27993));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1339 (.I0(n14289), .I1(n26500), .I2(n23701), 
            .I3(n13890), .O(n26581));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_816), 
            .I2(\data_in_frame[8] [5]), .I3(GND_net), .O(n6_adj_3748));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1341 (.I0(\data_out_frame[15] [5]), .I1(n24722), 
            .I2(n26167), .I3(GND_net), .O(n24614));
    defparam i1_3_lut_adj_1341.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_816), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n6_adj_3710));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1343 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3855));
    defparam i2_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1344 (.I0(n7_adj_3855), .I1(\data_out_frame[20] [0]), 
            .I2(n16570), .I3(n26413), .O(n26347));
    defparam i4_4_lut_adj_1344.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26532));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26320));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1347 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[15] [2]), .I3(\data_out_frame[12] [6]), 
            .O(n26642));   // verilog/coms.v(97[12:26])
    defparam i3_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_24_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n21989), .O(n2_adj_3803)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26696));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i11431_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n15236));
    defparam i11431_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1349 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n26621));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1349.LUT_INIT = 16'h9696;
    SB_CARRY add_43_24 (.CI(n21989), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n21990));
    SB_LUT4 i4_4_lut_adj_1350 (.I0(\data_out_frame[13] [3]), .I1(n26621), 
            .I2(n26126), .I3(\data_out_frame[10] [7]), .O(n10_adj_3819));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26269));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(\data_out_frame[11] [1]), .I1(n26120), 
            .I2(n26532), .I3(n6_adj_3818), .O(n14011));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i11432_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n15237));
    defparam i11432_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11433_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n15238));
    defparam i11433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1353 (.I0(n14011), .I1(n26167), .I2(\data_out_frame[15] [4]), 
            .I3(GND_net), .O(n13970));
    defparam i2_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1354 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n14_adj_3856));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1355 (.I0(n13970), .I1(n14011), .I2(n26467), 
            .I3(\data_out_frame[5] [7]), .O(n15_adj_3857));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n15024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n15023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n15022));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11434_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n15239));
    defparam i11434_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1356 (.I0(n15_adj_3857), .I1(n26618), .I2(n14_adj_3856), 
            .I3(n26120), .O(n26373));   // verilog/coms.v(74[16:27])
    defparam i8_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n15021));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1357 (.I0(n26642), .I1(\data_out_frame[11] [0]), 
            .I2(n26320), .I3(\data_out_frame[13] [0]), .O(n14_adj_3858));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n15020));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1358 (.I0(\data_out_frame[17] [4]), .I1(n14_adj_3858), 
            .I2(n10_adj_3817), .I3(n26126), .O(n23661));   // verilog/coms.v(85[17:63])
    defparam i7_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1359 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n13538), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_3682));
    defparam i1_3_lut_4_lut_adj_1359.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(n23661), .I1(n16570), .I2(GND_net), 
            .I3(GND_net), .O(n13291));
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1361 (.I0(n26217), .I1(\data_out_frame[16] [4]), 
            .I2(n13178), .I3(n13221), .O(n26323));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i11435_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n15240));
    defparam i11435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1362 (.I0(n26402), .I1(n13291), .I2(\data_out_frame[23] [7]), 
            .I3(n6_adj_3816), .O(n28172));
    defparam i4_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1363 (.I0(n23800), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n26314));
    defparam i2_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i11436_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n15241));
    defparam i11436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1364 (.I0(n23877), .I1(n26314), .I2(n28172), 
            .I3(n24737), .O(n28031));
    defparam i3_4_lut_adj_1364.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3812));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1365 (.I0(n13503), .I1(n11166), .I2(n31_adj_3653), 
            .I3(GND_net), .O(n27156));
    defparam i2_3_lut_adj_1365.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3811));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1366 (.I0(n13998), .I1(n24314), .I2(\data_out_frame[16] [6]), 
            .I3(n23654), .O(n24630));
    defparam i1_2_lut_3_lut_4_lut_adj_1366.LUT_INIT = 16'h9669;
    SB_LUT4 i11437_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n15242));
    defparam i11437_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1367 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n26200));
    defparam i2_3_lut_adj_1367.LUT_INIT = 16'h9696;
    SB_LUT4 i11438_3_lut_4_lut (.I0(n8_adj_3650), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n15243));
    defparam i11438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_23_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n21988), .O(n2_adj_3802)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1368 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26639));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1368.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1369 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[13] [0]), .I3(\data_out_frame[15] [1]), 
            .O(n26633));
    defparam i3_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26470));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'h6666;
    SB_CARRY add_43_23 (.CI(n21988), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n21989));
    SB_LUT4 i2_3_lut_adj_1371 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26618));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1372 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n8_adj_3859));
    defparam i3_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1373 (.I0(\data_out_frame[10] [2]), .I1(n24463), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3860));
    defparam i2_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1374 (.I0(\data_out_frame[12] [7]), .I1(n7_adj_3860), 
            .I2(\data_out_frame[7] [7]), .I3(n8_adj_3859), .O(n8_adj_3861));
    defparam i3_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1375 (.I0(n26470), .I1(\data_out_frame[10] [5]), 
            .I2(n8_adj_3861), .I3(n26193), .O(n6_adj_3862));
    defparam i1_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1376 (.I0(n26633), .I1(n26511), .I2(n26639), 
            .I3(n6_adj_3862), .O(n24622));
    defparam i4_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1377 (.I0(\data_out_frame[15] [1]), .I1(n26236), 
            .I2(\data_out_frame[13] [1]), .I3(n26618), .O(n16_adj_3863));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1378 (.I0(\data_out_frame[7] [7]), .I1(n26584), 
            .I2(n26686), .I3(n26200), .O(n17_adj_3864));   // verilog/coms.v(85[17:63])
    defparam i7_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1379 (.I0(n17_adj_3864), .I1(\data_out_frame[6] [1]), 
            .I2(n16_adj_3863), .I3(\data_out_frame[5] [5]), .O(n27507));   // verilog/coms.v(85[17:63])
    defparam i9_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1380 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(n27507), .I3(\data_out_frame[14] [7]), .O(n16570));   // verilog/coms.v(97[12:26])
    defparam i6_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1381 (.I0(n16570), .I1(n24622), .I2(GND_net), 
            .I3(GND_net), .O(n24770));
    defparam i1_2_lut_adj_1381.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1382 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[19] [2]), 
            .I2(n26303), .I3(GND_net), .O(n26311));
    defparam i2_3_lut_adj_1382.LUT_INIT = 16'h6969;
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n15019));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11423_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n15228));
    defparam i11423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1383 (.I0(n9_adj_3755), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n88), .I3(\FRAME_MATCHER.state [1]), .O(n19405));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1383.LUT_INIT = 16'hfefb;
    SB_LUT4 i11424_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n15229));
    defparam i11424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1384 (.I0(n13998), .I1(n24314), .I2(GND_net), 
            .I3(GND_net), .O(n24620));
    defparam i1_2_lut_adj_1384.LUT_INIT = 16'h6666;
    SB_LUT4 i11425_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n15230));
    defparam i11425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1385 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n26241));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26603));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n15018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n15017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n15016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n15015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n15014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n15013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n15012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n15011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n15010));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n15009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n15008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n15007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n15006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n15005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n15004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n15003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n15002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n15001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n15000));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n14999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n14998));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n14997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n14996));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n14995));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n14994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n14993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n14992));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n14991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n14990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n14989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n14830));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11426_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n15231));
    defparam i11426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n14829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n14828));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n14827));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n14988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n14987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n14986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n14985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n14984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n14983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n14982));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11427_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n15232));
    defparam i11427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n14818));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n14981));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n14980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n14979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n14978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n14977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n14976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n14975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n14974));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1387 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[10] [3]), .O(n26584));
    defparam i1_2_lut_3_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n14973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n14972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n14971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n14970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n14969));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n14968));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n14967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n14966));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n14965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n14964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n14963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n14962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n14961));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1388 (.I0(n26603), .I1(\data_out_frame[5] [6]), 
            .I2(n26102), .I3(\data_out_frame[7] [4]), .O(n14_adj_3865));
    defparam i6_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1389 (.I0(\data_out_frame[14] [4]), .I1(n14_adj_3865), 
            .I2(n10), .I3(n26083), .O(n13998));
    defparam i7_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i11428_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n15233));
    defparam i11428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1390 (.I0(n26193), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[10] [4]), .I3(\data_out_frame[6] [0]), .O(n14002));
    defparam i3_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_22_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n21987), .O(n2_adj_3801)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n14960));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1391 (.I0(\data_out_frame[7] [6]), .I1(n26665), 
            .I2(\data_out_frame[8] [0]), .I3(\data_out_frame[6] [0]), .O(n26511));
    defparam i3_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n14959));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11429_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n15234));
    defparam i11429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_1392 (.I0(n26511), .I1(n14002), .I2(n13998), 
            .I3(GND_net), .O(n8_adj_3866));
    defparam i3_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i11430_3_lut_4_lut (.I0(n8_adj_3666), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n15235));
    defparam i11430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1393 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(n26170), .O(n26495));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n26489));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(n13685), .I3(GND_net), .O(n6_adj_3652));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1396 (.I0(n26603), .I1(n4_adj_3813), .I2(n8_adj_3866), 
            .I3(n26677), .O(n26303));   // verilog/coms.v(85[17:28])
    defparam i2_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1397 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n14192));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n14958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n14957));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n14956));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1398 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[8] [3]), .O(n26193));
    defparam i1_2_lut_3_lut_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n14955));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n14954));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_22 (.CI(n21987), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n21988));
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n14953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n14952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n14951));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1399 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[4] [2]), .O(n26113));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i11415_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n15220));
    defparam i11415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_21_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n21986), .O(n2_adj_3800)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(n13998), .I1(n14360), .I2(GND_net), 
            .I3(GND_net), .O(n13990));
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'h6666;
    SB_LUT4 i11416_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n15221));
    defparam i11416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11417_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n15222));
    defparam i11417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1401 (.I0(n24630), .I1(n26303), .I2(\data_out_frame[18] [7]), 
            .I3(GND_net), .O(n13236));
    defparam i2_3_lut_adj_1401.LUT_INIT = 16'h6969;
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n14950));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11418_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n15223));
    defparam i11418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26211));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h6666;
    SB_LUT4 i11419_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n15224));
    defparam i11419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1403 (.I0(\data_out_frame[9] [4]), .I1(n26211), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[5] [2]), .O(n13788));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i11420_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n15225));
    defparam i11420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26600));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1405 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[1] [3]), .O(n6_adj_3651));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i11421_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n15226));
    defparam i11421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11422_3_lut_4_lut (.I0(n8_adj_3697), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n15227));
    defparam i11422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1406 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26116));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1406.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26680));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1408 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[9] [7]), .O(n14446));   // verilog/coms.v(74[16:27])
    defparam i1_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i11407_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n15212));
    defparam i11407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_21 (.CI(n21986), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n21987));
    SB_LUT4 i11408_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n15213));
    defparam i11408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11409_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n15214));
    defparam i11409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26102));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n17125), .I3(GND_net), .O(n83));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'hfefe;
    SB_LUT4 i11410_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n15215));
    defparam i11410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1411 (.I0(n26110), .I1(n26461), .I2(\data_out_frame[14] [3]), 
            .I3(\data_out_frame[9] [6]), .O(n12_adj_3867));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n14949));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n14948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n14947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n14946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n14945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n14944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n14943));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n14942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n14941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n14940));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n14939));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n14938));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11411_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n15216));
    defparam i11411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1412 (.I0(\data_out_frame[8] [0]), .I1(n12_adj_3867), 
            .I2(n26612), .I3(\data_out_frame[7] [3]), .O(n14360));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n14937));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11412_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n15217));
    defparam i11412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n14936));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n14935));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n14934));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n14933));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n14932));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n14931));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n14930));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n14929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n14928));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1413 (.I0(n13788), .I1(\data_out_frame[5] [3]), 
            .I2(n26464), .I3(\data_out_frame[7] [4]), .O(n26668));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i11413_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n15218));
    defparam i11413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1414 (.I0(n26668), .I1(n26454), .I2(n14360), 
            .I3(n26674), .O(n10_adj_3868));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i11414_3_lut_4_lut (.I0(n8_adj_3708), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n15219));
    defparam i11414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1415 (.I0(n14446), .I1(n10_adj_3868), .I2(\data_out_frame[12] [0]), 
            .I3(GND_net), .O(n13178));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_LUT4 i11399_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n15204));
    defparam i11399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11400_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n15205));
    defparam i11400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1416 (.I0(\data_out_frame[16] [4]), .I1(n13178), 
            .I2(GND_net), .I3(GND_net), .O(n23715));
    defparam i1_2_lut_adj_1416.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1417 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(n26157));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1418 (.I0(\data_in_frame[21] [7]), .I1(n26275), 
            .I2(n24414), .I3(GND_net), .O(n27369));
    defparam i2_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i11401_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n15206));
    defparam i11401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26236));
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'h6666;
    SB_LUT4 i11402_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n15207));
    defparam i11402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26686));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1421 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26612));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1421.LUT_INIT = 16'h6666;
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n14927));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n14926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n14925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n14924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n14923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n14922));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1422 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n26665));
    defparam i2_3_lut_adj_1422.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n14921));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n14920));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n14919));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11403_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n15208));
    defparam i11403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n14918));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n14917));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n14916));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1423 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n14240));
    defparam i1_2_lut_adj_1423.LUT_INIT = 16'h6666;
    SB_LUT4 i11404_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n15209));
    defparam i11404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n30289_bdd_4_lut (.I0(n30289), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30292));
    defparam n30289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1424 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26482));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1424.LUT_INIT = 16'h6666;
    SB_LUT4 i11405_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n15210));
    defparam i11405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11406_3_lut_4_lut (.I0(n8_adj_3716), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n15211));
    defparam i11406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25226 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30283));
    defparam byte_transmit_counter_0__bdd_4_lut_25226.LUT_INIT = 16'he4aa;
    SB_LUT4 i11391_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n15196));
    defparam i11391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n30283_bdd_4_lut (.I0(n30283), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30286));
    defparam n30283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_4_lut_adj_1425 (.I0(n23824), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[19] [2]), .I3(n26303), .O(n7_c));
    defparam i2_2_lut_4_lut_adj_1425.LUT_INIT = 16'h9669;
    SB_LUT4 i25076_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n9_adj_3755), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n88), .O(n14641));   // verilog/coms.v(127[12] 300[6])
    defparam i25076_2_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_adj_1426 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3869));
    defparam i1_2_lut_adj_1426.LUT_INIT = 16'h6666;
    SB_LUT4 i11392_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n15197));
    defparam i11392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1427 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[8] [0]), .I3(n6_adj_3869), .O(n26083));
    defparam i4_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1428 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26514));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1428.LUT_INIT = 16'h6666;
    SB_LUT4 i11393_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n15198));
    defparam i11393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11394_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n15199));
    defparam i11394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n14915));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n14914));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n14913));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_20_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n21985), .O(n2_adj_3799)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n14912));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_20 (.CI(n21985), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n21986));
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n14911));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1429 (.I0(n26083), .I1(n26584), .I2(\data_out_frame[14] [5]), 
            .I3(\data_out_frame[6] [1]), .O(n12_adj_3870));
    defparam i5_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n14910));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_19_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n21984), .O(n2_adj_3798)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n14909));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n14908));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n14907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n14906));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1430 (.I0(\data_out_frame[7] [5]), .I1(n12_adj_3870), 
            .I2(n26665), .I3(\data_out_frame[10] [1]), .O(n24314));
    defparam i6_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n14905));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n14904));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n14903));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11395_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n15200));
    defparam i11395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n14902));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n14901));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11396_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n15201));
    defparam i11396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1431 (.I0(n26686), .I1(\data_out_frame[15] [0]), 
            .I2(\data_out_frame[8] [2]), .I3(n26677), .O(n15_adj_3871));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1432 (.I0(n15_adj_3871), .I1(n26514), .I2(n14_adj_3788), 
            .I3(\data_out_frame[8] [4]), .O(n24463));   // verilog/coms.v(85[17:63])
    defparam i8_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1433 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(n24463), .I3(n24314), .O(n23824));
    defparam i1_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i12779_3_lut (.I0(\data_out_frame[20]_c [1]), .I1(\displacement[1] ), 
            .I2(n10896), .I3(GND_net), .O(n15078));
    defparam i12779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1434 (.I0(\data_out_frame[19] [0]), .I1(n13236), 
            .I2(n4_adj_3787), .I3(n23654), .O(n26386));
    defparam i2_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n14900));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11397_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n15202));
    defparam i11397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11398_3_lut_4_lut (.I0(n8_adj_3691), .I1(n26057), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n15203));
    defparam i11398_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1435 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[19] [2]), 
            .I2(n26386), .I3(n23824), .O(n27908));
    defparam i3_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i11383_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n15188));
    defparam i11383_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(\data_out_frame[25] [6]), .I1(n27908), 
            .I2(GND_net), .I3(GND_net), .O(n26377));
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'h9999;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n14899));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n14898));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n14897));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n14896));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_19 (.CI(n21984), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n21985));
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n14895));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11384_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n15189));
    defparam i11384_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n14894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n14893));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1437 (.I0(n26164), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[4] [2]), .O(n14279));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_18_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n21983), .O(n2_adj_3797)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n14892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n14891));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n14890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n14889));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_18 (.CI(n21983), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n21984));
    SB_LUT4 i11385_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n15190));
    defparam i11385_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n14888));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n14887));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11386_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n15191));
    defparam i11386_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n14886));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_17_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n21982), .O(n2_adj_3796)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_3_lut_4_lut_adj_1438 (.I0(\FRAME_MATCHER.state [1]), .I1(n83), 
            .I2(n1656), .I3(\FRAME_MATCHER.state [2]), .O(n2272));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1438.LUT_INIT = 16'h0f0e;
    SB_LUT4 i11387_3_lut_4_lut (.I0(n19251), .I1(n26035), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n15192));
    defparam i11387_3_lut_4_lut.LUT_INIT = 16'hfd20;
    uart_tx tx (.n26856(n26856), .clk32MHz(clk32MHz), .n26880(n26880), 
            .\r_SM_Main_2__N_3336[0] (r_SM_Main_2__N_3336[0]), .r_SM_Main({r_SM_Main}), 
            .\r_SM_Main_2__N_3333[1] (\r_SM_Main_2__N_3333[1] ), .GND_net(GND_net), 
            .tx_o(tx_o), .tx_data({tx_data}), .n14872(n14872), .VCC_net(VCC_net), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n7375(n7375), .n14835(n14835), 
            .tx_active(tx_active), .n4(n4_adj_4), .n30875(n30875), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.n14672(n14672), .clk32MHz(clk32MHz), .n14766(n14766), 
            .\r_SM_Main_2__N_3262[2] (\r_SM_Main_2__N_3262[2] ), .r_SM_Main({r_SM_Main_adj_12}), 
            .n26029(n26029), .GND_net(GND_net), .r_Rx_Data(r_Rx_Data), 
            .RX_N_2(RX_N_2), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_8 ), 
            .n13551(n13551), .n4(n4_adj_9), .VCC_net(VCC_net), .n15342(n15342), 
            .n25777(n25777), .rx_data_ready(rx_data_ready), .n15346(n15346), 
            .rx_data({rx_data}), .n18789(n18789), .n4_adj_1(n4_adj_10), 
            .n4_adj_2(n4_adj_11), .n13556(n13556), .n14826(n14826), .n14825(n14825), 
            .n14824(n14824), .n14823(n14823), .n14822(n14822), .n14821(n14821), 
            .n14820(n14820)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n26856, clk32MHz, n26880, \r_SM_Main_2__N_3336[0] , 
            r_SM_Main, \r_SM_Main_2__N_3333[1] , GND_net, tx_o, tx_data, 
            n14872, VCC_net, \r_Bit_Index[0] , n7375, n14835, tx_active, 
            n4, n30875, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output n26856;
    input clk32MHz;
    output n26880;
    input \r_SM_Main_2__N_3336[0] ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3333[1] ;
    input GND_net;
    output tx_o;
    input [7:0]tx_data;
    input n14872;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n7375;
    input n14835;
    output tx_active;
    output n4;
    input n30875;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [8:0]n41;
    
    wire n4063;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n14749, n19210, n8772, n8773, n30484, n30376, o_Tx_Serial_N_3364, 
        n3, n10886;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n10, n27095, n3_adj_3580, n30481, n30373, n22424, n22423, 
        n22422, n22421, n22420, n22419, n22418, n22417;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n26856), 
            .D(n307[2]), .R(n26880));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n26856), 
            .D(n307[1]), .R(n26880));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1127__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n4063), .D(n41[8]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n4063), .D(n41[7]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n4063), .D(n41[6]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n4063), .D(n41[5]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n4063), .D(n41[4]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n4063), .D(n41[3]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n4063), .D(n41[2]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1127__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n4063), .D(n41[1]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i5037_4_lut (.I0(\r_SM_Main_2__N_3336[0] ), .I1(n19210), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3333[1] ), .O(n8772));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5037_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i5038_3_lut (.I0(n8772), .I1(\r_SM_Main_2__N_3333[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n8773));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5038_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1572264_i1_3_lut (.I0(n30484), .I1(n30376), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3364));
    defparam i1572264_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3364), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n4063), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n8773), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .E(VCC_net), 
            .D(n14872));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1127__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n4063), .D(n41[0]), .R(n14749));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i25141_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3333[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n14749));
    defparam i25141_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1055_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4063));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1055_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1210_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1210_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n27095));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n27095), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3333[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n19210));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i25180_3_lut (.I0(n26856), .I1(n19210), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n26880));
    defparam i25180_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1217_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1217_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i6953_2_lut_3_lut (.I0(\r_SM_Main_2__N_3333[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3580));
    defparam i6953_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i3652_2_lut (.I0(\r_SM_Main_2__N_3336[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n7375));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i3652_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n30481));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30481_bdd_4_lut (.I0(n30481), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n30484));
    defparam n30481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_25381 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n30373));
    defparam r_Bit_Index_0__bdd_4_lut_25381.LUT_INIT = 16'he4aa;
    SB_LUT4 n30373_bdd_4_lut (.I0(n30373), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n30376));
    defparam n30373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3336[0] ), 
            .I3(r_SM_Main[1]), .O(n10886));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i25185_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3333[1] ), .O(n26856));
    defparam i25185_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n10886), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3580), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1127_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n22424), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1127_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n22423), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_9 (.CI(n22423), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n22424));
    SB_LUT4 r_Clock_Count_1127_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n22422), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_8 (.CI(n22422), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n22423));
    SB_LUT4 r_Clock_Count_1127_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n22421), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_7 (.CI(n22421), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n22422));
    SB_LUT4 r_Clock_Count_1127_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n22420), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n14835));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY r_Clock_Count_1127_add_4_6 (.CI(n22420), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n22421));
    SB_LUT4 r_Clock_Count_1127_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n22419), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_5 (.CI(n22419), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n22420));
    SB_LUT4 r_Clock_Count_1127_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n22418), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_4 (.CI(n22418), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n22419));
    SB_LUT4 r_Clock_Count_1127_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n22417), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_3 (.CI(n22417), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n22418));
    SB_LUT4 r_Clock_Count_1127_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1127_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1127_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n22417));
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3333[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n30875));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n14672, clk32MHz, n14766, \r_SM_Main_2__N_3262[2] , 
            r_SM_Main, n26029, GND_net, r_Rx_Data, RX_N_2, \r_Bit_Index[0] , 
            n13551, n4, VCC_net, n15342, n25777, rx_data_ready, 
            n15346, rx_data, n18789, n4_adj_1, n4_adj_2, n13556, 
            n14826, n14825, n14824, n14823, n14822, n14821, n14820) /* synthesis syn_module_defined=1 */ ;
    output n14672;
    input clk32MHz;
    output n14766;
    output \r_SM_Main_2__N_3262[2] ;
    output [2:0]r_SM_Main;
    input n26029;
    input GND_net;
    output r_Rx_Data;
    input RX_N_2;
    output \r_Bit_Index[0] ;
    output n13551;
    output n4;
    input VCC_net;
    input n15342;
    input n25777;
    output rx_data_ready;
    input n15346;
    output [7:0]rx_data;
    output n18789;
    output n4_adj_1;
    output n4_adj_2;
    output n13556;
    input n14826;
    input n14825;
    input n14824;
    input n14823;
    input n14822;
    input n14821;
    input n14820;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [7:0]n37;
    
    wire n14636;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n14747, n19064, n19265;
    wire [2:0]r_SM_Main_2__N_3268;
    
    wire n1, n3, r_Rx_Data_R, n12, n26054, n26830, n6, n10, 
        n13384, n29299, n19321, n22411, n22410, n22409, n22408, 
        n22407, n22406, n22405;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n14672), 
            .D(n326[2]), .R(n14766));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n14672), 
            .D(n326[1]), .R(n14766));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1125__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n14636), .D(n37[7]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1125__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n14636), .D(n37[6]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1125__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n14636), .D(n37[5]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1125__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n14636), .D(n37[4]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1125__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n14636), .D(n37[3]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1125__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n14636), .D(n37[2]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3262[2] ), 
            .R(n26029));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n19064), .I1(\r_SM_Main_2__N_3262[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n19265));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3268[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n19265), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR r_Clock_Count_1125__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n14636), .D(n37[1]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_2));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1125__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n14636), .D(n37[0]), .R(n14747));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[4]), 
            .I3(r_Clock_Count[1]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i6_4_lut (.I0(r_Clock_Count[3]), .I1(n12), .I2(n26054), .I3(r_Clock_Count[0]), 
            .O(r_SM_Main_2__N_3268[0]));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i21773_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_3268[0]), 
            .I3(GND_net), .O(n26830));
    defparam i21773_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n26830), .I2(\r_SM_Main_2__N_3262[2] ), 
            .I3(r_SM_Main[1]), .O(n14747));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3268[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i25079_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n14636));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i25079_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 i1188_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1188_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(GND_net), .O(n26054));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_833 (.I0(r_Clock_Count[3]), .I1(n26054), .I2(n10), 
            .I3(r_Clock_Count[4]), .O(\r_SM_Main_2__N_3262[2] ));
    defparam i1_4_lut_adj_833.LUT_INIT = 16'heccc;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n19064));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i10961_3_lut (.I0(n14672), .I1(n19064), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n14766));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10961_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3262[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n14672));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1195_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1195_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(\r_SM_Main_2__N_3262[2] ), .O(n13384));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_834 (.I0(\r_Bit_Index[0] ), .I1(n13384), .I2(GND_net), 
            .I3(GND_net), .O(n13551));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_834.LUT_INIT = 16'heeee;
    SB_LUT4 equal_95_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_95_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24492_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3268[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n29299));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i24492_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n29299), .I1(\r_SM_Main_2__N_3262[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n19321));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n19321), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1125_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n22411), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1125_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n22410), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_8 (.CI(n22410), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n22411));
    SB_LUT4 r_Clock_Count_1125_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n22409), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_7 (.CI(n22409), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n22410));
    SB_LUT4 r_Clock_Count_1125_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n22408), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_6 (.CI(n22408), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n22409));
    SB_LUT4 r_Clock_Count_1125_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n22407), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_5 (.CI(n22407), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n22408));
    SB_LUT4 r_Clock_Count_1125_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n22406), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_4 (.CI(n22406), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n22407));
    SB_LUT4 r_Clock_Count_1125_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n22405), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_3 (.CI(n22405), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n22406));
    SB_LUT4 r_Clock_Count_1125_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1125_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1125_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n22405));
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n15342));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n25777));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n15346));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i14996_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n18789));
    defparam i14996_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_91_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_91_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_94_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_94_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_835 (.I0(n13384), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n13556));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_835.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n14826));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n14825));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n14824));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n14823));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n14822));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n14821));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n14820));   // verilog/uart_rx.v(49[10] 144[8])
    
endmodule
