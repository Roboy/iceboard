// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue May 19 19:36:35 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    
    wire n1901, n1899;
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(351[11:24])
    
    wire n28909;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(359[15:20])
    
    wire pwm_setpoint_23__N_207, n209, n211, n39, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, 
        n261, n262, n263, n264, n265, n266, n267, n268, n269, 
        n270, n296, n330, n57890, n334, n335, n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345, n1897, n1895, 
        n356, n379, n22497;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n418, n419, n420, n421, n422, n423, n424, n425, n426, 
        n427, n428, n429, n430, n431, n432, n433, n434, n435, 
        n436, n437, n438, n439, n440, n441;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n69011;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216, n1903, GHA_N_355, GLA_N_372, GHB_N_377, 
        GLB_N_386, GHC_N_391, GLC_N_400, dti_N_404, n29486, n29483, 
        RX_N_2, n1893, n1891, n1889, n1887, n69008, n1885, n1883, 
        n1881;
    wire [31:0]motor_state_23__N_91;
    wire [38:0]encoder1_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
        n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
        n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
        n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
        read_N_409, n51168, n57889, n1405, n25014, n67323, n19, 
        n17, n16, n15, n13, n11, n9, n8, n7, n6, n5, n4, 
        n30, n23, n68684, n68675, n68663, n1828, n1933;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n29480;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [1:0]state;   // verilog/neopixel.v(16[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    
    wire n5076, n5075, n5074, n5073, n5072, n5071, n57979, n5070, 
        n5068, n5067, n5066, n5065, n5064, n5063, n5062, n5061, 
        n5060, n5059, n12, n66094, n68795, n29477, n29474, n29471, 
        n21, n19_adj_5685, n17_adj_5686, n16_adj_5687, n15_adj_5688, 
        n13_adj_5689, n12_adj_5690, n11_adj_5691, n2952, n57966, n57888, 
        n57967;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n57968, n57893, n57965, n57894, n57887, n57886, n3, n4_adj_5692, 
        n5_adj_5693, n6_adj_5694, n7_adj_5695, n8_adj_5696, n9_adj_5697, 
        n10, n11_adj_5698, n12_adj_5699, n13_adj_5700, n14, n15_adj_5701, 
        n16_adj_5702, n17_adj_5703, n18, n19_adj_5704, n20, n21_adj_5705, 
        n22, n23_adj_5706, n24, n25, n2, n57895, n14_adj_5707, 
        n15_adj_5708, n16_adj_5709, n17_adj_5710, n18_adj_5711, n19_adj_5712, 
        n20_adj_5713, n21_adj_5714, n22_adj_5715, n23_adj_5716, n24_adj_5717, 
        n25_adj_5718, n51167, n51116, n29468, n22373, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    
    wire n4_adj_5719;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    
    wire n51115;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    
    wire n57885, \FRAME_MATCHER.rx_data_ready_prev , n57964, n57884, 
        n57978, n2961, n5058, n25004, n29465, n57969, n57883, 
        n29462, n3014, n51166, n51165, n51164, n51163, n51114, 
        n51162, n51161, n51160, n38965, n38922, n38907, n57971, 
        n60939, n1, n60887, n5754, n1130, n6_adj_5720, n1191, 
        n58608, n57882, n57881, n51159, n51100, n1510, n25488, 
        n57880, n2076, n6_adj_5721, n51158, n51157, n14_adj_5722, 
        n13_adj_5723, n57879, n68792, n68789, n68786, n68783, n29459, 
        n62904, n29456, n4894, n4891, n4883, n51113, n51156, n38869, 
        Kp_23__N_869, n38852, n38797, n51112, n38795, n4_adj_5724, 
        n29453, n15_adj_5725, n51155, n29450, n6_adj_5726, n8_adj_5727, 
        n7_adj_5728, n4_adj_5729, n51154, n29447, n29444, n29441, 
        n29438, n25007, n29435, n39313, n29432, n13_adj_5730, n51153, 
        n51099, n66078, \FRAME_MATCHER.i_31__N_2509 , n15_adj_5731, 
        n15_adj_5732, n57975, n39366, n29429, n29426, n29423, n29420, 
        n29417, n29414, n29411, n29408, n29405, n29402, n29399, 
        n29395, n29392, n29389, n29386, n29383, n29380, n29377, 
        n29374, n29371, n29368, n29365, n29362, n29359, n29356, 
        n29353, n29350, n29347, n29344, n29341, n29338, n29335, 
        n29332, n29329, n29326, n29323, n29320, n29317, n29314, 
        n29311, n29308, n29305, n29302, n29299, n29296, n29244, 
        n62, n57977, n29209, n29206, n29205, n29204, n29203, n29202, 
        n29201, n29200, n29199, n29198, n29197, n29194, n29191, 
        n29188, n29187, n29184, n29183, n29182, n29181, n29180, 
        n29179, n29178, n29177, n29176, n29175, n29174, n29173, 
        n29172, n29171, n29170, n29169, n29168, n29165, n29164, 
        n51152, n29160, n29159, n29158, n29157, n29156, n29155, 
        n29123, n29122, n29121, n29120, n29119, n29118, n29117, 
        n29116, n29113, n29110, n29107, n29103, n29102, n29101, 
        n29100, n29099, n29098, n29097, n29096, n29095, n29094, 
        n29093, n29053, n29052, n29051, n29044, n29043, n29040, 
        n29039, n29033, n29032, n29028, n10_adj_5733, n9_adj_5734, 
        n8_adj_5735, n7_adj_5736, n6_adj_5737, n4_adj_5738, n40, n32, 
        n24_adj_5739, n19_adj_5740, n17_adj_5741, n16_adj_5742, n15_adj_5743, 
        n13_adj_5744, n11_adj_5745, n9_adj_5746, n8_adj_5747, n7_adj_5748, 
        n6_adj_5749, n5_adj_5750, n4_adj_5751, n57878, n57877, n57982, 
        n57986, n57876, n57972, n57875, n57874, n4_adj_5752, n4_adj_5753, 
        n6_adj_5754, n5_adj_5755, n6_adj_5756, n5_adj_5757, n57873, 
        n57974, n57872, n57871, n57995, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    wire [23:0]\PID_CONTROLLER.integral_23__N_3715 ;
    
    wire n363, n11_adj_5758;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, position_31__N_3827, n5057, n5056, n5055, n5054, 
        n5053, n5052, n5051, n5050, n5049, n5048, n5047;
    wire [1:0]a_new_adj_5905;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5760, n25237, position_31__N_3827_adj_5761, n68993, 
        n29951, n26, n25_adj_5762, n24_adj_5763, n23_adj_5764, n4_adj_5765, 
        n3_adj_5766;
    wire [7:0]data_adj_5918;   // verilog/eeprom.v(23[12:16])
    
    wire ready_prev, rw;
    wire [7:0]state_adj_5919;   // verilog/eeprom.v(27[11:16])
    wire [7:0]state_7__N_3916;
    
    wire n24_adj_5769, n29948, n68774, n29945, n29942, n5093, n5091, 
        n5090, n5089, n5088, n57870, n2_adj_5770, n29920, n29919, 
        n29918, n29917, n29916, n29915, n29914, n29912, n29911, 
        n29910, n29909, n29908, n29907, n29906, n29904, n29903, 
        n29902, n29901, n29900, n29899, n29898, n29897, n29896, 
        n29895, n5087;
    wire [15:0]data_adj_5926;   // verilog/tli4970.v(27[14:18])
    
    wire n57970, n29894, n29893, n29892, n66060, n57869, n57868, 
        n57867, n53988, n5086, n5085, n5084, n5083, n5082, n5081, 
        n5080, n5079, n5078, n5077, state_7__N_4317, n51151, n66058, 
        n29024, n29023, n22_adj_5779, n21_adj_5780, n29020, n29018, 
        n29017, n29016, n6579, n57866, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n57865, n57990;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n68768, n68762, n68756, n20_adj_5781, n19_adj_5782, n18_adj_5783, 
        n17_adj_5784, n16_adj_5785;
    wire [2:0]r_SM_Main_adj_5939;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5940;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_5941;   // verilog/uart_tx.v(34[16:27])
    
    wire n14_adj_5797, n22362, n29778, n29777, n29776, n29775, n29774, 
        n29773, n29772, n15_adj_5798, n29771, n14_adj_5799, n13_adj_5800, 
        n12_adj_5801, n11_adj_5802, n29770, n29769, n29768, n29767, 
        n29765, n29763, n29762, n29761, n29760, n29759, n29758, 
        n29757, n29756, n29755, n29754, n57864, n29753, n29752;
    wire [7:0]state_adj_5949;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire enable_slow_N_4211, n29751, n29750, n29749, n10_adj_5804, 
        n9_adj_5805, n8_adj_5806, n7_adj_5807, n29748, n6_adj_5808, 
        n5_adj_5809, n29747, n29745, n29744, n29743, n29742;
    wire [7:0]state_7__N_4108;
    
    wire n29740, n29739, n29738, n5_adj_5810, n29737, n29736, n29735, 
        n25136, n6388;
    wire [7:0]state_7__N_4124;
    
    wire n57863, n10_adj_5811, n29704, n29013, n29009, n62903, n57356, 
        n60747, n57862, n29683, n57861, n57860, n57994, n60858, 
        n27429, n57859, n57892, n57989, n57961, n57988, n57858, 
        n51486, n57857, n57987, n28782, n29667, n57963, n57856, 
        n28780, n57996, n66054, n35, n68990, n57855, n57891, n57854, 
        n57998, n57853, n51485, n57852, n57984, n57851, n29663, 
        n57850, n57983, n57849, n57901, n28772, n57897, n57848, 
        n57847, n57981, n28768, n28767, n51484, n68229, n13051, 
        n51483, n51482, n51481, n51480, n13052, n51150, n51479, 
        n51149, n51478, n51477, n51476, n51148, n51147, n51475, 
        n51474, n51473, n57846, n51472, n51471, n51470, n51469, 
        n13053, n51468, n51467, n51466, n51465, n51464, n51463, 
        n51462, n51461, n51460, n62052, n51459, n57558, n51111, 
        n51146, n51145, n51458, n51457, n51456, n51455, n24_adj_5812, 
        n51454, n51453, n20_adj_5813, n51452, n21_adj_5814, n51451, 
        n51450, n57845, n20_adj_5815, n19_adj_5816, n25141, n51449, 
        n51448, n51447, n51446, n13054, n51445, n51444, n10_adj_5817, 
        n51443, n51442, n51441, n51440, n17_adj_5818, n16_adj_5819, 
        n13055, n29000, n58000, n51439, n28969, n51438, n51437, 
        n51110, n51144, n51098, n51436, n51435, n51434, n51433, 
        n13056, n51432, n51431, n51990, n51430, n51429, n51989, 
        n51988, n51987, n25112, n51986, n51985, n51984, n28764, 
        n57844, n25148, n57980, n51143, n51142, n51141, n9941, 
        n9942, n9943, n9946, n9945, n9944, n68741, n9936, n9937, 
        n9938, n9940, n9939, n9931, n9932, n25145, n9935, n9934, 
        n9933, n9928, n25151, n51406, n51405, n9930, n9929, n51404, 
        n51403, n51402, n51401, n68738, n51400, n51399, n51398, 
        n51397, n51396, n9927, n51395, n51394, n26180, n51140, 
        n51393, n51109, n51392, n51097, n51139, n51391, n51390, 
        n51389, n51388, n51387, n51386, n51385, n51384, n51383, 
        n51138, n51137, n51136, n51382, n51381, n51380, n57973, 
        n25996, n51379, n51378, n51377, n51096, n57843, n57842, 
        n57999, n51376, n51375, n51374, n51373, n4_adj_5820, n6_adj_5821, 
        n8_adj_5822, n9_adj_5823, n11_adj_5824, n13_adj_5825, n15_adj_5826, 
        n25269, n51372, n4_adj_5827, n6_adj_5828, n8_adj_5829, n9_adj_5830, 
        n68179, n51371, n111, n57985, n57841, n51135, n51370, 
        n27295, n51369, n27292, n51368, n51134, n29653, n27288, 
        n51367, n51366, n51365, n51364, n51363, n48, n49, n50, 
        n51, n52, n53, n54, n55, n51362, n51361, n27270, n57997, 
        n51360, n27262, n51359, n51133, n51132, n51358, n9618, 
        n51357, n29647, n57840, n57839, n27211, n57992, n57838, 
        n57837, n57836, n57993, n57900, n57962, n28927, n57835, 
        n58004, n58003, n58002, n58001, n57960, n57959, n57958, 
        n57957, n57956, n58022, n57955, n57954, n57953, n57952, 
        n57951, n57950, n57949, n57948, n57947, n57946, n57945, 
        n57944, n57943, n57942, n57941, n57940, n57939, n57938, 
        n57937, n57936, n58321, n57935, n57934, n57933, n57932, 
        n57931, n57930, n58245, n57929, n57928, n57927, n57926, 
        n57925, n57924, n57923, n57922, n57921, n57920, n57919, 
        n57918, n68924, n57917, n57916, n57915, n57914, n57913, 
        n57899, n57912, n57911, n57910, n57898, n28838, n28837, 
        n57909, n57908, n57907, n57905, n28671, n57906, n28831, 
        n57834, n57904, n57903, n28827, n57902, n28825, n28009, 
        n28002, n27997, n27994, n58145, n58144, n58143, n58142, 
        n58141, n27972, n27968, n28417, n27924, n27920, n57991, 
        n51356, n51355, n51354, n51353, n57896, n51352, n51351, 
        n27187, n51108, n51350, n25117, n51349, n51348, n62902, 
        n68726, n68720, n68714, n68702, n68699, n57286, n57370, 
        n57628, n51107, n51106, n67678, n51131, n13040, n54370, 
        n13038, n13039, n68645, n68642, n68639, n68633, n68624, 
        n68969, n68966, n68963, n13043, n51130, n13042, n13041, 
        n51105, n29608, n29605, n29602, n29599, n25119, n13045, 
        n51129, n13044, n29593, n51128, n51095, n13046, n13048, 
        n38, n13047, n57372, n57374, n28993, n57376, n13049, n57378, 
        n57380, n29516, n13050, n28987, n29510, n29507, n29504, 
        n28982, n28979, n28976, n29501, n29498, n29495, n14_adj_5831, 
        n51104, n10_adj_5832, n51127, n68960, n57976, n51126, n51125, 
        n68303, n68302, n68289, n68288, n66692, n51124, n51103, 
        n10_adj_5833, n53279, n38105, n53_adj_5834, n62_adj_5835, 
        n51123, n6_adj_5836, n51102, n51122, n68948, n58436, n68942, 
        n24998, n51101, n51121, n38106, n68936, n53121, n51120, 
        n53862, n51119, n68180, n68930, n58238, n51118, n57833, 
        n68918, n51094, n58312, n51093, n27600, n7_adj_5837, n25133, 
        n25130, n7_adj_5838, n7_adj_5839, n66612, n28972, n51117, 
        n68104, n68098, n68094, n68083, n68082, n66592, n68064, 
        n68912, n68043, n58970, n58968, n29, n27, n23_adj_5840, 
        n67870, n67869, n10_adj_5841, n67860, n67859, n68906, n67792, 
        n67791, n6_adj_5842, n61676, n68900, n14_adj_5843, n26_adj_5844, 
        n13_adj_5845, n61658, n67427, n66451, n68894, n6_adj_5846, 
        n61640, n61622, n15_adj_5847, n14_adj_5848, n66958, n66400, 
        n61604, n4_adj_5849, n66388, n62649, n68888, n7_adj_5850, 
        n17_adj_5851, n25_adj_5852, n56586, n24_adj_5853, n61586, 
        n61568, n66342, n68882, n56676, n66333, n61550, n59879, 
        n59877, n67429, n68876, n67431, n67433, n15_adj_5854, n58185, 
        n62531, n14_adj_5855, n68870, n58276, n58264, n58653, n58446, 
        n58225, n58363, n59845, n59843, n58742, n60510, n65592, 
        n67952, n5_adj_5856, n57832, n65590, n59823, n59821, n65575, 
        n68864, n58707, n58698, n65569, n65562, n58147, n58748, 
        n60892, n69042, n25_adj_5857, n68861, n65556, n60645, n65553, 
        n65551, n65548, n58819, n58777, n67561, n65537, n58867, 
        n58857, n58845, n58835, n58828, n65536, n65535, n65534, 
        n65533, n65532, n65531, n58096, n62535, n65488, n68228, 
        n68855, n65475, n65474, n67563, n65449, n61280, n61278, 
        n58644, n57342, n12_adj_5858, n57346, n57350, n57354, n4_adj_5859, 
        n8_adj_5860, n58632, n69032, n7_adj_5861, n58952, n68849, 
        n57504, n7_adj_5862, n69026, n12_adj_5863, n11_adj_5864, n67180, 
        n69020, n62677, n60966, n23_adj_5865, n65385, n58140, n58680, 
        n4_adj_5866, n58922, n58139, n58391, n58919, n68604, n65376, 
        n57676, n58925, n6_adj_5867, n6_adj_5868, n6_adj_5869, n65364;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dir_189 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 n9618_bdd_4_lut_51826 (.I0(n9618), .I1(n428), .I2(current[15]), 
            .I3(duty[23]), .O(n68888));
    defparam n9618_bdd_4_lut_51826.LUT_INIT = 16'he4aa;
    SB_DFFE dti_191 (.Q(dti), .C(clk16MHz), .E(n27187), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i14008_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n22362), .I3(GND_net), .O(n29751));   // verilog/coms.v(130[12] 305[6])
    defparam i14008_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13352_3_lut (.I0(current[9]), .I1(data_adj_5926[9]), .I2(n27270), 
            .I3(GND_net), .O(n29095));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13352_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13353_3_lut (.I0(current[8]), .I1(data_adj_5926[8]), .I2(n27270), 
            .I3(GND_net), .O(n29096));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13353_3_lut.LUT_INIT = 16'hcaca;
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4124[3])) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n51348), .I0(GND_net), 
            .I1(n24_adj_5763), .CO(n51349));
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_5762), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.GND_net(GND_net), .clk16MHz(clk16MHz), 
            .n111(n111), .state({state}), .neopxl_color({neopxl_color}), 
            .\bit_ctr[1] (bit_ctr[1]), .\bit_ctr[0] (bit_ctr[0]), .n29244(n29244), 
            .VCC_net(VCC_net), .n5(n5_adj_5856), .n25(n25_adj_5857), .timer({timer}), 
            .n29205(n29205), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n29204(n29204), .n29203(n29203), .n27429(n27429), .n29202(n29202), 
            .n29201(n29201), .n29200(n29200), .n29199(n29199), .n29198(n29198), 
            .n29197(n29197), .n29187(n29187), .n29043(n29043), .NEOPXL_c(NEOPXL_c), 
            .n23(n23_adj_5865), .n39366(n39366), .LED_c(LED_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_5762), .CO(n51348));
    SB_LUT4 i14009_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n22362), .I3(GND_net), .O(n29752));   // verilog/coms.v(130[12] 305[6])
    defparam i14009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(n4883), .I1(GND_net), .I2(n15_adj_5701), 
            .I3(n51154), .O(n5061)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_12 (.CI(n51154), .I0(GND_net), .I1(n15_adj_5701), 
            .CO(n51155));
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(n4883), .I1(GND_net), .I2(n16_adj_5702), 
            .I3(n51153), .O(n5062)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n51153), .I0(GND_net), .I1(n16_adj_5702), 
            .CO(n51154));
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(n4883), .I1(GND_net), .I2(n17_adj_5703), 
            .I3(n51152), .O(n5063)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n51152), .I0(GND_net), .I1(n17_adj_5703), 
            .CO(n51153));
    SB_LUT4 i14010_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n22362), .I3(GND_net), .O(n29753));   // verilog/coms.v(130[12] 305[6])
    defparam i14010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13354_3_lut (.I0(current[7]), .I1(data_adj_5926[7]), .I2(n27270), 
            .I3(GND_net), .O(n29097));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(n4883), .I1(GND_net), .I2(n18), 
            .I3(n51151), .O(n5064)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n51151), .I0(GND_net), .I1(n18), 
            .CO(n51152));
    SB_LUT4 i13355_3_lut (.I0(current[6]), .I1(data_adj_5926[6]), .I2(n27270), 
            .I3(GND_net), .O(n29098));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14011_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n22362), .I3(GND_net), .O(n29754));   // verilog/coms.v(130[12] 305[6])
    defparam i14011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13356_3_lut (.I0(current[5]), .I1(data_adj_5926[5]), .I2(n27270), 
            .I3(GND_net), .O(n29099));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13357_3_lut (.I0(current[4]), .I1(data_adj_5926[4]), .I2(n27270), 
            .I3(GND_net), .O(n29100));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(n4883), .I1(GND_net), .I2(n19_adj_5704), 
            .I3(n51150), .O(n5065)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n51150), .I0(GND_net), .I1(n19_adj_5704), 
            .CO(n51151));
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(n4883), .I1(GND_net), .I2(n20), 
            .I3(n51149), .O(n5066)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_157_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n51129), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_7 (.CI(n51149), .I0(GND_net), .I1(n20), 
            .CO(n51150));
    SB_CARRY add_157_18 (.CI(n51129), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n51130));
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(n4883), .I1(GND_net), .I2(n21_adj_5705), 
            .I3(n51148), .O(n5067)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n68888_bdd_4_lut (.I0(n68888), .I1(duty[13]), .I2(n257), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[13]));
    defparam n68888_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY unary_minus_21_add_3_6 (.CI(n51148), .I0(GND_net), .I1(n21_adj_5705), 
            .CO(n51149));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(n296), .I1(GND_net), .I2(n22), 
            .I3(n51147), .O(n5068)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_238_13_lut (.I0(current[11]), .I1(duty[14]), .I2(n68604), 
            .I3(n51103), .O(n259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_13_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_157_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n51128), .O(n1310)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13358_3_lut (.I0(current[3]), .I1(data_adj_5926[3]), .I2(n27270), 
            .I3(GND_net), .O(n29101));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13358_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n51147), .I0(GND_net), .I1(n22), 
            .CO(n51148));
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(n379), .I1(GND_net), .I2(n23_adj_5706), 
            .I3(n51146), .O(n4_adj_5849)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_238_5_lut (.I0(current[3]), .I1(duty[6]), .I2(n68604), 
            .I3(n51095), .O(n267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58264));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_21_add_3_4 (.CI(n51146), .I0(GND_net), .I1(n23_adj_5706), 
            .CO(n51147));
    SB_CARRY add_238_13 (.CI(n51103), .I0(duty[14]), .I1(n68604), .CO(n51104));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n51145), .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n51145), .I0(GND_net), .I1(n24), 
            .CO(n51146));
    SB_CARRY add_157_17 (.CI(n51128), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n51129));
    SB_LUT4 add_157_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n51127), .O(n1311)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_16 (.CI(n51127), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n51128));
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[1] [4]), .I1(n25488), .I2(\data_in_frame[2] [0]), 
            .I3(n58264), .O(n10_adj_5817));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[1] [7]), .I1(n10_adj_5817), .I2(\data_in_frame[4] [1]), 
            .I3(GND_net), .O(Kp_23__N_869));   // verilog/coms.v(99[12:25])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14012_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n22362), .I3(GND_net), .O(n29755));   // verilog/coms.v(130[12] 305[6])
    defparam i14012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14013_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n22373), .I3(GND_net), .O(n29756));   // verilog/coms.v(130[12] 305[6])
    defparam i14013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13359_3_lut (.I0(current[2]), .I1(data_adj_5926[2]), .I2(n27270), 
            .I3(GND_net), .O(n29102));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13360_3_lut (.I0(current[1]), .I1(data_adj_5926[1]), .I2(n27270), 
            .I3(GND_net), .O(n29103));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19101_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n22373), .I3(GND_net), .O(n29757));
    defparam i19101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19121_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n22373), .I3(GND_net), .O(n29758));
    defparam i19121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n4_adj_5849), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(n65376)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i19128_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n22373), .I3(GND_net), .O(n29759));
    defparam i19128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13373_3_lut (.I0(baudrate[31]), .I1(data_adj_5918[7]), .I2(n60892), 
            .I3(GND_net), .O(n29116));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13373_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n51145));
    SB_LUT4 add_157_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n51144), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n51143), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_32 (.CI(n51143), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n51144));
    SB_LUT4 add_157_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n51142), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_31 (.CI(n51142), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n51143));
    SB_LUT4 i14017_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n22373), .I3(GND_net), .O(n29760));   // verilog/coms.v(130[12] 305[6])
    defparam i14017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_157_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n51141), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_30 (.CI(n51141), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n51142));
    SB_LUT4 add_157_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n51140), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_29 (.CI(n51140), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n51141));
    SB_LUT4 i14018_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n22373), .I3(GND_net), .O(n29761));   // verilog/coms.v(130[12] 305[6])
    defparam i14018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13374_3_lut (.I0(baudrate[30]), .I1(data_adj_5918[6]), .I2(n60892), 
            .I3(GND_net), .O(n29117));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13375_3_lut (.I0(baudrate[29]), .I1(data_adj_5918[5]), .I2(n60892), 
            .I3(GND_net), .O(n29118));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14019_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n22373), .I3(GND_net), .O(n29762));   // verilog/coms.v(130[12] 305[6])
    defparam i14019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13376_3_lut (.I0(baudrate[28]), .I1(data_adj_5918[4]), .I2(n60892), 
            .I3(GND_net), .O(n29119));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_157_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n51139), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14020_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n22373), .I3(GND_net), .O(n29763));   // verilog/coms.v(130[12] 305[6])
    defparam i14020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13377_3_lut (.I0(baudrate[27]), .I1(data_adj_5918[3]), .I2(n60892), 
            .I3(GND_net), .O(n29120));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_238_12_lut (.I0(current[10]), .I1(duty[13]), .I2(n68604), 
            .I3(n51102), .O(n260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_12_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i14022_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n22373), .I3(GND_net), .O(n29765));   // verilog/coms.v(130[12] 305[6])
    defparam i14022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13378_3_lut (.I0(baudrate[26]), .I1(data_adj_5918[2]), .I2(n60892), 
            .I3(GND_net), .O(n29121));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13379_3_lut (.I0(baudrate[25]), .I1(data_adj_5918[1]), .I2(n60892), 
            .I3(GND_net), .O(n29122));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_4_lut (.I0(n53862), .I1(n58363), .I2(n58391), .I3(n58698), 
            .O(n12_adj_5863));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14024_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n22373), .I3(GND_net), .O(n29767));   // verilog/coms.v(130[12] 305[6])
    defparam i14024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13380_3_lut (.I0(baudrate[24]), .I1(data_adj_5918[0]), .I2(n60892), 
            .I3(GND_net), .O(n29123));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14025_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n22373), .I3(GND_net), .O(n29768));   // verilog/coms.v(130[12] 305[6])
    defparam i14025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14026_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n22373), .I3(GND_net), .O(n29769));   // verilog/coms.v(130[12] 305[6])
    defparam i14026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14027_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n22373), .I3(GND_net), .O(n29770));   // verilog/coms.v(130[12] 305[6])
    defparam i14027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14028_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n22373), .I3(GND_net), .O(n29771));   // verilog/coms.v(130[12] 305[6])
    defparam i14028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14029_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n22373), .I3(GND_net), .O(n29772));   // verilog/coms.v(130[12] 305[6])
    defparam i14029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19067_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n22373), .I3(GND_net), .O(n29773));
    defparam i19067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14031_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n22373), .I3(GND_net), .O(n29774));   // verilog/coms.v(130[12] 305[6])
    defparam i14031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14032_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n22373), .I3(GND_net), .O(n29775));   // verilog/coms.v(130[12] 305[6])
    defparam i14032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14033_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n22373), .I3(GND_net), .O(n29776));   // verilog/coms.v(130[12] 305[6])
    defparam i14033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14034_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n22373), .I3(GND_net), .O(n29777));   // verilog/coms.v(130[12] 305[6])
    defparam i14034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14035_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n22373), .I3(GND_net), .O(n29778));   // verilog/coms.v(130[12] 305[6])
    defparam i14035_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_157_28 (.CI(n51139), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n51140));
    SB_LUT4 add_157_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n51126), .O(n1312)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_238_5 (.CI(n51095), .I0(duty[6]), .I1(n68604), .CO(n51096));
    SB_LUT4 add_157_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n51138), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_27 (.CI(n51138), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n51139));
    SB_CARRY add_238_12 (.CI(n51102), .I0(duty[13]), .I1(n68604), .CO(n51103));
    SB_LUT4 add_157_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n51137), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_15 (.CI(n51126), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n51127));
    SB_CARRY add_157_26 (.CI(n51137), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n51138));
    SB_LUT4 add_157_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n51125), .O(n1313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n51136), .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_25 (.CI(n51136), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n51137));
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51891 (.I0(byte_transmit_counter[3]), 
            .I1(n67433), .I2(n65553), .I3(byte_transmit_counter[4]), .O(n68882));
    defparam byte_transmit_counter_3__bdd_4_lut_51891.LUT_INIT = 16'he4aa;
    SB_LUT4 n68882_bdd_4_lut (.I0(n68882), .I1(n68861), .I2(n7_adj_5839), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n68882_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_157_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n51135), .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_14 (.CI(n51125), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n51126));
    SB_LUT4 add_157_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n51124), .O(n1314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_24 (.CI(n51135), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n51136));
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 LessThan_1069_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5828));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1069_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51816 (.I0(byte_transmit_counter[3]), 
            .I1(n67431), .I2(n65562), .I3(byte_transmit_counter[4]), .O(n68876));
    defparam byte_transmit_counter_3__bdd_4_lut_51816.LUT_INIT = 16'he4aa;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n68876_bdd_4_lut (.I0(n68876), .I1(n68855), .I2(n7_adj_5838), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n68876_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49038_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n66054));   // verilog/uart_rx.v(119[17:57])
    defparam i49038_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i23369_2_lut_2_lut (.I0(n296), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n5047));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i23369_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_157_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n51134), .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY add_157_23 (.CI(n51134), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n51135));
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 add_157_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n51133), .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_22 (.CI(n51133), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n51134));
    SB_LUT4 i13692_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n60939), .I3(GND_net), .O(n29435));   // verilog/coms.v(130[12] 305[6])
    defparam i13692_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_157_13 (.CI(n51124), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n51125));
    SB_LUT4 add_157_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n51132), .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_21 (.CI(n51132), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n51133));
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51811 (.I0(byte_transmit_counter[3]), 
            .I1(n67429), .I2(n65590), .I3(byte_transmit_counter[4]), .O(n68870));
    defparam byte_transmit_counter_3__bdd_4_lut_51811.LUT_INIT = 16'he4aa;
    SB_LUT4 n9618_bdd_4_lut_51856 (.I0(n9618), .I1(n422), .I2(current[15]), 
            .I3(duty[23]), .O(n68924));
    defparam n9618_bdd_4_lut_51856.LUT_INIT = 16'he4aa;
    SB_LUT4 i48845_2_lut (.I0(n68663), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65562));
    defparam i48845_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_157_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n51131), .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_157_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n51123), .O(n1315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_20 (.CI(n51131), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n51132));
    SB_LUT4 i50415_3_lut (.I0(n68993), .I1(n68741), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67431));
    defparam i50415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_157_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n51130), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n68924_bdd_4_lut (.I0(n68924), .I1(duty[19]), .I2(n251), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[19]));
    defparam n68924_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_238_11_lut (.I0(current[9]), .I1(duty[12]), .I2(n68604), 
            .I3(n51101), .O(n261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_11_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_157_12 (.CI(n51123), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n51124));
    SB_LUT4 i13412_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .I2(control_update), .I3(GND_net), .O(n29155));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n68870_bdd_4_lut (.I0(n68870), .I1(n68639), .I2(n68849), .I3(byte_transmit_counter[4]), 
            .O(tx_data[3]));
    defparam n68870_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_157_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n51122), .O(n1316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49062_3_lut_4_lut (.I0(r_Clock_Count_adj_5940[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5940[2]), .O(n66078));   // verilog/uart_tx.v(117[17:57])
    defparam i49062_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_238_4_lut (.I0(current[2]), .I1(duty[5]), .I2(n68604), 
            .I3(n51094), .O(n268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i13413_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I2(control_update), .I3(GND_net), .O(n29156));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13413_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_238_11 (.CI(n51101), .I0(duty[12]), .I1(n68604), .CO(n51102));
    SB_CARRY add_157_11 (.CI(n51122), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n51123));
    SB_LUT4 i13414_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .I2(control_update), .I3(GND_net), .O(n29157));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13415_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I2(control_update), .I3(GND_net), .O(n29158));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13415_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13416_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(control_update), .I3(GND_net), .O(n29159));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1072_i13_2_lut (.I0(r_Clock_Count_adj_5940[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5825));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13417_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I2(control_update), .I3(GND_net), .O(n29160));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51806 (.I0(byte_transmit_counter[3]), 
            .I1(n67427), .I2(n65592), .I3(byte_transmit_counter[4]), .O(n68864));
    defparam byte_transmit_counter_3__bdd_4_lut_51806.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_1072_i15_2_lut (.I0(r_Clock_Count_adj_5940[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5826));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1072_i9_2_lut (.I0(r_Clock_Count_adj_5940[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5823));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n68864_bdd_4_lut (.I0(n68864), .I1(n68675), .I2(n7_adj_5837), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n68864_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_1072_i11_2_lut (.I0(r_Clock_Count_adj_5940[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5824));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i11_2_lut.LUT_INIT = 16'h6666;
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 LessThan_1072_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5940[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5821));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i13421_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(control_update), .I3(GND_net), .O(n29164));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13421_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 LessThan_1072_i4_4_lut (.I0(r_Clock_Count_adj_5940[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5940[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5820));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i13425_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(control_update), .I3(GND_net), .O(n29168));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50775_3_lut (.I0(n4_adj_5820), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5824), 
            .I3(GND_net), .O(n67791));   // verilog/uart_tx.v(117[17:57])
    defparam i50775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50776_3_lut (.I0(n67791), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5825), 
            .I3(GND_net), .O(n67792));   // verilog/uart_tx.v(117[17:57])
    defparam i50776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49942_4_lut (.I0(n13_adj_5825), .I1(n11_adj_5824), .I2(n9_adj_5823), 
            .I3(n66078), .O(n66958));
    defparam i49942_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1072_i8_3_lut (.I0(n6_adj_5821), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5823), .I3(GND_net), .O(n8_adj_5822));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1072_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49676_3_lut (.I0(n67792), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5826), 
            .I3(GND_net), .O(n66692));   // verilog/uart_tx.v(117[17:57])
    defparam i49676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50662_4_lut (.I0(n66692), .I1(n8_adj_5822), .I2(n15_adj_5826), 
            .I3(n66958), .O(n67678));   // verilog/uart_tx.v(117[17:57])
    defparam i50662_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50663_3_lut (.I0(n67678), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5940[8]), 
            .I3(GND_net), .O(n4894));   // verilog/uart_tx.v(117[17:57])
    defparam i50663_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13426_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(control_update), .I3(GND_net), .O(n29169));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13427_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(control_update), .I3(GND_net), .O(n29170));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_157_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n51121), .O(n1317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13428_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(control_update), .I3(GND_net), .O(n29171));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13428_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13429_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(control_update), .I3(GND_net), .O(n29172));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13429_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_157_10 (.CI(n51121), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n51122));
    SB_LUT4 add_157_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n51120), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1062_1_lut (.I0(n296), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n4883));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1062_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5701));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1069_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5830));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1069_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1069_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5827));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1069_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 n9618_bdd_4_lut_51831 (.I0(n9618), .I1(n427), .I2(current[15]), 
            .I3(duty[23]), .O(n68894));
    defparam n9618_bdd_4_lut_51831.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_1069_i8_3_lut (.I0(n6_adj_5828), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5830), .I3(GND_net), .O(n8_adj_5829));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1069_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51163_4_lut (.I0(n8_adj_5829), .I1(n4_adj_5827), .I2(n9_adj_5830), 
            .I3(n66054), .O(n68179));   // verilog/uart_rx.v(119[17:57])
    defparam i51163_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51164_3_lut (.I0(n68179), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n68180));   // verilog/uart_rx.v(119[17:57])
    defparam i51164_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51027_3_lut (.I0(n68180), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n68043));   // verilog/uart_rx.v(119[17:57])
    defparam i51027_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49680_3_lut (.I0(n68043), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4891));   // verilog/uart_rx.v(119[17:57])
    defparam i49680_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13257_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n7_adj_5861), 
            .I3(GND_net), .O(n29000));   // verilog/coms.v(130[12] 305[6])
    defparam i13257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13430_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(control_update), .I3(GND_net), .O(n29173));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13250_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n7_adj_5861), 
            .I3(GND_net), .O(n28993));   // verilog/coms.v(130[12] 305[6])
    defparam i13250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13431_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(control_update), .I3(GND_net), .O(n29174));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13431_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_157_9 (.CI(n51120), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n51121));
    SB_LUT4 add_157_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n51119), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13432_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(control_update), .I3(GND_net), .O(n29175));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13432_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i13433_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(control_update), .I3(GND_net), .O(n29176));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13434_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(control_update), .I3(GND_net), .O(n29177));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49146_4_lut (.I0(data_ready), .I1(n6579), .I2(n24_adj_5853), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n65548));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49146_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i49290_2_lut (.I0(n24_adj_5853), .I1(n6579), .I2(GND_net), 
            .I3(GND_net), .O(n65551));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49290_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13435_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(control_update), .I3(GND_net), .O(n29178));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49_4_lut (.I0(n65551), .I1(n65548), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5842), .O(n56586));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i13961_3_lut (.I0(\data_in_frame[23] [7]), .I1(rx_data[7]), 
            .I2(n28009), .I3(GND_net), .O(n29704));   // verilog/coms.v(130[12] 305[6])
    defparam i13961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[23] [6]), .I1(n27924), .I2(n28009), 
            .I3(rx_data[6]), .O(n57346));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13436_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(control_update), .I3(GND_net), .O(n29179));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13437_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(control_update), .I3(GND_net), .O(n29180));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1785 (.I0(\data_in_frame[23] [2]), .I1(n27924), 
            .I2(n28009), .I3(rx_data[2]), .O(n57350));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1785.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13438_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(control_update), .I3(GND_net), .O(n29181));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1786 (.I0(\data_in_frame[23] [1]), .I1(n27924), 
            .I2(n28009), .I3(rx_data[1]), .O(n57354));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1786.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13439_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(control_update), .I3(GND_net), .O(n29182));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13440_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(control_update), .I3(GND_net), .O(n29183));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1787 (.I0(\data_in_frame[23] [0]), .I1(n27924), 
            .I2(n28009), .I3(rx_data[0]), .O(n57356));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1787.LUT_INIT = 16'h3a0a;
    SB_CARRY add_157_8 (.CI(n51119), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n51120));
    SB_LUT4 add_157_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n51118), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9618_bdd_4_lut_51841 (.I0(n9618), .I1(n425), .I2(current[15]), 
            .I3(duty[23]), .O(n68906));
    defparam n9618_bdd_4_lut_51841.LUT_INIT = 16'he4aa;
    SB_LUT4 n68906_bdd_4_lut (.I0(n68906), .I1(duty[16]), .I2(n254), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[16]));
    defparam n68906_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51836 (.I0(n9618), .I1(n426), .I2(current[15]), 
            .I3(duty[23]), .O(n68900));
    defparam n9618_bdd_4_lut_51836.LUT_INIT = 16'he4aa;
    SB_LUT4 n68894_bdd_4_lut (.I0(n68894), .I1(duty[14]), .I2(n256), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[14]));
    defparam n68894_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13444_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29187));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13444_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_157_7 (.CI(n51118), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n51119));
    SB_LUT4 i13454_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29197));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13455_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29198));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13456_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29199));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13920_4_lut (.I0(n61280), .I1(r_Bit_Index[0]), .I2(n58970), 
            .I3(n27292), .O(n29663));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13920_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i13457_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29200));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_157_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n51117), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13458_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29201));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13458_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13459_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29202));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13459_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13910_4_lut (.I0(n61278), .I1(r_Bit_Index_adj_5941[0]), .I2(n58968), 
            .I3(n27295), .O(n29653));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13910_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i51394_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n38797), .I3(GND_net), .O(n27262));
    defparam i51394_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i48638_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n65449));
    defparam i48638_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5851));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_CARRY add_157_6 (.CI(n51117), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n51118));
    SB_LUT4 i13244_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n7_adj_5861), 
            .I3(GND_net), .O(n28987));   // verilog/coms.v(130[12] 305[6])
    defparam i13244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5729));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /media/letrend/icecube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n9618_bdd_4_lut (.I0(n9618), .I1(n439), .I2(current[2]), .I3(duty[23]), 
            .O(n69032));
    defparam n9618_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69032_bdd_4_lut (.I0(n69032), .I1(duty[2]), .I2(n268), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n69032_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51941 (.I0(n9618), .I1(n440), .I2(current[1]), 
            .I3(duty[23]), .O(n69026));
    defparam n9618_bdd_4_lut_51941.LUT_INIT = 16'he4aa;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 n9618_bdd_4_lut_51851 (.I0(n9618), .I1(n423), .I2(current[15]), 
            .I3(duty[23]), .O(n68918));
    defparam n9618_bdd_4_lut_51851.LUT_INIT = 16'he4aa;
    SB_LUT4 n69026_bdd_4_lut (.I0(n69026), .I1(duty[1]), .I2(n269), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n69026_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51747 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(byte_transmit_counter[1]), .O(n68792));
    defparam byte_transmit_counter_0__bdd_4_lut_51747.LUT_INIT = 16'he4aa;
    SB_LUT4 i23261_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n38797), .I3(GND_net), .O(n38907));
    defparam i23261_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 n68792_bdd_4_lut (.I0(n68792), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(byte_transmit_counter[1]), 
            .O(n68795));
    defparam n68792_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1788 (.I0(state_adj_5919[2]), .I1(state_adj_5919[1]), 
            .I2(state_adj_5919[0]), .I3(n38869), .O(n57286));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'ha8e8;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i14149_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[1]), .I2(n6_adj_5726), 
            .I3(n25148), .O(n29892));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14149_4_lut.LUT_INIT = 16'hccca;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i14150_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[2]), .I2(n6_adj_5726), 
            .I3(n25145), .O(n29893));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14150_4_lut.LUT_INIT = 16'hccca;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i13460_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29203));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13460_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i13461_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29204));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13461_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i2_2_lut (.I0(dti_counter[7]), .I1(dti_counter[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5867));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1789 (.I0(dti_counter[0]), .I1(dti_counter[3]), 
            .I2(n6_adj_5867), .I3(dti_counter[1]), .O(n6_adj_5868));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i14151_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[3]), .I2(n6_adj_5726), 
            .I3(n25112), .O(n29894));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14151_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4_4_lut_adj_1790 (.I0(dti_counter[2]), .I1(dti_counter[6]), 
            .I2(dti_counter[4]), .I3(n6_adj_5868), .O(n22497));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i4_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_DFF dti_counter_1929__i0 (.Q(dti_counter[0]), .C(clk16MHz), .D(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i14152_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[4]), .I2(n6_adj_5756), 
            .I3(n25151), .O(n29895));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14152_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51742 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n68786));
    defparam byte_transmit_counter_0__bdd_4_lut_51742.LUT_INIT = 16'he4aa;
    SB_LUT4 i14153_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[5]), .I2(n6_adj_5756), 
            .I3(n25148), .O(n29896));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14153_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n68786_bdd_4_lut (.I0(n68786), .I1(\data_out_frame[21] [3]), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n68789));
    defparam n68786_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51561_2_lut (.I0(n22497), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i51561_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i13462_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29205));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9618_bdd_4_lut_51821 (.I0(n9618), .I1(n429), .I2(current[15]), 
            .I3(duty[23]), .O(n68774));
    defparam n9618_bdd_4_lut_51821.LUT_INIT = 16'he4aa;
    SB_LUT4 n68774_bdd_4_lut (.I0(n68774), .I1(duty[12]), .I2(n258), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[12]));
    defparam n68774_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51727 (.I0(n9618), .I1(n430), .I2(current[11]), 
            .I3(duty[23]), .O(n68768));
    defparam n9618_bdd_4_lut_51727.LUT_INIT = 16'he4aa;
    SB_LUT4 n68768_bdd_4_lut (.I0(n68768), .I1(duty[11]), .I2(n259), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[11]));
    defparam n68768_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51722 (.I0(n9618), .I1(n431), .I2(current[10]), 
            .I3(duty[23]), .O(n68762));
    defparam n9618_bdd_4_lut_51722.LUT_INIT = 16'he4aa;
    SB_LUT4 n68762_bdd_4_lut (.I0(n68762), .I1(duty[10]), .I2(n260), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[10]));
    defparam n68762_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14154_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[6]), .I2(n6_adj_5756), 
            .I3(n25145), .O(n29897));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14154_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13740_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n58139), .I3(GND_net), .O(n29483));   // verilog/coms.v(130[12] 305[6])
    defparam i13740_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9618_bdd_4_lut_51717 (.I0(n9618), .I1(n432), .I2(current[9]), 
            .I3(duty[23]), .O(n68756));
    defparam n9618_bdd_4_lut_51717.LUT_INIT = 16'he4aa;
    SB_LUT4 n68756_bdd_4_lut (.I0(n68756), .I1(duty[9]), .I2(n261), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n68756_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(current[11]), .I1(current_limit[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14155_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[7]), .I2(n6_adj_5756), 
            .I3(n25112), .O(n29898));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14155_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14156_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[8]), .I2(n5_adj_5810), 
            .I3(n25141), .O(n29899));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14156_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14157_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[9]), .I2(n5_adj_5757), 
            .I3(n25141), .O(n29900));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14157_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48829_2_lut (.I0(n68783), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65553));
    defparam i48829_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14158_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[10]), .I2(n5_adj_5755), 
            .I3(n25141), .O(n29901));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14158_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14159_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[11]), .I2(n6_adj_5754), 
            .I3(n25112), .O(n29902));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14159_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50417_3_lut (.I0(n68963), .I1(n68645), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67433));
    defparam i50417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14160_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[12]), .I2(n38922), 
            .I3(n25151), .O(n29903));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14160_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5688));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50164_4_lut (.I0(n9_adj_5734), .I1(n7_adj_5736), .I2(current[2]), 
            .I3(current_limit[2]), .O(n67180));
    defparam i50164_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50547_4_lut (.I0(n15_adj_5688), .I1(n13_adj_5689), .I2(n11_adj_5691), 
            .I3(n67180), .O(n67563));
    defparam i50547_4_lut.LUT_INIT = 16'hfeff;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27262), 
            .D(n1324), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i14161_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[15]), .I2(n38922), 
            .I3(n25112), .O(n29904));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14161_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 n9618_bdd_4_lut_51936 (.I0(n9618), .I1(n441), .I2(current[0]), 
            .I3(duty[23]), .O(n69020));
    defparam n9618_bdd_4_lut_51936.LUT_INIT = 16'he4aa;
    SB_LUT4 i50545_4_lut (.I0(n21), .I1(n19_adj_5685), .I2(n17_adj_5686), 
            .I3(n67563), .O(n67561));
    defparam i50545_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1791 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n58022));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_1791.LUT_INIT = 16'h2222;
    SB_LUT4 n69020_bdd_4_lut (.I0(n69020), .I1(duty[0]), .I2(n270), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n69020_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_238_10_lut (.I0(current[8]), .I1(duty[11]), .I2(n68604), 
            .I3(n51100), .O(n262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_10_lut.LUT_INIT = 16'hA3AC;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27262), 
            .D(n1323), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27262), 
            .D(n1322), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i13310_3_lut_4_lut (.I0(n1881), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3827), .O(n29053));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13310_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i14163_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n61676), 
            .I3(n27), .O(n29906));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14163_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13309_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29052));   // verilog/coms.v(130[12] 305[6])
    defparam i13309_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13308_3_lut_4_lut (.I0(n1933), .I1(b_prev_adj_5760), .I2(a_new_adj_5905[1]), 
            .I3(position_31__N_3827_adj_5761), .O(n29051));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13308_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_DFF read_203 (.Q(state_7__N_3916[0]), .C(clk16MHz), .D(n60966));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i14164_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n61604), 
            .I3(n27), .O(n29907));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14164_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51702 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[1]), .O(n68738));
    defparam byte_transmit_counter_0__bdd_4_lut_51702.LUT_INIT = 16'he4aa;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n57628));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27262), 
            .D(n1321), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 n68738_bdd_4_lut (.I0(n68738), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20] [2]), .I3(byte_transmit_counter[1]), 
            .O(n68741));
    defparam n68738_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13297_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5939[1]), 
            .I2(r_SM_Main_adj_5939[2]), .I3(n6_adj_5836), .O(n29040));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13297_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_CARRY add_157_19 (.CI(n51130), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n51131));
    SB_LUT4 dti_counter_1929_add_4_9_lut (.I0(n65537), .I1(n38795), .I2(dti_counter[7]), 
            .I3(n51990), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 dti_counter_1929_add_4_8_lut (.I0(n65536), .I1(n38795), .I2(dti_counter[6]), 
            .I3(n51989), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 add_157_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n51116), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_157_5 (.CI(n51116), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n51117));
    SB_CARRY dti_counter_1929_add_4_8 (.CI(n51989), .I0(n38795), .I1(dti_counter[6]), 
            .CO(n51990));
    SB_LUT4 i14165_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n61658), 
            .I3(n27), .O(n29908));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14165_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 dti_counter_1929_add_4_7_lut (.I0(n65535), .I1(n38795), .I2(dti_counter[5]), 
            .I3(n51988), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i23139_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i23139_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY dti_counter_1929_add_4_7 (.CI(n51988), .I0(n38795), .I1(dti_counter[5]), 
            .CO(n51989));
    SB_LUT4 dti_counter_1929_add_4_6_lut (.I0(n65534), .I1(n38795), .I2(dti_counter[4]), 
            .I3(n51987), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i51588_1_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n59879), 
            .I3(n59877), .O(n68604));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51588_1_lut_4_lut.LUT_INIT = 16'h4c5d;
    SB_LUT4 i1_4_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n59879), 
            .I3(n59877), .O(n209));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb3a2;
    SB_LUT4 i23138_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i23138_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY dti_counter_1929_add_4_6 (.CI(n51987), .I0(n38795), .I1(dti_counter[4]), 
            .CO(n51988));
    SB_LUT4 i23221_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i23221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 dti_counter_1929_add_4_5_lut (.I0(n65533), .I1(n38795), .I2(dti_counter[3]), 
            .I3(n51986), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1929_add_4_5 (.CI(n51986), .I0(n38795), .I1(dti_counter[3]), 
            .CO(n51987));
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27262), 
            .D(n1325), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5749));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 dti_counter_1929_add_4_4_lut (.I0(n65532), .I1(n38795), .I2(dti_counter[2]), 
            .I3(n51985), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_1929_add_4_4 (.CI(n51985), .I0(n38795), .I1(dti_counter[2]), 
            .CO(n51986));
    SB_DFFESR GHC_198 (.Q(GHC), .C(clk16MHz), .E(n27211), .D(GHC_N_391), 
            .R(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_196 (.Q(GHB), .C(clk16MHz), .E(n27211), .D(GHB_N_377), 
            .R(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i49042_2_lut_4_lut (.I0(current[8]), .I1(duty[8]), .I2(current[4]), 
            .I3(duty[4]), .O(n66058));
    defparam i49042_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 dti_counter_1929_add_4_3_lut (.I0(n65531), .I1(n38795), .I2(dti_counter[1]), 
            .I3(n51984), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_DFFESR GHA_194 (.Q(GHA), .C(clk16MHz), .E(n27211), .D(GHA_N_355), 
            .R(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY dti_counter_1929_add_4_3 (.CI(n51984), .I0(n38795), .I1(dti_counter[1]), 
            .CO(n51985));
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_5869), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i14166_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n61640), 
            .I3(n27), .O(n29909));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14166_4_lut.LUT_INIT = 16'hccca;
    SB_DFFESR GLA_195 (.Q(INLA_c_0), .C(clk16MHz), .E(n27211), .D(GLA_N_372), 
            .R(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLB_197 (.Q(INLB_c_0), .C(clk16MHz), .E(n27211), .D(GLB_N_386), 
            .R(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27262), 
            .D(n1320), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 dti_counter_1929_add_4_2_lut (.I0(n65488), .I1(n2952), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1929_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5747));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR GLC_199 (.Q(INLC_c_0), .C(clk16MHz), .E(n27211), .D(GLC_N_400), 
            .R(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY dti_counter_1929_add_4_2 (.CI(VCC_net), .I0(n2952), .I1(dti_counter[0]), 
            .CO(n51984));
    SB_LUT4 add_157_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n51115), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27262), 
            .D(n1319), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    GND i1 (.Y(GND_net));
    SB_LUT4 i14167_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n61586), 
            .I3(n27), .O(n29910));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14167_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13695_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n60939), .I3(GND_net), .O(n29438));   // verilog/coms.v(130[12] 305[6])
    defparam i13695_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13466_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n27972), 
            .I3(GND_net), .O(n29209));   // verilog/coms.v(130[12] 305[6])
    defparam i13466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1792 (.I0(n58777), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[24] [1]), .I3(n58819), .O(n10_adj_5841));
    defparam i4_4_lut_adj_1792.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5762));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13463_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n27972), 
            .I3(GND_net), .O(n29206));   // verilog/coms.v(130[12] 305[6])
    defparam i13463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1793 (.I0(state[0]), .I1(n23_adj_5865), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5719));
    defparam i1_2_lut_adj_1793.LUT_INIT = 16'h2222;
    SB_LUT4 i13_4_lut (.I0(n111), .I1(n39366), .I2(state[1]), .I3(n4_adj_5719), 
            .O(n5_adj_5856));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i5217_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5217_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i14168_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n61622), 
            .I3(n27), .O(n29911));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14168_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5219_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5219_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i5221_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i5221_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i5223_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i5223_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(delay_counter[28]), .I1(delay_counter[30]), 
            .I2(delay_counter[25]), .I3(delay_counter[24]), .O(n6_adj_5720));
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i14169_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n61550), 
            .I3(n27), .O(n29912));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14169_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4_4_lut_adj_1795 (.I0(delay_counter[27]), .I1(delay_counter[26]), 
            .I2(delay_counter[29]), .I3(n6_adj_5720), .O(n24998));
    defparam i4_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i4193_4_lut (.I0(n25007), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5769));
    defparam i4193_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5769), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n60887));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5691));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5689));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5734));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5686));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5736));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5685));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(current[10]), .I1(current_limit[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_238_10 (.CI(n51100), .I0(duty[11]), .I1(n68604), .CO(n51101));
    SB_LUT4 LessThan_20_i9_2_lut (.I0(duty[4]), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(n60887), .I1(delay_counter[18]), .I2(n25004), 
            .I3(GND_net), .O(n60510));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_20_i7_2_lut (.I0(duty[3]), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_157_4 (.CI(n51115), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n51116));
    SB_LUT4 LessThan_20_i11_2_lut (.I0(duty[5]), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i13_2_lut (.I0(duty[6]), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(duty[8]), .I1(n338), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(duty[7]), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(duty[9]), .I1(n337), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1796 (.I0(delay_counter[23]), .I1(n60510), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5850));
    defparam i2_4_lut_adj_1796.LUT_INIT = 16'heaaa;
    SB_CARRY add_238_4 (.CI(n51094), .I0(duty[5]), .I1(n68604), .CO(n51095));
    SB_LUT4 add_157_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n51114), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1797 (.I0(n7_adj_5850), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n24998), .O(n62));
    defparam i4_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1798 (.I0(r_SM_Main_adj_5939[0]), .I1(o_Rx_DV_N_3488[24]), 
            .I2(n27), .I3(GND_net), .O(n14_adj_5855));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i5_3_lut_adj_1798.LUT_INIT = 16'h0202;
    SB_LUT4 i2_3_lut_adj_1799 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25004));
    defparam i2_3_lut_adj_1799.LUT_INIT = 16'hfefe;
    SB_LUT4 add_238_9_lut (.I0(current[7]), .I1(duty[10]), .I2(n68604), 
            .I3(n51099), .O(n263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i5_3_lut_adj_1800 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14_adj_5848));
    defparam i5_3_lut_adj_1800.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(delay_counter[8]), .I1(delay_counter[7]), .I2(delay_counter[1]), 
            .I3(delay_counter[0]), .O(n15_adj_5847));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5847), .I1(delay_counter[2]), .I2(n14_adj_5848), 
            .I3(delay_counter[6]), .O(n25007));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1801 (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5722));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i6_4_lut_adj_1801.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1802 (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5723));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i5_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5738));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i6_4_lut_adj_1803 (.I0(n29), .I1(o_Rx_DV_N_3488[12]), .I2(n23_adj_5840), 
            .I3(n4894), .O(n15_adj_5854));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i6_4_lut_adj_1803.LUT_INIT = 16'h0001;
    SB_LUT4 i23151_4_lut (.I0(n13_adj_5723), .I1(baudrate[0]), .I2(n14_adj_5722), 
            .I3(n25117), .O(n38797));
    defparam i23151_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 i1_2_lut_adj_1804 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5859));
    defparam i1_2_lut_adj_1804.LUT_INIT = 16'heeee;
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27262), 
            .D(n1318), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i8_4_lut_adj_1805 (.I0(n15_adj_5854), .I1(n1), .I2(n14_adj_5855), 
            .I3(r_SM_Main_adj_5939[1]), .O(n69042));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i8_4_lut_adj_1805.LUT_INIT = 16'h8000;
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27262), 
            .D(n1317), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27262), 
            .D(n1316), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i2_4_lut_adj_1806 (.I0(delay_counter[9]), .I1(n4_adj_5859), 
            .I2(delay_counter[10]), .I3(n25007), .O(n60858));
    defparam i2_4_lut_adj_1806.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1807 (.I0(n60858), .I1(n25004), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n60747));
    defparam i2_4_lut_adj_1807.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5727));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY add_238_9 (.CI(n51099), .I0(duty[10]), .I1(n68604), .CO(n51100));
    SB_CARRY add_157_3 (.CI(n51114), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n51115));
    SB_LUT4 i2_4_lut_adj_1808 (.I0(delay_counter[22]), .I1(n60747), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5728));
    defparam i2_4_lut_adj_1808.LUT_INIT = 16'ha8a0;
    SB_LUT4 add_238_8_lut (.I0(current[6]), .I1(duty[9]), .I2(n68604), 
            .I3(n51098), .O(n264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_157_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam add_157_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY add_157_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n51114));
    SB_LUT4 i23219_4_lut (.I0(n7_adj_5728), .I1(delay_counter[31]), .I2(n24998), 
            .I3(n8_adj_5727), .O(n1405));   // verilog/TinyFPGA_B.v(379[14:38])
    defparam i23219_4_lut.LUT_INIT = 16'h3230;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF dti_counter_1929__i1 (.Q(dti_counter[1]), .C(clk16MHz), .D(n54));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i23275_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(365[12:35])
    defparam i23275_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45887_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n62903));
    defparam i45887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45888_4_lut (.I0(n62903), .I1(n27600), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n62904));
    defparam i45888_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45886_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n62902));
    defparam i45886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i592_2_lut (.I0(n1405), .I1(n38797), .I2(GND_net), .I3(GND_net), 
            .O(n2961));   // verilog/TinyFPGA_B.v(383[18] 385[12])
    defparam i592_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14171_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[1]), 
            .I2(n10_adj_5833), .I3(n25119), .O(n29914));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14171_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i45670_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n62677));
    defparam i45670_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51568_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6579), .I2(n62677), 
            .I3(n25_adj_5852), .O(n17_adj_5851));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i51568_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i14172_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[2]), 
            .I2(n4_adj_5752), .I3(n25136), .O(n29915));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14172_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_238_3_lut (.I0(current[1]), .I1(duty[4]), .I2(n68604), 
            .I3(n51093), .O(n269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i14173_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[3]), 
            .I2(n4_adj_5752), .I3(n25119), .O(n29916));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14173_4_lut.LUT_INIT = 16'hccca;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
           .D(n57676));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i13451_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n27972), 
            .I3(GND_net), .O(n29194));   // verilog/coms.v(130[12] 305[6])
    defparam i13451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13448_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n27972), 
            .I3(GND_net), .O(n29191));   // verilog/coms.v(130[12] 305[6])
    defparam i13448_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27262), 
            .D(n1315), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27262), 
            .D(n1314), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10_adj_5733), .I1(current_limit[7]), 
            .I2(n15_adj_5688), .I3(GND_net), .O(n12_adj_5690));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n56586));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i13445_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n27972), 
            .I3(GND_net), .O(n29188));   // verilog/coms.v(130[12] 305[6])
    defparam i13445_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27262), 
            .D(n1313), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 add_238_23_lut (.I0(current[15]), .I1(duty[23]), .I2(n68604), 
            .I3(n51113), .O(n249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_23_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i14174_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[4]), 
            .I2(n4_adj_5753), .I3(n25136), .O(n29917));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14174_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_238_22_lut (.I0(current[15]), .I1(duty[23]), .I2(n68604), 
            .I3(n51112), .O(n250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_22_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_238_22 (.CI(n51112), .I0(duty[23]), .I1(n68604), .CO(n51113));
    SB_LUT4 add_238_21_lut (.I0(current[15]), .I1(duty[22]), .I2(n68604), 
            .I3(n51111), .O(n251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_21_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_238_8 (.CI(n51098), .I0(duty[9]), .I1(n68604), .CO(n51099));
    SB_LUT4 i13441_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n7_adj_5862), 
            .I3(GND_net), .O(n29184));   // verilog/coms.v(130[12] 305[6])
    defparam i13441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13422_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n7_adj_5862), 
            .I3(GND_net), .O(n29165));   // verilog/coms.v(130[12] 305[6])
    defparam i13422_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14175_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[5]), 
            .I2(n4_adj_5753), .I3(n25119), .O(n29918));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14175_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51350_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[4] [5]), .I2(n7_adj_5862), 
            .I3(GND_net), .O(n57504));   // verilog/coms.v(94[13:20])
    defparam i51350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13370_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n7_adj_5862), 
            .I3(GND_net), .O(n29113));   // verilog/coms.v(130[12] 305[6])
    defparam i13370_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27262), 
            .D(n1312), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i14176_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[6]), 
            .I2(n38965), .I3(n25136), .O(n29919));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14176_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13367_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n7_adj_5862), 
            .I3(GND_net), .O(n29110));   // verilog/coms.v(130[12] 305[6])
    defparam i13367_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_238_21 (.CI(n51111), .I0(duty[22]), .I1(n68604), .CO(n51112));
    SB_LUT4 i13364_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n7_adj_5862), 
            .I3(GND_net), .O(n29107));   // verilog/coms.v(130[12] 305[6])
    defparam i13364_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_238_7_lut (.I0(current[5]), .I1(duty[8]), .I2(n68604), 
            .I3(n51097), .O(n265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_238_3 (.CI(n51093), .I0(duty[4]), .I1(n68604), .CO(n51094));
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27262), 
            .D(n1311), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27262), 
            .D(n1310), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_CARRY add_238_7 (.CI(n51097), .I0(duty[8]), .I1(n68604), .CO(n51098));
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27262), 
            .D(n1309), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 add_238_2_lut (.I0(GND_net), .I1(duty[3]), .I2(n211), .I3(GND_net), 
            .O(n1828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14177_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[7]), 
            .I2(n38965), .I3(n25119), .O(n29920));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14177_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 add_238_20_lut (.I0(current[15]), .I1(duty[21]), .I2(n68604), 
            .I3(n51110), .O(n252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_20_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_238_20 (.CI(n51110), .I0(duty[21]), .I1(n68604), .CO(n51111));
    SB_DFF dti_counter_1929__i2 (.Q(dti_counter[2]), .C(clk16MHz), .D(n53));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 n9618_bdd_4_lut_51712 (.I0(n9618), .I1(n433), .I2(current[8]), 
            .I3(duty[23]), .O(n68726));
    defparam n9618_bdd_4_lut_51712.LUT_INIT = 16'he4aa;
    SB_LUT4 n68726_bdd_4_lut (.I0(n68726), .I1(duty[8]), .I2(n262), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n68726_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51687 (.I0(n9618), .I1(n434), .I2(current[7]), 
            .I3(duty[23]), .O(n68720));
    defparam n9618_bdd_4_lut_51687.LUT_INIT = 16'he4aa;
    SB_LUT4 n68720_bdd_4_lut (.I0(n68720), .I1(duty[7]), .I2(n263), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n68720_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF dti_counter_1929__i3 (.Q(dti_counter[3]), .C(clk16MHz), .D(n52));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1929__i4 (.Q(dti_counter[4]), .C(clk16MHz), .D(n51));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1929__i5 (.Q(dti_counter[5]), .C(clk16MHz), .D(n50));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1929__i6 (.Q(dti_counter[6]), .C(clk16MHz), .D(n49));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_1929__i7 (.Q(dti_counter[7]), .C(clk16MHz), .D(n48));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27262), 
            .D(n1308), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27262), 
            .D(n1307), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27262), 
            .D(n1306), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27262), 
            .D(n1305), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27262), 
            .D(n1304), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27262), 
            .D(n1303), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27262), 
            .D(n1302), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27262), 
            .D(n1301), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27262), 
            .D(n1300), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27262), 
            .D(n1299), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27262), 
            .D(n1298), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27262), 
            .D(n1297), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27262), 
            .D(n1296), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27262), 
            .D(n1295), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27262), 
            .D(n1294), .R(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i1_2_lut_adj_1809 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5721));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1809.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1810 (.I0(n58680), .I1(n58312), .I2(n58857), 
            .I3(n6_adj_5721), .O(n58185));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1810.LUT_INIT = 16'h6996;
    SB_DFF reset_204 (.Q(reset), .C(clk16MHz), .D(n56676));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_238_19_lut (.I0(current[15]), .I1(duty[20]), .I2(n68604), 
            .I3(n51109), .O(n253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_19_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i23150_1_lut_2_lut (.I0(n22497), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n2952));
    defparam i23150_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 n9618_bdd_4_lut_51682 (.I0(n9618), .I1(n435), .I2(current[6]), 
            .I3(duty[23]), .O(n68714));
    defparam n9618_bdd_4_lut_51682.LUT_INIT = 16'he4aa;
    SB_LUT4 i14199_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n58147), 
            .I3(GND_net), .O(n29942));   // verilog/coms.v(130[12] 305[6])
    defparam i14199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14202_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n58147), 
            .I3(GND_net), .O(n29945));   // verilog/coms.v(130[12] 305[6])
    defparam i14202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5764));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5779));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5780));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14205_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n58147), 
            .I3(GND_net), .O(n29948));   // verilog/coms.v(130[12] 305[6])
    defparam i14205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5781));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5782));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5783));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5784));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1811 (.I0(n25269), .I1(n58321), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n53279));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1811.LUT_INIT = 16'h9696;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5785));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13553_3_lut (.I0(\data_in_frame[8] [0]), .I1(rx_data[0]), .I2(n58140), 
            .I3(GND_net), .O(n29296));   // verilog/coms.v(130[12] 305[6])
    defparam i13553_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5798));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5799));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5800));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5801));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5802));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14208_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n58147), 
            .I3(GND_net), .O(n29951));   // verilog/coms.v(130[12] 305[6])
    defparam i14208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13556_3_lut (.I0(\data_in_frame[8] [1]), .I1(rx_data[1]), .I2(n58140), 
            .I3(GND_net), .O(n29299));   // verilog/coms.v(130[12] 305[6])
    defparam i13556_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5804));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5805));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5806));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5807));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5808));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5809));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5765));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5766));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5770));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13559_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n58140), 
            .I3(GND_net), .O(n29302));   // verilog/coms.v(130[12] 305[6])
    defparam i13559_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5718));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5717));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_238_19 (.CI(n51109), .I0(duty[20]), .I1(n68604), .CO(n51110));
    SB_LUT4 add_4749_21_lut (.I0(GND_net), .I1(n13038), .I2(encoder1_position[21]), 
            .I3(n51486), .O(n9927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4749_20_lut (.I0(GND_net), .I1(n13039), .I2(encoder1_position[20]), 
            .I3(n51485), .O(n9928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_20 (.CI(n51485), .I0(n13039), .I1(encoder1_position[20]), 
            .CO(n51486));
    SB_LUT4 unary_minus_19_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5716));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13562_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n58140), 
            .I3(GND_net), .O(n29305));   // verilog/coms.v(130[12] 305[6])
    defparam i13562_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13865_3_lut (.I0(\data_in_frame[20] [6]), .I1(rx_data[6]), 
            .I2(n28002), .I3(GND_net), .O(n29608));   // verilog/coms.v(130[12] 305[6])
    defparam i13865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_4749_19_lut (.I0(GND_net), .I1(n13040), .I2(encoder1_position[19]), 
            .I3(n51484), .O(n9929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13565_3_lut (.I0(\data_in_frame[8] [4]), .I1(rx_data[4]), .I2(n58140), 
            .I3(GND_net), .O(n29308));   // verilog/coms.v(130[12] 305[6])
    defparam i13565_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4749_19 (.CI(n51484), .I0(n13040), .I1(encoder1_position[19]), 
            .CO(n51485));
    SB_LUT4 add_4749_18_lut (.I0(GND_net), .I1(n13041), .I2(encoder1_position[18]), 
            .I3(n51483), .O(n9930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_18 (.CI(n51483), .I0(n13041), .I1(encoder1_position[18]), 
            .CO(n51484));
    SB_LUT4 add_4749_17_lut (.I0(GND_net), .I1(n13042), .I2(encoder1_position[17]), 
            .I3(n51482), .O(n9931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5715));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_238_6_lut (.I0(current[4]), .I1(duty[7]), .I2(n68604), 
            .I3(n51096), .O(n266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_19_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5712));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_238_18_lut (.I0(current[15]), .I1(duty[19]), .I2(n68604), 
            .I3(n51108), .O(n254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_18_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_4749_17 (.CI(n51482), .I0(n13042), .I1(encoder1_position[17]), 
            .CO(n51483));
    SB_LUT4 i13862_3_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(n28002), .I3(GND_net), .O(n29605));   // verilog/coms.v(130[12] 305[6])
    defparam i13862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5711));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5710));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5709));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4749_16_lut (.I0(GND_net), .I1(n13043), .I2(encoder1_position[16]), 
            .I3(n51481), .O(n9932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_16 (.CI(n51481), .I0(n13043), .I1(encoder1_position[16]), 
            .CO(n51482));
    SB_LUT4 unary_minus_19_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5708));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1812 (.I0(n58238), .I1(n58952), .I2(n1191), .I3(n58845), 
            .O(n20_adj_5815));   // verilog/coms.v(100[12:26])
    defparam i8_4_lut_adj_1812.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n58748), .I1(\data_out_frame[5] [5]), .I2(\data_out_frame[17] [3]), 
            .I3(n58925), .O(n19_adj_5816));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n58446), .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[11] [0]), 
            .I3(\data_out_frame[15] [2]), .O(n21_adj_5814));   // verilog/coms.v(100[12:26])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_19_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5707));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_1_lut (.I0(current[15]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4749_15_lut (.I0(GND_net), .I1(n13044), .I2(encoder1_position[15]), 
            .I3(n51480), .O(n9933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13568_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n58140), 
            .I3(GND_net), .O(n29311));   // verilog/coms.v(130[12] 305[6])
    defparam i13568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1089_i1_4_lut (.I0(n65376), .I1(n25), .I2(n296), .I3(n356), 
            .O(n5093));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam mux_1089_i1_4_lut.LUT_INIT = 16'hcac0;
    SB_CARRY add_4749_15 (.CI(n51480), .I0(n13044), .I1(encoder1_position[15]), 
            .CO(n51481));
    SB_LUT4 i13859_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n28002), .I3(GND_net), .O(n29602));   // verilog/coms.v(130[12] 305[6])
    defparam i13859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13571_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n58140), 
            .I3(GND_net), .O(n29314));   // verilog/coms.v(130[12] 305[6])
    defparam i13571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_4749_14_lut (.I0(GND_net), .I1(n13045), .I2(encoder1_position[14]), 
            .I3(n51479), .O(n9934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13856_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n28002), .I3(GND_net), .O(n29599));   // verilog/coms.v(130[12] 305[6])
    defparam i13856_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4749_14 (.CI(n51479), .I0(n13045), .I1(encoder1_position[14]), 
            .CO(n51480));
    SB_LUT4 i11_3_lut (.I0(n21_adj_5814), .I1(n19_adj_5816), .I2(n20_adj_5815), 
            .I3(GND_net), .O(n53988));   // verilog/coms.v(100[12:26])
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13574_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n58140), 
            .I3(GND_net), .O(n29317));   // verilog/coms.v(130[12] 305[6])
    defparam i13574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13577_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n58141), 
            .I3(GND_net), .O(n29320));   // verilog/coms.v(130[12] 305[6])
    defparam i13577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_4749_13_lut (.I0(GND_net), .I1(n13046), .I2(encoder1_position[13]), 
            .I3(n51478), .O(n9935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_13 (.CI(n51478), .I0(n13046), .I1(encoder1_position[13]), 
            .CO(n51479));
    SB_LUT4 add_4749_12_lut (.I0(GND_net), .I1(n13047), .I2(encoder1_position[12]), 
            .I3(n51477), .O(n9936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_12 (.CI(n51477), .I0(n13047), .I1(encoder1_position[12]), 
            .CO(n51478));
    SB_LUT4 add_4749_11_lut (.I0(GND_net), .I1(n13048), .I2(encoder1_position[11]), 
            .I3(n51476), .O(n9937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_11 (.CI(n51476), .I0(n13048), .I1(encoder1_position[11]), 
            .CO(n51477));
    SB_LUT4 add_4749_10_lut (.I0(GND_net), .I1(n13049), .I2(encoder1_position[10]), 
            .I3(n51475), .O(n9938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13580_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n58141), 
            .I3(GND_net), .O(n29323));   // verilog/coms.v(130[12] 305[6])
    defparam i13580_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4749_10 (.CI(n51475), .I0(n13049), .I1(encoder1_position[10]), 
            .CO(n51476));
    SB_LUT4 i13850_3_lut (.I0(\data_in_frame[20] [1]), .I1(rx_data[1]), 
            .I2(n28002), .I3(GND_net), .O(n29593));   // verilog/coms.v(130[12] 305[6])
    defparam i13850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13583_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n58141), 
            .I3(GND_net), .O(n29326));   // verilog/coms.v(130[12] 305[6])
    defparam i13583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n68714_bdd_4_lut (.I0(n68714), .I1(duty[6]), .I2(n264), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n68714_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_18_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5700));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_5699));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13586_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n58141), 
            .I3(GND_net), .O(n29329));   // verilog/coms.v(130[12] 305[6])
    defparam i13586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5698));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5697));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4749_9_lut (.I0(GND_net), .I1(n13050), .I2(encoder1_position[9]), 
            .I3(n51474), .O(n9939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_9 (.CI(n51474), .I0(n13050), .I1(encoder1_position[9]), 
            .CO(n51475));
    SB_LUT4 unary_minus_18_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5696));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4749_8_lut (.I0(GND_net), .I1(n13051), .I2(encoder1_position[8]), 
            .I3(n51473), .O(n9940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_8 (.CI(n51473), .I0(n13051), .I1(encoder1_position[8]), 
            .CO(n51474));
    SB_LUT4 unary_minus_18_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5695));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5694));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13589_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n58141), 
            .I3(GND_net), .O(n29332));   // verilog/coms.v(130[12] 305[6])
    defparam i13589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5693));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5692));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5735), .I1(current_limit[9]), 
            .I2(n19_adj_5685), .I3(GND_net), .O(n16_adj_5687));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4749_7_lut (.I0(GND_net), .I1(n13052), .I2(encoder1_position[7]), 
            .I3(n51472), .O(n9941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_7 (.CI(n51472), .I0(n13052), .I1(encoder1_position[7]), 
            .CO(n51473));
    SB_LUT4 add_4749_6_lut (.I0(GND_net), .I1(n13053), .I2(encoder1_position[6]), 
            .I3(n51471), .O(n9942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_6 (.CI(n51471), .I0(n13053), .I1(encoder1_position[6]), 
            .CO(n51472));
    SB_LUT4 add_4749_5_lut (.I0(GND_net), .I1(n13054), .I2(encoder1_position[5]), 
            .I3(n51470), .O(n9943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_5 (.CI(n51470), .I0(n13054), .I1(encoder1_position[5]), 
            .CO(n51471));
    SB_LUT4 add_4749_4_lut (.I0(GND_net), .I1(n13055), .I2(encoder1_position[4]), 
            .I3(n51469), .O(n9944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_4 (.CI(n51469), .I0(n13055), .I1(encoder1_position[4]), 
            .CO(n51470));
    SB_LUT4 i49484_2_lut (.I0(displacement[0]), .I1(n15_adj_5732), .I2(GND_net), 
            .I3(GND_net), .O(n65364));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam i49484_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13592_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n58141), 
            .I3(GND_net), .O(n29335));   // verilog/coms.v(130[12] 305[6])
    defparam i13592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_4749_3_lut (.I0(GND_net), .I1(n13056), .I2(encoder1_position[3]), 
            .I3(n51468), .O(n9945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4749_3 (.CI(n51468), .I0(n13056), .I1(encoder1_position[3]), 
            .CO(n51469));
    SB_CARRY add_238_2 (.CI(GND_net), .I0(duty[3]), .I1(n211), .CO(n51093));
    SB_LUT4 add_4749_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(n9946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4749_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48665_2_lut (.I0(displacement[1]), .I1(n15_adj_5732), .I2(GND_net), 
            .I3(GND_net), .O(n65475));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam i48665_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_4749_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n51468));
    SB_LUT4 add_4748_23_lut (.I0(GND_net), .I1(n9927), .I2(encoder1_position[23]), 
            .I3(n51467), .O(encoder1_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_238_6 (.CI(n51096), .I0(duty[7]), .I1(n68604), .CO(n51097));
    SB_CARRY add_238_18 (.CI(n51108), .I0(duty[19]), .I1(n68604), .CO(n51109));
    SB_LUT4 i48664_2_lut (.I0(displacement[2]), .I1(n15_adj_5732), .I2(GND_net), 
            .I3(GND_net), .O(n65474));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam i48664_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_4748_22_lut (.I0(GND_net), .I1(n9928), .I2(encoder1_position[22]), 
            .I3(n51466), .O(encoder1_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_22 (.CI(n51466), .I0(n9928), .I1(encoder1_position[22]), 
            .CO(n51467));
    SB_LUT4 add_4748_21_lut (.I0(GND_net), .I1(n9929), .I2(encoder1_position[21]), 
            .I3(n51465), .O(encoder1_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13595_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n58141), 
            .I3(GND_net), .O(n29338));   // verilog/coms.v(130[12] 305[6])
    defparam i13595_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4748_21 (.CI(n51465), .I0(n9929), .I1(encoder1_position[21]), 
            .CO(n51466));
    SB_LUT4 add_4748_20_lut (.I0(GND_net), .I1(n9930), .I2(encoder1_position[20]), 
            .I3(n51464), .O(encoder1_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_20 (.CI(n51464), .I0(n9930), .I1(encoder1_position[20]), 
            .CO(n51465));
    SB_LUT4 i27_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(100[12:26])
    defparam i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4748_19_lut (.I0(GND_net), .I1(n9931), .I2(encoder1_position[19]), 
            .I3(n51463), .O(encoder1_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_19 (.CI(n51463), .I0(n9931), .I1(encoder1_position[19]), 
            .CO(n51464));
    SB_LUT4 add_4748_18_lut (.I0(GND_net), .I1(n9932), .I2(encoder1_position[18]), 
            .I3(n51462), .O(encoder1_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_18 (.CI(n51462), .I0(n9932), .I1(encoder1_position[18]), 
            .CO(n51463));
    SB_LUT4 add_4748_17_lut (.I0(GND_net), .I1(n9933), .I2(encoder1_position[17]), 
            .I3(n51461), .O(encoder1_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_17 (.CI(n51461), .I0(n9933), .I1(encoder1_position[17]), 
            .CO(n51462));
    SB_LUT4 add_4748_16_lut (.I0(GND_net), .I1(n9934), .I2(encoder1_position[16]), 
            .I3(n51460), .O(encoder1_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_238_17_lut (.I0(current[15]), .I1(duty[18]), .I2(n68604), 
            .I3(n51107), .O(n255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_17_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n57886));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n58004));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_CARRY add_4748_16 (.CI(n51460), .I0(n9934), .I1(encoder1_position[16]), 
            .CO(n51461));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n57892));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_LUT4 mux_253_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_91[3]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1815 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n57893));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1815.LUT_INIT = 16'h2300;
    SB_LUT4 i13598_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n58141), 
            .I3(GND_net), .O(n29341));   // verilog/coms.v(130[12] 305[6])
    defparam i13598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1816 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n57885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1816.LUT_INIT = 16'h2300;
    SB_LUT4 mux_253_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_91[4]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_4748_15_lut (.I0(GND_net), .I1(n9935), .I2(encoder1_position[15]), 
            .I3(n51459), .O(encoder1_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_15 (.CI(n51459), .I0(n9935), .I1(encoder1_position[15]), 
            .CO(n51460));
    SB_LUT4 add_4748_14_lut (.I0(GND_net), .I1(n9936), .I2(encoder1_position[14]), 
            .I3(n51458), .O(encoder1_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_14 (.CI(n51458), .I0(n9936), .I1(encoder1_position[14]), 
            .CO(n51459));
    SB_LUT4 add_4748_13_lut (.I0(GND_net), .I1(n9937), .I2(encoder1_position[13]), 
            .I3(n51457), .O(encoder1_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_253_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13601_3_lut (.I0(\data_in_frame[10] [0]), .I1(rx_data[0]), 
            .I2(n58142), .I3(GND_net), .O(n29344));   // verilog/coms.v(130[12] 305[6])
    defparam i13601_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1817 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n57884));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1817.LUT_INIT = 16'h2300;
    SB_LUT4 mux_251_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_91[5]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n69008));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i13604_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n58142), .I3(GND_net), .O(n29347));   // verilog/coms.v(130[12] 305[6])
    defparam i13604_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4748_13 (.CI(n51457), .I0(n9937), .I1(encoder1_position[13]), 
            .CO(n51458));
    SB_LUT4 i1_4_lut_adj_1818 (.I0(hall3), .I1(commutation_state[1]), .I2(hall2), 
            .I3(hall1), .O(n57676));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hd054;
    SB_LUT4 mux_253_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_91[6]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_253_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_91[7]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_253_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1819 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58748));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1819.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1820 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n57894));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1820.LUT_INIT = 16'h2300;
    SB_LUT4 mux_251_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_91[8]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i9_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_238_17 (.CI(n51107), .I0(duty[18]), .I1(n68604), .CO(n51108));
    SB_LUT4 add_238_16_lut (.I0(current[15]), .I1(duty[17]), .I2(n68604), 
            .I3(n51106), .O(n256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_16_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i22446_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(n38105));
    defparam i22446_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i22447_3_lut (.I0(encoder0_position_scaled[9]), .I1(n38105), 
            .I2(n15_adj_5731), .I3(GND_net), .O(n38106));
    defparam i22447_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_4748_12_lut (.I0(GND_net), .I1(n9938), .I2(encoder1_position[12]), 
            .I3(n51456), .O(encoder1_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_253_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_91[10]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_253_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_91[11]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_253_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_91[12]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_253_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_91[13]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i14_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4748_12 (.CI(n51456), .I0(n9938), .I1(encoder1_position[12]), 
            .CO(n51457));
    SB_LUT4 mux_253_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_91[14]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i15_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_238_16 (.CI(n51106), .I0(duty[17]), .I1(n68604), .CO(n51107));
    SB_LUT4 mux_253_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_91[15]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_4748_11_lut (.I0(GND_net), .I1(n9939), .I2(encoder1_position[11]), 
            .I3(n51455), .O(encoder1_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_11 (.CI(n51455), .I0(n9939), .I1(encoder1_position[11]), 
            .CO(n51456));
    SB_LUT4 add_4748_10_lut (.I0(GND_net), .I1(n9940), .I2(encoder1_position[10]), 
            .I3(n51454), .O(encoder1_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_253_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_4748_10 (.CI(n51454), .I0(n9940), .I1(encoder1_position[10]), 
            .CO(n51455));
    SB_LUT4 mux_251_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_91[16]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_4748_9_lut (.I0(GND_net), .I1(n9941), .I2(encoder1_position[9]), 
            .I3(n51453), .O(encoder1_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_9 (.CI(n51453), .I0(n9941), .I1(encoder1_position[9]), 
            .CO(n51454));
    SB_LUT4 add_4748_8_lut (.I0(GND_net), .I1(n9942), .I2(encoder1_position[8]), 
            .I3(n51452), .O(encoder1_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_238_15_lut (.I0(current[15]), .I1(duty[16]), .I2(n68604), 
            .I3(n51105), .O(n257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_15_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n57883));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h2300;
    SB_LUT4 mux_253_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_91[17]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1822 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n57882));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1822.LUT_INIT = 16'h2300;
    SB_CARRY add_4748_8 (.CI(n51452), .I0(n9942), .I1(encoder1_position[8]), 
            .CO(n51453));
    SB_LUT4 add_4748_7_lut (.I0(GND_net), .I1(n9943), .I2(encoder1_position[7]), 
            .I3(n51451), .O(encoder1_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_7 (.CI(n51451), .I0(n9943), .I1(encoder1_position[7]), 
            .CO(n51452));
    SB_LUT4 i14_4_lut_adj_1823 (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(n13_adj_5845));
    defparam i14_4_lut_adj_1823.LUT_INIT = 16'h0aca;
    SB_LUT4 add_4748_6_lut (.I0(GND_net), .I1(n9944), .I2(encoder1_position[6]), 
            .I3(n51450), .O(encoder1_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_3_lut (.I0(encoder0_position_scaled[18]), .I1(n13_adj_5845), 
            .I2(n15_adj_5731), .I3(GND_net), .O(n14_adj_5843));
    defparam i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n57881));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h2300;
    SB_LUT4 mux_253_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_4748_6 (.CI(n51450), .I0(n9944), .I1(encoder1_position[6]), 
            .CO(n51451));
    SB_LUT4 mux_251_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_91[19]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1825 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n57880));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1825.LUT_INIT = 16'h2300;
    SB_LUT4 i13607_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n58142), .I3(GND_net), .O(n29350));   // verilog/coms.v(130[12] 305[6])
    defparam i13607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_4748_5_lut (.I0(GND_net), .I1(n9945), .I2(encoder1_position[5]), 
            .I3(n51449), .O(encoder1_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_5 (.CI(n51449), .I0(n9945), .I1(encoder1_position[5]), 
            .CO(n51450));
    SB_LUT4 mux_253_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_251_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_91[20]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_253_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_4748_4_lut (.I0(GND_net), .I1(n9946), .I2(encoder1_position[4]), 
            .I3(n51448), .O(encoder1_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4748_4 (.CI(n51448), .I0(n9946), .I1(encoder1_position[4]), 
            .CO(n51449));
    SB_LUT4 add_4748_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[3]), 
            .I3(n51447), .O(encoder1_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_251_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_91[21]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i22_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4748_3 (.CI(n51447), .I0(encoder1_position[1]), .I1(encoder1_position[3]), 
            .CO(n51448));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n57879));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h2300;
    SB_LUT4 add_4748_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4748_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13610_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n58142), .I3(GND_net), .O(n29353));   // verilog/coms.v(130[12] 305[6])
    defparam i13610_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4748_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n51447));
    SB_LUT4 add_4746_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(encoder1_position[19]), 
            .I3(n51446), .O(n13038)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_238_15 (.CI(n51105), .I0(duty[16]), .I1(n68604), .CO(n51106));
    SB_LUT4 add_4746_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(encoder1_position[18]), 
            .I3(n51445), .O(n13039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_19 (.CI(n51445), .I0(encoder1_position[17]), .I1(encoder1_position[18]), 
            .CO(n51446));
    SB_LUT4 add_4746_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(encoder1_position[17]), 
            .I3(n51444), .O(n13040)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_18 (.CI(n51444), .I0(encoder1_position[16]), .I1(encoder1_position[17]), 
            .CO(n51445));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n57878));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1828 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n57996));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1828.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1829 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n57995));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1829.LUT_INIT = 16'h2300;
    SB_LUT4 add_238_14_lut (.I0(current[15]), .I1(duty[15]), .I2(n68604), 
            .I3(n51104), .O(n258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_238_14_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_4746_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(encoder1_position[16]), 
            .I3(n51443), .O(n13041)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_17 (.CI(n51443), .I0(encoder1_position[15]), .I1(encoder1_position[16]), 
            .CO(n51444));
    SB_CARRY add_238_14 (.CI(n51104), .I0(duty[15]), .I1(n68604), .CO(n51105));
    SB_LUT4 add_4746_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(encoder1_position[15]), 
            .I3(n51442), .O(n13042)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_16 (.CI(n51442), .I0(encoder1_position[14]), .I1(encoder1_position[15]), 
            .CO(n51443));
    SB_LUT4 add_4746_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(encoder1_position[14]), 
            .I3(n51441), .O(n13043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_15 (.CI(n51441), .I0(encoder1_position[13]), .I1(encoder1_position[14]), 
            .CO(n51442));
    SB_LUT4 add_4746_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(encoder1_position[13]), 
            .I3(n51440), .O(n13044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_14 (.CI(n51440), .I0(encoder1_position[12]), .I1(encoder1_position[13]), 
            .CO(n51441));
    SB_LUT4 add_4746_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(encoder1_position[12]), 
            .I3(n51439), .O(n13045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_13 (.CI(n51439), .I0(encoder1_position[11]), .I1(encoder1_position[12]), 
            .CO(n51440));
    SB_LUT4 add_4746_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(encoder1_position[11]), 
            .I3(n51438), .O(n13046)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_12 (.CI(n51438), .I0(encoder1_position[10]), .I1(encoder1_position[11]), 
            .CO(n51439));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n57877));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h2300;
    SB_LUT4 add_4746_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(encoder1_position[10]), 
            .I3(n51437), .O(n13047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_11 (.CI(n51437), .I0(encoder1_position[9]), .I1(encoder1_position[10]), 
            .CO(n51438));
    SB_LUT4 add_4746_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(encoder1_position[9]), 
            .I3(n51436), .O(n13048)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_10 (.CI(n51436), .I0(encoder1_position[8]), .I1(encoder1_position[9]), 
            .CO(n51437));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n57876));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h2300;
    SB_LUT4 add_4746_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(encoder1_position[8]), 
            .I3(n51435), .O(n13049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_9 (.CI(n51435), .I0(encoder1_position[7]), .I1(encoder1_position[8]), 
            .CO(n51436));
    SB_LUT4 add_4746_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(encoder1_position[7]), 
            .I3(n51434), .O(n13050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_8 (.CI(n51434), .I0(encoder1_position[6]), .I1(encoder1_position[7]), 
            .CO(n51435));
    SB_LUT4 add_4746_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(encoder1_position[6]), 
            .I3(n51433), .O(n13051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_7 (.CI(n51433), .I0(encoder1_position[5]), .I1(encoder1_position[6]), 
            .CO(n51434));
    SB_LUT4 add_4746_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(encoder1_position[5]), 
            .I3(n51432), .O(n13052)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_6 (.CI(n51432), .I0(encoder1_position[4]), .I1(encoder1_position[5]), 
            .CO(n51433));
    SB_LUT4 add_4746_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position[4]), 
            .I3(n51431), .O(n13053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_5 (.CI(n51431), .I0(encoder1_position[3]), .I1(encoder1_position[4]), 
            .CO(n51432));
    SB_LUT4 add_4746_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[3]), 
            .I3(n51430), .O(n13054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_4 (.CI(n51430), .I0(encoder1_position[2]), .I1(encoder1_position[3]), 
            .CO(n51431));
    SB_LUT4 add_4746_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[2]), 
            .I3(n51429), .O(n13055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_3 (.CI(n51429), .I0(encoder1_position[1]), .I1(encoder1_position[2]), 
            .CO(n51430));
    SB_LUT4 add_4746_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n13056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4746_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4746_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n51429));
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n51168), .O(n356)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(n4883), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n51167), .O(n5048)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_25 (.CI(n51167), .I0(GND_net), .I1(pwm_setpoint_23__N_207), 
            .CO(n51168));
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(n4883), .I1(GND_net), .I2(n3), 
            .I3(n51166), .O(n5049)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_24 (.CI(n51166), .I0(GND_net), .I1(n3), 
            .CO(n51167));
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(n4883), .I1(GND_net), .I2(n4_adj_5692), 
            .I3(n51165), .O(n5050)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_23 (.CI(n51165), .I0(GND_net), .I1(n4_adj_5692), 
            .CO(n51166));
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(n4883), .I1(GND_net), .I2(n5_adj_5693), 
            .I3(n51164), .O(n5051)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n51164), .I0(GND_net), .I1(n5_adj_5693), 
            .CO(n51165));
    SB_LUT4 mux_253_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(n4883), .I1(GND_net), .I2(n6_adj_5694), 
            .I3(n51163), .O(n5052)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_21 (.CI(n51163), .I0(GND_net), .I1(n6_adj_5694), 
            .CO(n51164));
    SB_LUT4 mux_251_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_91[22]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(n4883), .I1(GND_net), .I2(n7_adj_5695), 
            .I3(n51162), .O(n5053)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_20 (.CI(n51162), .I0(GND_net), .I1(n7_adj_5695), 
            .CO(n51163));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n57875));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(n4883), .I1(GND_net), .I2(n8_adj_5696), 
            .I3(n51161), .O(n5054)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_19 (.CI(n51161), .I0(GND_net), .I1(n8_adj_5696), 
            .CO(n51162));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1833 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n57874));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1833.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(n4883), .I1(GND_net), .I2(n9_adj_5697), 
            .I3(n51160), .O(n5055)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_18 (.CI(n51160), .I0(GND_net), .I1(n9_adj_5697), 
            .CO(n51161));
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(n4883), .I1(GND_net), .I2(n10), 
            .I3(n51159), .O(n5056)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_17 (.CI(n51159), .I0(GND_net), .I1(n10), 
            .CO(n51160));
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(n4883), .I1(GND_net), .I2(n11_adj_5698), 
            .I3(n51158), .O(n5057)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_16 (.CI(n51158), .I0(GND_net), .I1(n11_adj_5698), 
            .CO(n51159));
    SB_LUT4 i13613_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n58142), .I3(GND_net), .O(n29356));   // verilog/coms.v(130[12] 305[6])
    defparam i13613_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(n4883), .I1(GND_net), .I2(n12_adj_5699), 
            .I3(n51157), .O(n5058)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_15 (.CI(n51157), .I0(GND_net), .I1(n12_adj_5699), 
            .CO(n51158));
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(n4883), .I1(GND_net), .I2(n13_adj_5700), 
            .I3(n51156), .O(n5059)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_14 (.CI(n51156), .I0(GND_net), .I1(n13_adj_5700), 
            .CO(n51157));
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(n4883), .I1(GND_net), .I2(n14), 
            .I3(n51155), .O(n5060)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_13 (.CI(n51155), .I0(GND_net), .I1(n14), 
            .CO(n51156));
    SB_LUT4 add_1091_25_lut (.I0(GND_net), .I1(n5047), .I2(n5070), .I3(n51406), 
            .O(n418)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1091_24_lut (.I0(GND_net), .I1(n5047), .I2(n5071), .I3(n51405), 
            .O(n419)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_24 (.CI(n51405), .I0(n5047), .I1(n5071), .CO(n51406));
    SB_LUT4 add_1091_23_lut (.I0(GND_net), .I1(n5047), .I2(n5072), .I3(n51404), 
            .O(n420)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_23 (.CI(n51404), .I0(n5047), .I1(n5072), .CO(n51405));
    SB_LUT4 add_1091_22_lut (.I0(GND_net), .I1(n5048), .I2(n5073), .I3(n51403), 
            .O(n421)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_22 (.CI(n51403), .I0(n5048), .I1(n5073), .CO(n51404));
    SB_LUT4 add_1091_21_lut (.I0(GND_net), .I1(n5049), .I2(n5074), .I3(n51402), 
            .O(n422)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_21 (.CI(n51402), .I0(n5049), .I1(n5074), .CO(n51403));
    SB_LUT4 add_1091_20_lut (.I0(GND_net), .I1(n5050), .I2(n5075), .I3(n51401), 
            .O(n423)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_20 (.CI(n51401), .I0(n5050), .I1(n5075), .CO(n51402));
    SB_LUT4 add_1091_19_lut (.I0(GND_net), .I1(n5051), .I2(n5076), .I3(n51400), 
            .O(n424)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_19 (.CI(n51400), .I0(n5051), .I1(n5076), .CO(n51401));
    SB_LUT4 add_1091_18_lut (.I0(GND_net), .I1(n5052), .I2(n5077), .I3(n51399), 
            .O(n425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1834 (.I0(control_mode[3]), .I1(control_mode[4]), 
            .I2(control_mode[2]), .I3(control_mode[6]), .O(n62052));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_CARRY add_1091_18 (.CI(n51399), .I0(n5052), .I1(n5077), .CO(n51400));
    SB_LUT4 add_1091_17_lut (.I0(GND_net), .I1(n5053), .I2(n5078), .I3(n51398), 
            .O(n426)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_17 (.CI(n51398), .I0(n5053), .I1(n5078), .CO(n51399));
    SB_LUT4 add_1091_16_lut (.I0(GND_net), .I1(n5054), .I2(n5079), .I3(n51397), 
            .O(n427)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(n62052), .I1(control_mode[7]), .I2(control_mode[5]), 
            .I3(GND_net), .O(n25130));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n57873));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h2300;
    SB_CARRY add_1091_16 (.CI(n51397), .I0(n5054), .I1(n5079), .CO(n51398));
    SB_LUT4 add_1091_15_lut (.I0(GND_net), .I1(n5055), .I2(n5080), .I3(n51396), 
            .O(n428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_15 (.CI(n51396), .I0(n5055), .I1(n5080), .CO(n51397));
    SB_LUT4 add_1091_14_lut (.I0(GND_net), .I1(n5056), .I2(n5081), .I3(n51395), 
            .O(n429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_14 (.CI(n51395), .I0(n5056), .I1(n5081), .CO(n51396));
    SB_LUT4 add_1091_13_lut (.I0(GND_net), .I1(n5057), .I2(n5082), .I3(n51394), 
            .O(n430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_13 (.CI(n51394), .I0(n5057), .I1(n5082), .CO(n51395));
    SB_LUT4 add_1091_12_lut (.I0(GND_net), .I1(n5058), .I2(n5083), .I3(n51393), 
            .O(n431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_12 (.CI(n51393), .I0(n5058), .I1(n5083), .CO(n51394));
    SB_LUT4 add_1091_11_lut (.I0(GND_net), .I1(n5059), .I2(n5084), .I3(n51392), 
            .O(n432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_11 (.CI(n51392), .I0(n5059), .I1(n5084), .CO(n51393));
    SB_LUT4 add_1091_10_lut (.I0(GND_net), .I1(n5060), .I2(n5085), .I3(n51391), 
            .O(n433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_10 (.CI(n51391), .I0(n5060), .I1(n5085), .CO(n51392));
    SB_LUT4 add_1091_9_lut (.I0(GND_net), .I1(n5061), .I2(n5086), .I3(n51390), 
            .O(n434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_9 (.CI(n51390), .I0(n5061), .I1(n5086), .CO(n51391));
    SB_LUT4 add_1091_8_lut (.I0(GND_net), .I1(n5062), .I2(n5087), .I3(n51389), 
            .O(n435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_8 (.CI(n51389), .I0(n5062), .I1(n5087), .CO(n51390));
    SB_LUT4 add_1091_7_lut (.I0(GND_net), .I1(n5063), .I2(n5088), .I3(n51388), 
            .O(n436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1836 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n57872));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1836.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1837 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n57871));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1837.LUT_INIT = 16'h2300;
    SB_CARRY add_1091_7 (.CI(n51388), .I0(n5063), .I1(n5088), .CO(n51389));
    SB_LUT4 add_1091_6_lut (.I0(GND_net), .I1(n5064), .I2(n5089), .I3(n51387), 
            .O(n437)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_6 (.CI(n51387), .I0(n5064), .I1(n5089), .CO(n51388));
    SB_LUT4 add_1091_5_lut (.I0(GND_net), .I1(n5065), .I2(n5090), .I3(n51386), 
            .O(n438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_5 (.CI(n51386), .I0(n5065), .I1(n5090), .CO(n51387));
    SB_LUT4 add_1091_4_lut (.I0(GND_net), .I1(n5066), .I2(n5091), .I3(n51385), 
            .O(n439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_4 (.CI(n51385), .I0(n5066), .I1(n5091), .CO(n51386));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1838 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n57994));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1838.LUT_INIT = 16'h2300;
    SB_LUT4 add_1091_3_lut (.I0(GND_net), .I1(n5067), .I2(n13_adj_5730), 
            .I3(n51384), .O(n440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1091_3 (.CI(n51384), .I0(n5067), .I1(n13_adj_5730), .CO(n51385));
    SB_LUT4 i1_3_lut_adj_1839 (.I0(control_mode[0]), .I1(n25130), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5725));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut_adj_1839.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_253_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5725), .I3(n15_adj_5732), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_253_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_1091_2_lut (.I0(GND_net), .I1(n5068), .I2(n5093), .I3(GND_net), 
            .O(n441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1091_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_251_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_91[23]), 
            .I2(n15_adj_5731), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_251_i24_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_1091_2 (.CI(GND_net), .I0(n5068), .I1(n5093), .CO(n51384));
    SB_LUT4 unary_minus_19_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n51383), .O(n330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n51382), .O(n334)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_14 (.CI(n51382), .I0(GND_net), .I1(n2), 
            .CO(n51383));
    SB_LUT4 unary_minus_19_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5707), 
            .I3(n51381), .O(n335)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_13 (.CI(n51381), .I0(GND_net), .I1(n14_adj_5707), 
            .CO(n51382));
    SB_LUT4 unary_minus_19_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5708), 
            .I3(n51380), .O(n336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_12 (.CI(n51380), .I0(GND_net), .I1(n15_adj_5708), 
            .CO(n51381));
    SB_LUT4 i13616_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n58142), .I3(GND_net), .O(n29359));   // verilog/coms.v(130[12] 305[6])
    defparam i13616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5709), 
            .I3(n51379), .O(n337)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_11 (.CI(n51379), .I0(GND_net), .I1(n16_adj_5709), 
            .CO(n51380));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n57870));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_19_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5710), 
            .I3(n51378), .O(n338)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_10 (.CI(n51378), .I0(GND_net), .I1(n17_adj_5710), 
            .CO(n51379));
    SB_LUT4 unary_minus_19_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5711), 
            .I3(n51377), .O(n339)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_9 (.CI(n51377), .I0(GND_net), .I1(n18_adj_5711), 
            .CO(n51378));
    SB_LUT4 unary_minus_19_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5712), 
            .I3(n51376), .O(n340)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_8 (.CI(n51376), .I0(GND_net), .I1(n19_adj_5712), 
            .CO(n51377));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n57869));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_19_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5713), 
            .I3(n51375), .O(n341)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_7 (.CI(n51375), .I0(GND_net), .I1(n20_adj_5713), 
            .CO(n51376));
    SB_LUT4 unary_minus_19_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5714), 
            .I3(n51374), .O(n342)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_6 (.CI(n51374), .I0(GND_net), .I1(n21_adj_5714), 
            .CO(n51375));
    SB_LUT4 unary_minus_19_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5715), 
            .I3(n51373), .O(n343)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_5 (.CI(n51373), .I0(GND_net), .I1(n22_adj_5715), 
            .CO(n51374));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1842 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n57868));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1842.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_19_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5716), 
            .I3(n51372), .O(n344)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_4 (.CI(n51372), .I0(GND_net), .I1(n23_adj_5716), 
            .CO(n51373));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n57867));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_19_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5717), 
            .I3(n51371), .O(n345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_3 (.CI(n51371), .I0(GND_net), .I1(n24_adj_5717), 
            .CO(n51372));
    SB_LUT4 unary_minus_19_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n25_adj_5718), 
            .I3(VCC_net), .O(n65385)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_19_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5718), 
            .CO(n51371));
    SB_LUT4 i13619_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n58142), .I3(GND_net), .O(n29362));   // verilog/coms.v(130[12] 305[6])
    defparam i13619_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5770), .I3(n51370), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5766), .I3(n51369), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n51369), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5766), .CO(n51370));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5765), .I3(n51368), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n51368), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5765), .CO(n51369));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5809), .I3(n51367), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n51367), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5809), .CO(n51368));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5808), .I3(n51366), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1844 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n57993));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1844.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n51366), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5808), .CO(n51367));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5807), .I3(n51365), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n51365), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5807), .CO(n51366));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5806), .I3(n51364), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n51364), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5806), .CO(n51365));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5805), .I3(n51363), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n51363), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5805), .CO(n51364));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5804), .I3(n51362), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n51362), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5804), .CO(n51363));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5802), .I3(n51361), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n51361), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5802), .CO(n51362));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5801), .I3(n51360), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1845 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n57992));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1845.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n51360), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5801), .CO(n51361));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5800), .I3(n51359), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n51359), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5800), .CO(n51360));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5799), .I3(n51358), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n51358), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5799), .CO(n51359));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5798), .I3(n51357), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n51357), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5798), .CO(n51358));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5785), .I3(n51356), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n51356), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5785), .CO(n51357));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5784), .I3(n51355), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n51355), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5784), .CO(n51356));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5783), .I3(n51354), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n51354), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5783), .CO(n51355));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5782), .I3(n51353), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n51353), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5782), .CO(n51354));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5781), .I3(n51352), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n51352), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5781), .CO(n51353));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5780), .I3(n51351), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49372_2_lut_4_lut (.I0(duty[8]), .I1(n338), .I2(duty[4]), 
            .I3(n342), .O(n66388));
    defparam i49372_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n51351), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5780), .CO(n51352));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5779), .I3(n51350), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n51350), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5779), .CO(n51351));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_5764), .I3(n51349), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n51349), .I0(GND_net), 
            .I1(n23_adj_5764), .CO(n51350));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_5763), .I3(n51348), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51066_4_lut (.I0(n16_adj_5687), .I1(n6_adj_5737), .I2(n19_adj_5685), 
            .I3(n66333), .O(n68082));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51066_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1846 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n57991));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1846.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1847 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n57990));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1847.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n28927));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1849 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n57989));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1849.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1850 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n57895));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1850.LUT_INIT = 16'h2300;
    SB_LUT4 i13301_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n27968), 
            .I3(GND_net), .O(n29044));   // verilog/coms.v(130[12] 305[6])
    defparam i13301_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1851 (.I0(\data_out_frame[8] [3]), .I1(n58828), 
            .I2(GND_net), .I3(GND_net), .O(n58312));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1851.LUT_INIT = 16'h6666;
    SB_LUT4 i51067_3_lut (.I0(n68082), .I1(current_limit[10]), .I2(n21), 
            .I3(GND_net), .O(n68083));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1852 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5724));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1852.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1853 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n57988));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1853.LUT_INIT = 16'h2300;
    SB_LUT4 i2_4_lut_adj_1854 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(\data_out_frame[15] [1]), .I3(n4_adj_5724), .O(n58925));   // verilog/coms.v(100[12:26])
    defparam i2_4_lut_adj_1854.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1855 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n57987));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1855.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n57866));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1857 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n57865));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1857.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n57864));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1859 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n57863));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1859.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1860 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n57862));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1860.LUT_INIT = 16'h2300;
    SB_LUT4 i13285_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n27968), 
            .I3(GND_net), .O(n29028));   // verilog/coms.v(130[12] 305[6])
    defparam i13285_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1861 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n57861));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1861.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1862 (.I0(\data_out_frame[6] [2]), .I1(n58238), 
            .I2(GND_net), .I3(GND_net), .O(n25237));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1862.LUT_INIT = 16'h6666;
    SB_LUT4 i50936_3_lut (.I0(n68083), .I1(current_limit[11]), .I2(n23), 
            .I3(GND_net), .O(n67952));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49207_3_lut (.I0(state_7__N_4108[0]), .I1(n38852), .I2(enable_slow_N_4211), 
            .I3(GND_net), .O(n65575));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i49207_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i16_4_lut (.I0(state_adj_5949[0]), .I1(n65575), .I2(n6388), 
            .I3(n6_adj_5846), .O(n8_adj_5860));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1863 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n57860));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1863.LUT_INIT = 16'h2300;
    SB_LUT4 i14_4_lut (.I0(duty[0]), .I1(duty[23]), .I2(duty[1]), .I3(duty[2]), 
            .O(n211));   // verilog/TinyFPGA_B.v(111[25:31])
    defparam i14_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i13904_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5918[0]), 
            .I2(n10_adj_5833), .I3(n25136), .O(n29647));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13904_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13281_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n27968), 
            .I3(GND_net), .O(n29024));   // verilog/coms.v(130[12] 305[6])
    defparam i13281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1864 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n57859));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1864.LUT_INIT = 16'h2300;
    SB_LUT4 i13924_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n61568), 
            .I3(n27), .O(n29667));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13924_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1865 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n57858));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1865.LUT_INIT = 16'h2300;
    SB_LUT4 i13940_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[0]), .I2(n11_adj_5758), 
            .I3(state_7__N_4317), .O(n29683));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13940_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13277_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n27968), 
            .I3(GND_net), .O(n29020));   // verilog/coms.v(130[12] 305[6])
    defparam i13277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1866 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n57857));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1866.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1867 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n57856));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1867.LUT_INIT = 16'h2300;
    SB_LUT4 i30_4_lut (.I0(state_7__N_3916[0]), .I1(n25014), .I2(state_adj_5919[1]), 
            .I3(n4_adj_5866), .O(n12_adj_5858));   // verilog/eeprom.v(35[8] 81[4])
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12_adj_5858), .I1(n65569), .I2(state_adj_5919[0]), 
            .I3(state_adj_5919[2]), .O(n57342));   // verilog/eeprom.v(35[8] 81[4])
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i13270_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n27968), 
            .I3(GND_net), .O(n29013));   // verilog/coms.v(130[12] 305[6])
    defparam i13270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13266_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n27968), 
            .I3(GND_net), .O(n29009));   // verilog/coms.v(130[12] 305[6])
    defparam i13266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n57855));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1869 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n28782));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1869.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1870 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n57854));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1870.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1871 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n28780));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1871.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1872 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n57853));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1872.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1873 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n57852));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1873.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1874 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58653));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1874.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1875 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n57986));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1875.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[6] [6]), .O(n58245));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n57985));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1877 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n57984));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1877.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_1878 (.I0(n38), .I1(n25996), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n58680));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1878.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n57983));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h2300;
    SB_LUT4 i14338_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3014));   // verilog/coms.v(130[12] 305[6])
    defparam i14338_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n57982));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n57981));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n57980));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n57979));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n57978));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h2300;
    SB_LUT4 i6_4_lut_adj_1885 (.I0(n58922), .I1(\data_out_frame[8] [7]), 
            .I2(n58245), .I3(n1130), .O(n14_adj_5797));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1885.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1886 (.I0(\data_out_frame[13] [2]), .I1(n14_adj_5797), 
            .I2(n10_adj_5811), .I3(\data_out_frame[10] [6]), .O(n25269));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut_adj_1886.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n57851));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n57977));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n57976));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h2300;
    SB_LUT4 i13992_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n22362), .I3(GND_net), .O(n29735));   // verilog/coms.v(130[12] 305[6])
    defparam i13992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n57975));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 i13993_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n22362), .I3(GND_net), .O(n29736));   // verilog/coms.v(130[12] 305[6])
    defparam i13993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13994_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n22362), .I3(GND_net), .O(n29737));   // verilog/coms.v(130[12] 305[6])
    defparam i13994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1891 (.I0(\data_in_frame[17] [6]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[6]), .O(n57370));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_1891.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13995_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n22362), .I3(GND_net), .O(n29738));   // verilog/coms.v(130[12] 305[6])
    defparam i13995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13996_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n22362), .I3(GND_net), .O(n29739));   // verilog/coms.v(130[12] 305[6])
    defparam i13996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13997_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n22362), .I3(GND_net), .O(n29740));   // verilog/coms.v(130[12] 305[6])
    defparam i13997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n57974));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h2300;
    SB_LUT4 i13999_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n22362), .I3(GND_net), .O(n29742));   // verilog/coms.v(130[12] 305[6])
    defparam i13999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n28909));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n57850));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h2300;
    SB_LUT4 i14000_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n22362), .I3(GND_net), .O(n29743));   // verilog/coms.v(130[12] 305[6])
    defparam i14000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13622_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n58142), .I3(GND_net), .O(n29365));   // verilog/coms.v(130[12] 305[6])
    defparam i13622_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14001_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n22362), .I3(GND_net), .O(n29744));   // verilog/coms.v(130[12] 305[6])
    defparam i14001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1895 (.I0(\data_in_frame[17] [5]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[5]), .O(n57372));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1895.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14002_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n22362), .I3(GND_net), .O(n29745));   // verilog/coms.v(130[12] 305[6])
    defparam i14002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14004_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n22362), .I3(GND_net), .O(n29747));   // verilog/coms.v(130[12] 305[6])
    defparam i14004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14005_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n22362), .I3(GND_net), .O(n29748));   // verilog/coms.v(130[12] 305[6])
    defparam i14005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14006_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n22362), .I3(GND_net), .O(n29749));   // verilog/coms.v(130[12] 305[6])
    defparam i14006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13625_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n58143), .I3(GND_net), .O(n29368));   // verilog/coms.v(130[12] 305[6])
    defparam i13625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1896 (.I0(\data_in_frame[17] [4]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[4]), .O(n57374));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1896.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13628_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n58143), .I3(GND_net), .O(n29371));   // verilog/coms.v(130[12] 305[6])
    defparam i13628_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1897 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58225));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1897.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n57849));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n57848));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n57847));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n28772));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i6_4_lut_adj_1902 (.I0(\data_out_frame[9] [1]), .I1(n26180), 
            .I2(n58225), .I3(\data_out_frame[11] [3]), .O(n14_adj_5831));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1902.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1903 (.I0(\data_out_frame[13] [5]), .I1(n14_adj_5831), 
            .I2(n10_adj_5832), .I3(n58644), .O(n58707));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut_adj_1903.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n57896));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n57846));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_LUT4 i13631_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n58143), .I3(GND_net), .O(n29374));   // verilog/coms.v(130[12] 305[6])
    defparam i13631_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1906 (.I0(\data_in_frame[17] [3]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[3]), .O(n57376));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1906.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n57845));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n28768));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_1909 (.I0(\data_out_frame[15] [2]), .I1(n53121), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n58321));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1909.LUT_INIT = 16'h9696;
    SB_LUT4 i13239_3_lut (.I0(\data_in_frame[2] [0]), .I1(rx_data[0]), .I2(n7_adj_5861), 
            .I3(GND_net), .O(n28982));   // verilog/coms.v(130[12] 305[6])
    defparam i13239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n28767));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1911 (.I0(\data_in_frame[17] [2]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[2]), .O(n57378));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1911.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n57844));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n57843));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1914 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58276));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1914.LUT_INIT = 16'h6666;
    SB_LUT4 i13773_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n27997), .I3(GND_net), .O(n29516));   // verilog/coms.v(130[12] 305[6])
    defparam i13773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n28764));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1916 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58742));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1916.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1917 (.I0(\data_out_frame[10] [0]), .I1(n58436), 
            .I2(\data_out_frame[10] [1]), .I3(\data_out_frame[9] [6]), .O(n12));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut_adj_1917.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1918 (.I0(\data_out_frame[7] [5]), .I1(n12), .I2(n58742), 
            .I3(\data_out_frame[5] [6]), .O(n1510));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1918.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n62_adj_5835), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_5834));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1919 (.I0(\data_out_frame[10] [5]), .I1(n58952), 
            .I2(GND_net), .I3(GND_net), .O(n58857));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1919.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n57842));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_1921 (.I0(\data_in_frame[17] [0]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[0]), .O(n57380));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1921.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_adj_1922 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58436));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1922.LUT_INIT = 16'h6666;
    SB_LUT4 n69008_bdd_4_lut (.I0(n69008), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n69011));
    defparam n69008_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51088_4_lut (.I0(current[15]), .I1(n23), .I2(current_limit[12]), 
            .I3(n67561), .O(n68104));
    defparam i51088_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i13767_3_lut (.I0(\data_in_frame[16] [7]), .I1(rx_data[7]), 
            .I2(n27994), .I3(GND_net), .O(n29510));   // verilog/coms.v(130[12] 305[6])
    defparam i13767_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13764_3_lut (.I0(\data_in_frame[16] [6]), .I1(rx_data[6]), 
            .I2(n27994), .I3(GND_net), .O(n29507));   // verilog/coms.v(130[12] 305[6])
    defparam i13764_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13634_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n58143), .I3(GND_net), .O(n29377));   // verilog/coms.v(130[12] 305[6])
    defparam i13634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13236_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n58147), 
            .I3(GND_net), .O(n28979));   // verilog/coms.v(130[12] 305[6])
    defparam i13236_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n57841));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_LUT4 i13233_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n58147), 
            .I3(GND_net), .O(n28976));   // verilog/coms.v(130[12] 305[6])
    defparam i13233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n57840));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 i13761_3_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(n27994), .I3(GND_net), .O(n29504));   // verilog/coms.v(130[12] 305[6])
    defparam i13761_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1925 (.I0(n58238), .I1(n58919), .I2(n58835), 
            .I3(n58632), .O(n60645));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1925.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1926 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(n60645), .I3(\data_out_frame[7] [6]), .O(n16_adj_5819));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1926.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1927 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[14] [5]), .I3(\data_out_frame[10] [5]), 
            .O(n17_adj_5818));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut_adj_1927.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1928 (.I0(n17_adj_5818), .I1(\data_out_frame[8] [4]), 
            .I2(n16_adj_5819), .I3(\data_out_frame[5] [6]), .O(n58608));   // verilog/coms.v(100[12:26])
    defparam i9_4_lut_adj_1928.LUT_INIT = 16'h6996;
    SB_LUT4 i51078_4_lut (.I0(n12_adj_5690), .I1(n4_adj_5738), .I2(n15_adj_5688), 
            .I3(n66342), .O(n68094));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51078_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13758_3_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(n27994), .I3(GND_net), .O(n29501));   // verilog/coms.v(130[12] 305[6])
    defparam i13758_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13229_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n58147), 
            .I3(GND_net), .O(n28972));   // verilog/coms.v(130[12] 305[6])
    defparam i13229_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n57839));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h2300;
    SB_LUT4 i13637_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n58143), .I3(GND_net), .O(n29380));   // verilog/coms.v(130[12] 305[6])
    defparam i13637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13226_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n58147), 
            .I3(GND_net), .O(n28969));   // verilog/coms.v(130[12] 305[6])
    defparam i13226_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [5]), .O(n58952));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n57838));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h2300;
    SB_LUT4 i13755_3_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(n27994), .I3(GND_net), .O(n29498));   // verilog/coms.v(130[12] 305[6])
    defparam i13755_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1931 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n57837));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1931.LUT_INIT = 16'h2300;
    SB_LUT4 i13640_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n58143), .I3(GND_net), .O(n29383));   // verilog/coms.v(130[12] 305[6])
    defparam i13640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13698_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n58145), .I3(GND_net), .O(n29441));   // verilog/coms.v(130[12] 305[6])
    defparam i13698_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13752_3_lut (.I0(\data_in_frame[16] [2]), .I1(rx_data[2]), 
            .I2(n27994), .I3(GND_net), .O(n29495));   // verilog/coms.v(130[12] 305[6])
    defparam i13752_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n57836));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n57835));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n57973));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n57834));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n57972));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n57971));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n57970));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n10_adj_5811));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n57969));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n57968));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_LUT4 i13743_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n58139), .I3(GND_net), .O(n29486));   // verilog/coms.v(130[12] 305[6])
    defparam i13743_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1941 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n57967));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1941.LUT_INIT = 16'h2300;
    SB_LUT4 i49363_2_lut_3_lut (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(state_adj_5919[1]), .I3(GND_net), .O(n65569));   // verilog/eeprom.v(35[8] 81[4])
    defparam i49363_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1942 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n57966));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1942.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n57965));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 i50307_3_lut (.I0(n67952), .I1(current_limit[12]), .I2(current[15]), 
            .I3(GND_net), .O(n67323));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50307_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n57964));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n57963));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n57832));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n57962));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n57961));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_4_lut_adj_1949 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n38797), .O(n56676));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_4_lut_4_lut_adj_1949.LUT_INIT = 16'hb1f1;
    SB_LUT4 i13643_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n58143), .I3(GND_net), .O(n29386));   // verilog/coms.v(130[12] 305[6])
    defparam i13643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n57960));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n57959));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_LUT4 i51213_3_lut (.I0(n67323), .I1(n68094), .I2(n68104), .I3(GND_net), 
            .O(n68229));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n57958));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i13646_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n58143), .I3(GND_net), .O(n29389));   // verilog/coms.v(130[12] 305[6])
    defparam i13646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n57957));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 i51117_4_lut (.I0(n68229), .I1(current_limit[14]), .I2(current[15]), 
            .I3(current_limit[13]), .O(n30));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51117_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n58003));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n58002));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n58001));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n58000));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n57999));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n57998));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n57997));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_LUT4 i13701_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n58145), .I3(GND_net), .O(n29444));   // verilog/coms.v(130[12] 305[6])
    defparam i13701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n57956));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 i13704_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n58145), .I3(GND_net), .O(n29447));   // verilog/coms.v(130[12] 305[6])
    defparam i13704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n57955));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i13649_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n58144), .I3(GND_net), .O(n29392));   // verilog/coms.v(130[12] 305[6])
    defparam i13649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13707_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n58145), .I3(GND_net), .O(n29450));   // verilog/coms.v(130[12] 305[6])
    defparam i13707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n26_adj_5844));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n57954));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 i13710_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n58145), .I3(GND_net), .O(n29453));   // verilog/coms.v(130[12] 305[6])
    defparam i13710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n57953));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 i13713_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n58145), .I3(GND_net), .O(n29456));   // verilog/coms.v(130[12] 305[6])
    defparam i13713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13652_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n58144), .I3(GND_net), .O(n29395));   // verilog/coms.v(130[12] 305[6])
    defparam i13652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n57952));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_20_i5_2_lut (.I0(duty[2]), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49435_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n66451));
    defparam i49435_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n57951));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n342), .I1(n338), .I2(n17), .I3(GND_net), 
            .O(n8));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n57950));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_20_i6_3_lut (.I0(n344), .I1(n343), .I2(n7), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i16_3_lut (.I0(n8), .I1(n337), .I2(n19), .I3(GND_net), 
            .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n57949));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i45524_3_lut (.I0(duty[19]), .I1(duty[21]), .I2(n330), .I3(GND_net), 
            .O(n62531));
    defparam i45524_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i13656_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n58144), .I3(GND_net), .O(n29399));   // verilog/coms.v(130[12] 305[6])
    defparam i13656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i45528_3_lut (.I0(duty[14]), .I1(duty[17]), .I2(n330), .I3(GND_net), 
            .O(n62535));
    defparam i45528_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i13716_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n58145), .I3(GND_net), .O(n29459));   // verilog/coms.v(130[12] 305[6])
    defparam i13716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i45642_4_lut (.I0(duty[20]), .I1(n62531), .I2(duty[22]), .I3(n330), 
            .O(n62649));
    defparam i45642_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 LessThan_20_i4_3_lut (.I0(n65385), .I1(n345), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n68918_bdd_4_lut (.I0(n68918), .I1(duty[18]), .I2(n252), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[18]));
    defparam n68918_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50853_3_lut (.I0(n4), .I1(n341), .I2(n11), .I3(GND_net), 
            .O(n67869));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i50853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n57948));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i13659_3_lut (.I0(\data_in_frame[12] [3]), .I1(rx_data[3]), 
            .I2(n58144), .I3(GND_net), .O(n29402));   // verilog/coms.v(130[12] 305[6])
    defparam i13659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n57947));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i50854_3_lut (.I0(n67869), .I1(n340), .I2(n13), .I3(GND_net), 
            .O(n67870));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i50854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n57946));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n57945));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n57944));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n57943));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n57942));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n57941));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n57940));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 i49384_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n66451), 
            .O(n66400));
    defparam i49384_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5763));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n57939));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 i51082_4_lut (.I0(n16), .I1(n6), .I2(n19), .I3(n66388), 
            .O(n68098));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51082_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13719_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n58145), .I3(GND_net), .O(n29462));   // verilog/coms.v(130[12] 305[6])
    defparam i13719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n57938));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n57937));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n57936));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n57935));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n57934));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i13722_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n58139), .I3(GND_net), .O(n29465));   // verilog/coms.v(130[12] 305[6])
    defparam i13722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49576_3_lut (.I0(n67870), .I1(n339), .I2(n15), .I3(GND_net), 
            .O(n66592));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i49576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51286_4_lut (.I0(n66592), .I1(n68098), .I2(n19), .I3(n66400), 
            .O(n68302));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51286_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n57933));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n57932));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n57931));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n57930));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n57929));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n57928));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n57927));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n57926));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_1993 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_3_lut_adj_1993.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n57925));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n57924));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_5869));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1996 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1996.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n57923));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i13662_3_lut (.I0(\data_in_frame[12] [4]), .I1(rx_data[4]), 
            .I2(n58144), .I3(GND_net), .O(n29405));   // verilog/coms.v(130[12] 305[6])
    defparam i13662_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n57922));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h2300;
    SB_LUT4 i51287_3_lut (.I0(n68302), .I1(n336), .I2(duty[10]), .I3(GND_net), 
            .O(n68303));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51287_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n57921));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 i51212_3_lut (.I0(n68303), .I1(n335), .I2(duty[11]), .I3(GND_net), 
            .O(n68228));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51212_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n57920));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5737));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n57919));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 i23439_2_lut_2_lut (.I0(duty[23]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5070));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23439_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23440_2_lut_2_lut (.I0(duty[22]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5071));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23440_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13665_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n58144), .I3(GND_net), .O(n29408));   // verilog/coms.v(130[12] 305[6])
    defparam i13665_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13668_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n58144), .I3(GND_net), .O(n29411));   // verilog/coms.v(130[12] 305[6])
    defparam i13668_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23441_2_lut_2_lut (.I0(duty[21]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5072));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23441_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23442_2_lut_2_lut (.I0(duty[20]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5073));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23442_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23443_2_lut_2_lut (.I0(duty[19]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5074));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23443_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n57918));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n57917));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i23444_2_lut_2_lut (.I0(duty[18]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5075));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23444_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23445_2_lut_2_lut (.I0(duty[17]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5076));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23445_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23446_2_lut_2_lut (.I0(duty[16]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5077));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23446_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23447_2_lut_2_lut (.I0(duty[15]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5078));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23447_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23448_2_lut_2_lut (.I0(duty[14]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5079));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23448_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 LessThan_20_i26_3_lut (.I0(n68228), .I1(n334), .I2(duty[12]), 
            .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i23452_2_lut_2_lut (.I0(duty[13]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5080));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23452_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23453_2_lut_2_lut (.I0(duty[12]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5081));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23453_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23454_2_lut_2_lut (.I0(duty[11]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5082));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23454_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23455_2_lut_2_lut (.I0(duty[10]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5083));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23455_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23456_2_lut_2_lut (.I0(duty[9]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5084));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23456_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23457_2_lut_2_lut (.I0(duty[8]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5085));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23457_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13671_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n58144), .I3(GND_net), .O(n29414));   // verilog/coms.v(130[12] 305[6])
    defparam i13671_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23458_2_lut_2_lut (.I0(duty[7]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5086));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23458_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12668_2_lut (.I0(n27211), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28417));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i12668_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13674_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n60939), .I3(GND_net), .O(n29417));   // verilog/coms.v(130[12] 305[6])
    defparam i13674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51340_4_lut (.I0(commutation_state[1]), .I1(n22497), .I2(dti), 
            .I3(commutation_state[2]), .O(n27211));
    defparam i51340_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i13677_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n60939), .I3(GND_net), .O(n29420));   // verilog/coms.v(130[12] 305[6])
    defparam i13677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23459_2_lut_2_lut (.I0(duty[6]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5087));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23459_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23460_2_lut_2_lut (.I0(duty[5]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5088));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23460_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i13273_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n22373), .I3(GND_net), .O(n29016));   // verilog/coms.v(130[12] 305[6])
    defparam i13273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23461_2_lut_2_lut (.I0(duty[4]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5089));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23461_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23462_2_lut_2_lut (.I0(duty[3]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5090));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23462_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i48767_2_lut (.I0(n68699), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65592));
    defparam i48767_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i23463_2_lut_2_lut (.I0(duty[2]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5091));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i23463_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7_4_lut_adj_2004 (.I0(duty[18]), .I1(n26), .I2(n330), .I3(duty[23]), 
            .O(n20_adj_5813));
    defparam i7_4_lut_adj_2004.LUT_INIT = 16'h2100;
    SB_LUT4 i50411_3_lut (.I0(n68969), .I1(n68795), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67427));
    defparam i50411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_2_lut_adj_2005 (.I0(n296), .I1(duty[1]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5730));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_2_lut_2_lut_adj_2005.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n57916));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n57915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 i13725_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n58139), .I3(GND_net), .O(n29468));   // verilog/coms.v(130[12] 305[6])
    defparam i13725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n57914));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 i11_4_lut (.I0(n330), .I1(n62649), .I2(n62535), .I3(duty[13]), 
            .O(n24_adj_5812));
    defparam i11_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n57913));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n57912));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 i13680_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n60939), .I3(GND_net), .O(n29423));   // verilog/coms.v(130[12] 305[6])
    defparam i13680_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13728_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n58139), .I3(GND_net), .O(n29471));   // verilog/coms.v(130[12] 305[6])
    defparam i13728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n57911));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n57898));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h2300;
    SB_LUT4 i13683_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n60939), .I3(GND_net), .O(n29426));   // verilog/coms.v(130[12] 305[6])
    defparam i13683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n57910));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 i48940_4_lut (.I0(duty[16]), .I1(n20_adj_5813), .I2(duty[15]), 
            .I3(n330), .O(n65556));
    defparam i48940_4_lut.LUT_INIT = 16'h8004;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n57909));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n57908));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 i14_4_lut_adj_2016 (.I0(n65556), .I1(pwm_setpoint_23__N_207), 
            .I2(n296), .I3(n24_adj_5812), .O(n9618));
    defparam i14_4_lut_adj_2016.LUT_INIT = 16'hcac0;
    SB_LUT4 i49317_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n66333));
    defparam i49317_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n57897));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5735));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2018 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n28838));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2018.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2019 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n28837));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2019.LUT_INIT = 16'h2300;
    SB_LUT4 i13731_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n58139), .I3(GND_net), .O(n29474));   // verilog/coms.v(130[12] 305[6])
    defparam i13731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2020 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n57907));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2020.LUT_INIT = 16'h2300;
    SB_LUT4 i13274_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n22362), .I3(GND_net), .O(n29017));   // verilog/coms.v(130[12] 305[6])
    defparam i13274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2021 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n57906));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2021.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n57904));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2023 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n57905));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2023.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2024 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n57833));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2024.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2025 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n28831));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2025.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2026 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n57903));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2026.LUT_INIT = 16'h2300;
    SB_LUT4 i10_1_lut_adj_2027 (.I0(duty[23]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut_adj_2027.LUT_INIT = 16'h5555;
    SB_LUT4 i13275_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n22362), .I3(GND_net), .O(n29018));   // verilog/coms.v(130[12] 305[6])
    defparam i13275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n57902));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2029 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n57901));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2029.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n28827));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2031 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n57900));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2031.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n28825));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2033 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n57899));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2033.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2034 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n57891));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2034.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2035 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n57890));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2035.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n57889));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h2300;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51916 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n68990));
    defparam byte_transmit_counter_0__bdd_4_lut_51916.LUT_INIT = 16'he4aa;
    SB_LUT4 n68990_bdd_4_lut (.I0(n68990), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n68993));
    defparam n68990_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5227_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5227_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i13737_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n58139), .I3(GND_net), .O(n29480));   // verilog/coms.v(130[12] 305[6])
    defparam i13737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5225_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5225_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2037 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n57888));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2037.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n57887));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h2300;
    SB_LUT4 i1848_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1405), .I3(n38797), .O(n6579));   // verilog/TinyFPGA_B.v(361[5] 387[12])
    defparam i1848_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i49326_2_lut_4_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(current[5]), .I3(current_limit[5]), .O(n66342));
    defparam i49326_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i13501_4_lut_4_lut (.I0(n27429), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n29244));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13501_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 i13280_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(control_update), .I3(GND_net), .O(n29023));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i10_3_lut_3_lut (.I0(current_limit[5]), .I1(current_limit[6]), 
            .I2(current[6]), .I3(GND_net), .O(n10_adj_5733));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n9618_bdd_4_lut_51677 (.I0(n9618), .I1(n436), .I2(current[5]), 
            .I3(duty[23]), .O(n68702));
    defparam n9618_bdd_4_lut_51677.LUT_INIT = 16'he4aa;
    SB_LUT4 n68702_bdd_4_lut (.I0(n68702), .I1(duty[5]), .I2(n265), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n68702_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n58922));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_2039 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n58238));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_2039.LUT_INIT = 16'h9696;
    SB_LUT4 unary_minus_18_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5706));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5743));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_2040 (.I0(state_adj_5919[2]), .I1(data_ready), 
            .I2(n39313), .I3(n25133), .O(n57558));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_2040.LUT_INIT = 16'hcca8;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5740));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5744));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5741));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5748));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5746));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5745));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i5_2_lut (.I0(current[2]), .I1(duty[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5750));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49078_4_lut (.I0(n11_adj_5745), .I1(n9_adj_5746), .I2(n7_adj_5748), 
            .I3(n5_adj_5750), .O(n66094));
    defparam i49078_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13289_3_lut (.I0(current[0]), .I1(data_adj_5926[0]), .I2(n27270), 
            .I3(GND_net), .O(n29032));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5747), .I1(duty[9]), .I2(n19_adj_5740), 
            .I3(GND_net), .O(n16_adj_5742));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50843_3_lut (.I0(n4_adj_5751), .I1(duty[5]), .I2(n11_adj_5745), 
            .I3(GND_net), .O(n67859));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50844_3_lut (.I0(n67859), .I1(duty[6]), .I2(n13_adj_5744), 
            .I3(GND_net), .O(n67860));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49044_4_lut (.I0(n17_adj_5741), .I1(n15_adj_5743), .I2(n13_adj_5744), 
            .I3(n66094), .O(n66060));
    defparam i49044_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51048_4_lut (.I0(n16_adj_5742), .I1(n6_adj_5749), .I2(n19_adj_5740), 
            .I3(n66058), .O(n68064));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51048_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i23149_2_lut (.I0(n22497), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n38795));
    defparam i23149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49596_3_lut (.I0(n67860), .I1(duty[7]), .I2(n15_adj_5743), 
            .I3(GND_net), .O(n66612));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i49596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51272_4_lut (.I0(n66612), .I1(n68064), .I2(n19_adj_5740), 
            .I3(n66060), .O(n68288));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51272_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51273_3_lut (.I0(n68288), .I1(duty[10]), .I2(current[10]), 
            .I3(GND_net), .O(n68289));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51273_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_2041 (.I0(control_mode[0]), .I1(n25130), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_5731));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_3_lut_adj_2041.LUT_INIT = 16'hfefe;
    SB_LUT4 i51218_3_lut (.I0(n68289), .I1(duty[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5739));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51218_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_2042 (.I0(control_mode[0]), .I1(n25130), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_5732));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_3_lut_adj_2042.LUT_INIT = 16'hefef;
    SB_LUT4 i3_4_lut_adj_2043 (.I0(duty[14]), .I1(n24_adj_5739), .I2(duty[12]), 
            .I3(duty[13]), .O(n59821));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_2043.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_2044 (.I0(duty[14]), .I1(n24_adj_5739), .I2(duty[12]), 
            .I3(duty[13]), .O(n59823));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_2044.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_2045 (.I0(duty[15]), .I1(current[15]), .I2(n59823), 
            .I3(n59821), .O(n32));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_2045.LUT_INIT = 16'hb3a2;
    SB_LUT4 i3_4_lut_adj_2046 (.I0(duty[18]), .I1(n32), .I2(duty[16]), 
            .I3(duty[17]), .O(n59843));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_2046.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_2047 (.I0(duty[18]), .I1(n32), .I2(duty[16]), 
            .I3(duty[17]), .O(n59845));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_2047.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_2048 (.I0(duty[19]), .I1(current[15]), .I2(n59845), 
            .I3(n59843), .O(n40));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_2048.LUT_INIT = 16'hb3a2;
    SB_LUT4 i3_4_lut_adj_2049 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n59877));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_2049.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_2050 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n59879));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_2050.LUT_INIT = 16'h8000;
    SB_LUT4 i13686_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n60939), .I3(GND_net), .O(n29429));   // verilog/coms.v(130[12] 305[6])
    defparam i13686_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49430_2_lut (.I0(n68633), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65590));
    defparam i49430_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50413_3_lut (.I0(n69011), .I1(n68789), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67429));
    defparam i50413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5705));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13290_4_lut (.I0(rw), .I1(state_adj_5919[1]), .I2(state_adj_5919[2]), 
            .I3(n5754), .O(n29033));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13290_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 unary_minus_18_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27288), .O(n54370));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 n9618_bdd_4_lut_51667 (.I0(n9618), .I1(n437), .I2(current[4]), 
            .I3(duty[23]), .O(n68684));
    defparam n9618_bdd_4_lut_51667.LUT_INIT = 16'he4aa;
    SB_LUT4 n68684_bdd_4_lut (.I0(n68684), .I1(duty[4]), .I2(n266), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n68684_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51906 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n68966));
    defparam byte_transmit_counter_0__bdd_4_lut_51906.LUT_INIT = 16'he4aa;
    SB_LUT4 i13296_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(n58096), .I3(state_7__N_4108[0]), 
            .O(n29039));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13296_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 n68966_bdd_4_lut (.I0(n68966), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n68969));
    defparam n68966_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_2051 (.I0(hall1), .I1(commutation_state[2]), .I2(hall3), 
            .I3(hall2), .O(n57628));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_2051.LUT_INIT = 16'hd054;
    SB_LUT4 unary_minus_18_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5704));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13300_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n25_adj_5857), .I3(GND_net), .O(n29043));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13300_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_2052 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n60966));
    defparam i3_4_lut_adj_2052.LUT_INIT = 16'h0004;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5842));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i1_2_lut_4_lut_adj_2053 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1405), .I3(n38797), .O(n24_adj_5853));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_adj_2053.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_4_lut_4_lut_adj_2054 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2961), .O(n25_adj_5852));   // verilog/TinyFPGA_B.v(376[7:11])
    defparam i1_4_lut_4_lut_adj_2054.LUT_INIT = 16'h5450;
    SB_LUT4 i13689_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n60939), .I3(GND_net), .O(n29432));   // verilog/coms.v(130[12] 305[6])
    defparam i13689_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13734_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n58139), .I3(GND_net), .O(n29477));   // verilog/coms.v(130[12] 305[6])
    defparam i13734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9618_bdd_4_lut_51846 (.I0(n9618), .I1(n424), .I2(current[15]), 
            .I3(duty[23]), .O(n68912));
    defparam n9618_bdd_4_lut_51846.LUT_INIT = 16'he4aa;
    SB_LUT4 n68912_bdd_4_lut (.I0(n68912), .I1(duty[17]), .I2(n253), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[17]));
    defparam n68912_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_18_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5703));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5702));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51886 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n68960));
    defparam byte_transmit_counter_0__bdd_4_lut_51886.LUT_INIT = 16'he4aa;
    SB_LUT4 n68960_bdd_4_lut (.I0(n68960), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n68963));
    defparam n68960_bdd_4_lut.LUT_INIT = 16'haad8;
    \quadrature_decoder(1)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1928(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .n1883(n1883), 
            .GND_net(GND_net), .n1885(n1885), .n1887(n1887), .n1889(n1889), 
            .n1891(n1891), .n1893(n1893), .n1895(n1895), .n1897(n1897), 
            .n1899(n1899), .n1901(n1901), .n1903(n1903), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net), .\a_new[1] (a_new[1]), .position_31__N_3827(position_31__N_3827), 
            .b_prev(b_prev), .n29053(n29053), .n1881(n1881)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(304[49] 310[6])
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    \quadrature_decoder(1)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1928(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .\a_new[1] (a_new_adj_5905[1]), 
            .position_31__N_3827(position_31__N_3827_adj_5761), .n29051(n29051), 
            .n1933(n1933), .b_prev(b_prev_adj_5760)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[49] 318[6])
    SB_LUT4 n68900_bdd_4_lut (.I0(n68900), .I1(duty[15]), .I2(n255), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[15]));
    defparam n68900_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51657 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(byte_transmit_counter[1]), .O(n68642));
    defparam byte_transmit_counter_0__bdd_4_lut_51657.LUT_INIT = 16'he4aa;
    SB_LUT4 n68642_bdd_4_lut (.I0(n68642), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(byte_transmit_counter[1]), 
            .O(n68645));
    defparam n68642_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51931 (.I0(n9618), .I1(n418), .I2(current[15]), 
            .I3(duty[23]), .O(n68948));
    defparam n9618_bdd_4_lut_51931.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_3_lut_4_lut (.I0(\data_in_frame[8] [1]), .I1(n58867), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[3] [6]), .O(n11_adj_5864));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n68948_bdd_3_lut (.I0(n68948), .I1(duty[23]), .I2(n249), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam n68948_bdd_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 i48800_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n65488));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48800_2_lut_4_lut.LUT_INIT = 16'h2100;
    TLI4970 tli (.GND_net(GND_net), .VCC_net(VCC_net), .clk16MHz(clk16MHz), 
            .n27270(n27270), .\current[15] (current[15]), .state_7__N_4317(state_7__N_4317), 
            .n6(n6_adj_5756), .n5(n5_adj_5757), .n5_adj_23(n5_adj_5755), 
            .n6_adj_24(n6_adj_5754), .n29103(n29103), .\current[1] (current[1]), 
            .n29102(n29102), .\current[2] (current[2]), .n29101(n29101), 
            .\current[3] (current[3]), .n29100(n29100), .\current[4] (current[4]), 
            .n29099(n29099), .\current[5] (current[5]), .n29098(n29098), 
            .\current[6] (current[6]), .n29097(n29097), .\current[7] (current[7]), 
            .n29096(n29096), .\current[8] (current[8]), .n29095(n29095), 
            .\current[9] (current[9]), .n29094(n29094), .\current[10] (current[10]), 
            .n29093(n29093), .\current[11] (current[11]), .n38922(n38922), 
            .CS_c(CS_c), .n29032(n29032), .\current[0] (current[0]), .n11(n11_adj_5758), 
            .CS_CLK_c(CS_CLK_c), .n29904(n29904), .\data[15] (data_adj_5926[15]), 
            .n29903(n29903), .\data[12] (data_adj_5926[12]), .n29902(n29902), 
            .\data[11] (data_adj_5926[11]), .n29901(n29901), .\data[10] (data_adj_5926[10]), 
            .n29900(n29900), .\data[9] (data_adj_5926[9]), .n29899(n29899), 
            .\data[8] (data_adj_5926[8]), .n29898(n29898), .\data[7] (data_adj_5926[7]), 
            .n29897(n29897), .\data[6] (data_adj_5926[6]), .n29896(n29896), 
            .\data[5] (data_adj_5926[5]), .n29895(n29895), .\data[4] (data_adj_5926[4]), 
            .n29894(n29894), .\data[3] (data_adj_5926[3]), .n29893(n29893), 
            .\data[2] (data_adj_5926[2]), .n29892(n29892), .\data[1] (data_adj_5926[1]), 
            .n29683(n29683), .\data[0] (data_adj_5926[0]), .\duty[0] (duty[0]), 
            .\duty[1] (duty[1]), .n4(n4_adj_5751), .n25112(n25112), .n25151(n25151), 
            .n25141(n25141), .n25145(n25145), .n25148(n25148), .n6_adj_25(n6_adj_5726), 
            .n5_adj_26(n5_adj_5810)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(404[11] 410[4])
    SB_LUT4 i49261_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n65531));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i49261_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i48745_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n65532));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48745_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i48698_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n65533));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48698_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 n9618_bdd_4_lut_51652 (.I0(n9618), .I1(n438), .I2(current[3]), 
            .I3(duty[23]), .O(n68624));
    defparam n9618_bdd_4_lut_51652.LUT_INIT = 16'he4aa;
    SB_LUT4 n68624_bdd_4_lut (.I0(n68624), .I1(duty[3]), .I2(n267), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n68624_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9618_bdd_4_lut_51871 (.I0(n9618), .I1(n419), .I2(current[15]), 
            .I3(duty[23]), .O(n68942));
    defparam n9618_bdd_4_lut_51871.LUT_INIT = 16'he4aa;
    SB_LUT4 n68942_bdd_4_lut (.I0(n68942), .I1(duty[22]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam n68942_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48844_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n65534));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48844_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i48744_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n65535));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48744_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i48743_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n65536));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48743_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i48742_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n65537));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i48742_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_4_lut_adj_2055 (.I0(commutation_state[0]), .I1(n4_adj_5729), 
            .I2(commutation_state_prev[0]), .I3(dti_N_404), .O(n27187));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_2055.LUT_INIT = 16'hdeff;
    coms neopxl_color_23__I_0 (.\data_in_frame[5] ({Open_0, Open_1, Open_2, 
         \data_in_frame[5] [4], Open_3, Open_4, \data_in_frame[5] [1], 
         Open_5}), .n3014(n3014), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .clk16MHz(clk16MHz), .n57886(n57886), .n58004(n58004), .n29483(n29483), 
         .VCC_net(VCC_net), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .n57892(n57892), .n57893(n57893), .n57885(n57885), .n29480(n29480), 
         .n57884(n57884), .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[2] ({Open_6, 
         Open_7, Open_8, Open_9, Open_10, Open_11, \data_in_frame[2] [1:0]}), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .n57894(n57894), .n57883(n57883), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n57882(n57882), 
         .n57881(n57881), .n57880(n57880), .n57879(n57879), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .GND_net(GND_net), .\data_in_frame[3] ({Open_12, \data_in_frame[3] [6], 
         Open_13, Open_14, Open_15, Open_16, \data_in_frame[3] [1], 
         Open_17}), .n57878(n57878), .\data_out_frame[1][6] (\data_out_frame[1] [6]), 
         .n57996(n57996), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .n57995(n57995), .n57877(n57877), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), 
         .pwm_setpoint({pwm_setpoint}), .n57876(n57876), .n57875(n57875), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n57874(n57874), 
         .n57873(n57873), .n25488(n25488), .n57872(n57872), .n57871(n57871), 
         .\data_in_frame[14] ({\data_in_frame[14] }), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .n29477(n29477), .Kp_23__N_869(Kp_23__N_869), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n57994(n57994), .n57870(n57870), .n57869(n57869), .n58867(n58867), 
         .n58698(n58698), .n53862(n53862), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n57868(n57868), .n57867(n57867), .\data_out_frame[3][3] (\data_out_frame[3] [3]), 
         .n57993(n57993), .\data_in_frame[2][5] (\data_in_frame[2] [5]), 
         .n29474(n29474), .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .n57992(n57992), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .n57991(n57991), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n57990(n57990), 
         .\data_in_frame[3][4] (\data_in_frame[3] [4]), .n29471(n29471), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .n28927(n28927), .n57989(n57989), 
         .n57895(n57895), .\data_in_frame[5][6] (\data_in_frame[5] [6]), 
         .n29468(n29468), .n57988(n57988), .n57987(n57987), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n57866(n57866), .n57865(n57865), .n57864(n57864), .n57863(n57863), 
         .n57862(n57862), .n57861(n57861), .n57860(n57860), .n57859(n57859), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .n57858(n57858), 
         .n57857(n57857), .n57856(n57856), .n57855(n57855), .n28782(n28782), 
         .n57854(n57854), .n28780(n28780), .n57853(n57853), .n57852(n57852), 
         .n57986(n57986), .n29465(n29465), .n57985(n57985), .n62(n62_adj_5835), 
         .n57984(n57984), .\data_out_frame[5] ({\data_out_frame[5] }), .n57983(n57983), 
         .n29462(n29462), .n57982(n57982), .n57981(n57981), .n57980(n57980), 
         .n29459(n29459), .n57979(n57979), .n57978(n57978), .n57851(n57851), 
         .n29456(n29456), .n57977(n57977), .n29453(n29453), .n57976(n57976), 
         .n29450(n29450), .\data_out_frame[6] ({\data_out_frame[6] }), .\encoder0_position_scaled[22] (encoder0_position_scaled[22]), 
         .n57975(n57975), .n29447(n29447), .n57974(n57974), .n29444(n29444), 
         .n28909(n28909), .n57850(n57850), .n57849(n57849), .n57848(n57848), 
         .n57847(n57847), .n28772(n28772), .n57896(n57896), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n57846(n57846), .n57845(n57845), .n28768(n28768), .n28767(n28767), 
         .n57844(n57844), .n57843(n57843), .n28764(n28764), .n57842(n57842), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .n57841(n57841), 
         .n57840(n57840), .n57839(n57839), .n57838(n57838), .n57837(n57837), 
         .n57836(n57836), .n57835(n57835), .n57973(n57973), .n29441(n29441), 
         .n57834(n57834), .neopxl_color({neopxl_color}), .n22373(n22373), 
         .n58391(n58391), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .\data_in_frame[5][3] (\data_in_frame[5] [3]), .n11(n11_adj_5864), 
         .n12(n12_adj_5863), .\data_in_frame[20] ({Open_18, Open_19, Open_20, 
         \data_in_frame[20] [4:2], Open_21, Open_22}), .n29438(n29438), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[21] ({\data_in_frame[21] [7:4], 
         Open_23, \data_in_frame[21] [2:0]}), .\data_in_frame[23][2] (\data_in_frame[23] [2]), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_in_frame[23][6] (\data_in_frame[23] [6]), .\data_in_frame[16] ({Open_24, 
         \data_in_frame[16] [6], Open_25, Open_26, \data_in_frame[16] [3:2], 
         Open_27, Open_28}), .\data_in_frame[20][1] (\data_in_frame[20] [1]), 
         .n57972(n57972), .\data_in_frame[3][0] (\data_in_frame[3] [0]), 
         .\data_in_frame[5][2] (\data_in_frame[5] [2]), .n57971(n57971), 
         .\data_in_frame[23][1] (\data_in_frame[23] [1]), .\data_in_frame[23][7] (\data_in_frame[23] [7]), 
         .\data_in_frame[23][0] (\data_in_frame[23] [0]), .\data_in_frame[20][5] (\data_in_frame[20] [5]), 
         .reset(reset), .\data_in_frame[5][0] (\data_in_frame[5] [0]), .n29435(n29435), 
         .setpoint({setpoint}), .\data_in_frame[20][6] (\data_in_frame[20] [6]), 
         .byte_transmit_counter({Open_29, Open_30, Open_31, byte_transmit_counter[4:1], 
         Open_32}), .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[3][2] (\data_in_frame[3] [2]), 
         .n57970(n57970), .\data_in_frame[16][5] (\data_in_frame[16] [5]), 
         .\data_in_frame[16][4] (\data_in_frame[16] [4]), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .n29432(n29432), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_in_frame[17] ({Open_33, 
         \data_in_frame[17] [6:1], Open_34}), .n29429(n29429), .n57969(n57969), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .n29426(n29426), 
         .n57968(n57968), .n29423(n29423), .n57967(n57967), .rx_data({rx_data}), 
         .n7(n7_adj_5861), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n29420(n29420), .n29417(n29417), .n29414(n29414), .n57966(n57966), 
         .n29411(n29411), .n29408(n29408), .n29405(n29405), .n68861(n68861), 
         .n68855(n68855), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n29402(n29402), .n57965(n57965), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .displacement({displacement}), .\encoder0_position_scaled[21] (encoder0_position_scaled[21]), 
         .n29399(n29399), .\data_in_frame[17][0] (\data_in_frame[17] [0]), 
         .PWMLimit({PWMLimit}), .n29395(n29395), .n57964(n57964), .n29392(n29392), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .encoder1_position_scaled({encoder1_position_scaled}), 
         .n29389(n29389), .n29386(n29386), .n27924(n27924), .\data_in_frame[16][7] (\data_in_frame[16] [7]), 
         .n28009(n28009), .n29383(n29383), .n29380(n29380), .n68849(n68849), 
         .n29377(n29377), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n29374(n29374), .\encoder0_position_scaled[20] (encoder0_position_scaled[20]), 
         .n29371(n29371), .n29368(n29368), .n29365(n29365), .n29362(n29362), 
         .n29359(n29359), .\data_out_frame[9] ({\data_out_frame[9] }), .n57963(n57963), 
         .n29356(n29356), .n29353(n29353), .n29350(n29350), .n29347(n29347), 
         .n29344(n29344), .n29341(n29341), .n29338(n29338), .n29335(n29335), 
         .n29332(n29332), .n29329(n29329), .n29326(n29326), .n29323(n29323), 
         .n29320(n29320), .n29317(n29317), .n29314(n29314), .n29311(n29311), 
         .n29308(n29308), .n29305(n29305), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n29302(n29302), .n29299(n29299), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n29296(n29296), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n57832(n57832), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n29107(n29107), .n29110(n29110), .n29113(n29113), .n57504(n57504), 
         .n29165(n29165), .n29184(n29184), .n29188(n29188), .n29191(n29191), 
         .n29194(n29194), .n29206(n29206), .n29209(n29209), .n57962(n57962), 
         .\data_out_frame[8][3] (\data_out_frame[8] [3]), .n57961(n57961), 
         .\data_out_frame[8][4] (\data_out_frame[8] [4]), .n57960(n57960), 
         .\data_out_frame[8][5] (\data_out_frame[8] [5]), .n57959(n57959), 
         .\data_out_frame[8][6] (\data_out_frame[8] [6]), .n57958(n57958), 
         .\data_out_frame[8][7] (\data_out_frame[8] [7]), .n57957(n57957), 
         .rx_data_ready(rx_data_ready), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n68783(n68783), .\encoder0_position_scaled[7] (encoder0_position_scaled[7]), 
         .\encoder0_position_scaled[6] (encoder0_position_scaled[6]), .\encoder0_position_scaled[5] (encoder0_position_scaled[5]), 
         .\encoder0_position_scaled[4] (encoder0_position_scaled[4]), .\encoder0_position_scaled[3] (encoder0_position_scaled[3]), 
         .\encoder0_position_scaled[15] (encoder0_position_scaled[15]), .n58003(n58003), 
         .n58002(n58002), .n58001(n58001), .n58000(n58000), .n57999(n57999), 
         .n57998(n57998), .n57997(n57997), .n57956(n57956), .n57955(n57955), 
         .n26(n26_adj_5844), .n57954(n57954), .n57953(n57953), .n57952(n57952), 
         .n57951(n57951), .n57950(n57950), .n57949(n57949), .n57948(n57948), 
         .n57947(n57947), .n57946(n57946), .n57945(n57945), .n57944(n57944), 
         .n57943(n57943), .n57942(n57942), .n57941(n57941), .n57940(n57940), 
         .n57939(n57939), .n57938(n57938), .n57937(n57937), .n57936(n57936), 
         .n57935(n57935), .n57934(n57934), .n57933(n57933), .n57932(n57932), 
         .n57931(n57931), .n57930(n57930), .n57929(n57929), .n57928(n57928), 
         .n57927(n57927), .n57926(n57926), .n57925(n57925), .n57924(n57924), 
         .n57923(n57923), .n57922(n57922), .n57921(n57921), .n57920(n57920), 
         .n57919(n57919), .n57918(n57918), .n57917(n57917), .n57916(n57916), 
         .n57915(n57915), .n57914(n57914), .n57913(n57913), .n57912(n57912), 
         .n57911(n57911), .n57898(n57898), .n57910(n57910), .n57909(n57909), 
         .n57908(n57908), .n57897(n57897), .n28838(n28838), .n28837(n28837), 
         .n57907(n57907), .n57906(n57906), .n57904(n57904), .n57905(n57905), 
         .n57833(n57833), .n28831(n28831), .n57903(n57903), .n57902(n57902), 
         .n57901(n57901), .n28827(n28827), .n57900(n57900), .n28825(n28825), 
         .n57899(n57899), .n57891(n57891), .n57890(n57890), .LED_c(LED_c), 
         .n29052(n29052), .n22362(n22362), .n58147(n58147), .n27920(n27920), 
         .DE_c(DE_c), .n57889(n57889), .n29018(n29018), .current_limit({Open_35, 
         current_limit[14:0]}), .n29017(n29017), .control_mode({control_mode}), 
         .n29016(n29016), .n58819(n58819), .\Ki[0] (Ki[0]), .n10(n10_adj_5832), 
         .n38(n38), .n27972(n27972), .n1510(n1510), .n10_adj_6(n10_adj_5841), 
         .n58707(n58707), .n58653(n58653), .n2076(n2076), .n57888(n57888), 
         .n29486(n29486), .n27600(n27600), .n363(n363), .n35(n35), .n29495(n29495), 
         .n29498(n29498), .n28969(n28969), .n28972(n28972), .n29501(n29501), 
         .n29504(n29504), .n28976(n28976), .n28979(n28979), .n29507(n29507), 
         .n29510(n29510), .n57380(n57380), .n29516(n29516), .n57378(n57378), 
         .n28982(n28982), .n57376(n57376), .n57374(n57374), .n57372(n57372), 
         .n57370(n57370), .n29593(n29593), .n29599(n29599), .n29602(n29602), 
         .n29605(n29605), .n29608(n29608), .n29951(n29951), .n29948(n29948), 
         .n29945(n29945), .n29942(n29942), .\Kp[0] (Kp[0]), .n28987(n28987), 
         .n57356(n57356), .n57354(n57354), .n57350(n57350), .n57346(n57346), 
         .n29704(n29704), .n28993(n28993), .\data_in_frame[2][3] (\data_in_frame[2] [3]), 
         .n29000(n29000), .deadband({deadband}), .IntegralLimit({IntegralLimit}), 
         .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), 
         .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), 
         .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), 
         .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[1] (Ki[1]), 
         .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
         .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), 
         .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
         .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .n29778(n29778), .n29777(n29777), 
         .n29776(n29776), .n29775(n29775), .n29774(n29774), .n29773(n29773), 
         .n29772(n29772), .n29771(n29771), .n29770(n29770), .n29769(n29769), 
         .n29768(n29768), .n29767(n29767), .n29765(n29765), .n29763(n29763), 
         .n29762(n29762), .n29761(n29761), .n29760(n29760), .n29759(n29759), 
         .n29758(n29758), .n29757(n29757), .n29756(n29756), .n29755(n29755), 
         .n29754(n29754), .n29753(n29753), .n29752(n29752), .n29751(n29751), 
         .n29750(n29750), .n29749(n29749), .n29748(n29748), .n29747(n29747), 
         .n29745(n29745), .n29744(n29744), .n29743(n29743), .n29742(n29742), 
         .n29740(n29740), .n29739(n29739), .n29738(n29738), .n29737(n29737), 
         .n29736(n29736), .n29735(n29735), .n57887(n57887), .n29009(n29009), 
         .n29013(n29013), .n29020(n29020), .n29024(n29024), .n29028(n29028), 
         .n7_adj_7(n7_adj_5862), .n29044(n29044), .n27968(n27968), .\encoder0_position_scaled[14] (encoder0_position_scaled[14]), 
         .n53279(n53279), .n28002(n28002), .n53121(n53121), .n58777(n58777), 
         .tx_active(tx_active), .n58922(n58922), .n1130(n1130), .n58644(n58644), 
         .\encoder0_position_scaled[13] (encoder0_position_scaled[13]), .n58225(n58225), 
         .n58436(n58436), .n58919(n58919), .n58245(n58245), .n25237(n25237), 
         .n25996(n25996), .n58312(n58312), .n58828(n58828), .n58446(n58446), 
         .n58680(n58680), .n27997(n27997), .n27994(n27994), .n58835(n58835), 
         .n1191(n1191), .n58845(n58845), .n58276(n58276), .n58742(n58742), 
         .n58321(n58321), .n25269(n25269), .n58925(n58925), .n58857(n58857), 
         .n58363(n58363), .n58608(n58608), .n26180(n26180), .\encoder0_position_scaled[19] (encoder0_position_scaled[19]), 
         .\encoder0_position_scaled[18] (encoder0_position_scaled[18]), .\encoder0_position_scaled[17] (encoder0_position_scaled[17]), 
         .\encoder0_position_scaled[16] (encoder0_position_scaled[16]), .\encoder0_position_scaled[12] (encoder0_position_scaled[12]), 
         .\current[15] (current[15]), .n30(n30), .n296(n296), .\encoder0_position_scaled[11] (encoder0_position_scaled[11]), 
         .ID({ID}), .\current[7] (current[7]), .\current[6] (current[6]), 
         .\current[5] (current[5]), .\current[4] (current[4]), .\current[3] (current[3]), 
         .\current[2] (current[2]), .\current[1] (current[1]), .\encoder0_position_scaled[10] (encoder0_position_scaled[10]), 
         .\current[0] (current[0]), .\current[11] (current[11]), .\current[10] (current[10]), 
         .\current[9] (current[9]), .\current[8] (current[8]), .\encoder0_position_scaled[9] (encoder0_position_scaled[9]), 
         .\encoder0_position_scaled[8] (encoder0_position_scaled[8]), .\encoder0_position_scaled[23] (encoder0_position_scaled[23]), 
         .n21(n21_adj_5814), .n19(n19_adj_5816), .n20(n20_adj_5815), .n58143(n58143), 
         .n58632(n58632), .n68699(n68699), .n58142(n58142), .n53(n53_adj_5834), 
         .n58141(n58141), .n58185(n58185), .n53988(n53988), .n68675(n68675), 
         .n68663(n68663), .n58140(n58140), .n58144(n58144), .n58145(n58145), 
         .n58139(n58139), .n60939(n60939), .n68639(n68639), .n62904(n62904), 
         .n62902(n62902), .n7_adj_8(n7_adj_5837), .n7_adj_9(n7_adj_5839), 
         .n7_adj_10(n7_adj_5838), .n1828(n1828), .n209(n209), .n270(n270), 
         .n68633(n68633), .r_Clock_Count({r_Clock_Count_adj_5940}), .n1(n1), 
         .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_5939}), .\r_Bit_Index[0] (r_Bit_Index_adj_5941[0]), 
         .n27(n27), .\tx_data[6] (tx_data[6]), .\tx_data[3] (tx_data[3]), 
         .\tx_data[2] (tx_data[2]), .\tx_data[1] (tx_data[1]), .n58968(n58968), 
         .n29040(n29040), .n69042(n69042), .n29653(n29653), .n27295(n27295), 
         .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .n4894(n4894), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
         .n29(n29), .n23(n23_adj_5840), .n61278(n61278), .n6(n6_adj_5836), 
         .tx_enable(tx_enable), .baudrate({baudrate}), .r_Clock_Count_adj_22({r_Clock_Count}), 
         .n25117(n25117), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), .\r_SM_Main[2]_adj_19 (r_SM_Main[2]), 
         .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .r_Rx_Data(r_Rx_Data), 
         .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), 
         .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), 
         .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), 
         .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), .n4891(n4891), .\r_Bit_Index[0]_adj_20 (r_Bit_Index[0]), 
         .\r_SM_Main[1]_adj_21 (r_SM_Main[1]), .n58022(n58022), .n27288(n27288), 
         .n58970(n58970), .n61676(n61676), .n61604(n61604), .n61658(n61658), 
         .n61640(n61640), .n61586(n61586), .n61622(n61622), .n61550(n61550), 
         .n29912(n29912), .n29911(n29911), .n29910(n29910), .n29909(n29909), 
         .n29908(n29908), .n29907(n29907), .n29906(n29906), .n29663(n29663), 
         .n54370(n54370), .n29667(n29667), .n27292(n27292), .n61568(n61568), 
         .n61280(n61280)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i12957_4_lut (.I0(n27262), .I1(n1405), .I2(n65449), .I3(n38907), 
            .O(n28671));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i12957_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 n9618_bdd_4_lut_51866 (.I0(n9618), .I1(n420), .I2(current[15]), 
            .I3(duty[23]), .O(n68936));
    defparam n9618_bdd_4_lut_51866.LUT_INIT = 16'he4aa;
    SB_LUT4 n68936_bdd_4_lut (.I0(n68936), .I1(duty[21]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam n68936_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13350_3_lut (.I0(current[11]), .I1(data_adj_5926[11]), .I2(n27270), 
            .I3(GND_net), .O(n29093));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_2056 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[6] [7]), .I3(\data_in_frame[6] [1]), .O(n58867));
    defparam i2_3_lut_4_lut_adj_2056.LUT_INIT = 16'h6996;
    SB_LUT4 n9618_bdd_4_lut_51861 (.I0(n9618), .I1(n421), .I2(current[15]), 
            .I3(duty[23]), .O(n68930));
    defparam n9618_bdd_4_lut_51861.LUT_INIT = 16'he4aa;
    EEPROM eeprom (.GND_net(GND_net), .enable_slow_N_4211(enable_slow_N_4211), 
           .ready_prev(ready_prev), .clk16MHz(clk16MHz), .n5753({n5754}), 
           .\state[2] (state_adj_5919[2]), .\state[0] (state_adj_5919[0]), 
           .\state[1] (state_adj_5919[1]), .n58096(n58096), .data({data_adj_5918}), 
           .ID({ID}), .n25014(n25014), .\state[0]_adj_3 (state_adj_5949[0]), 
           .baudrate({baudrate}), .n29123(n29123), .n29122(n29122), .n29121(n29121), 
           .n29120(n29120), .n29119(n29119), .n29118(n29118), .n29117(n29117), 
           .n29116(n29116), .n39313(n39313), .n29033(n29033), .rw(rw), 
           .n57558(n57558), .data_ready(data_ready), .n57286(n57286), 
           .n57342(n57342), .n38869(n38869), .\state_7__N_3916[0] (state_7__N_3916[0]), 
           .n4(n4_adj_5866), .n25133(n25133), .n60892(n60892), .VCC_net(VCC_net), 
           .scl_enable(scl_enable), .\state_7__N_4108[0] (state_7__N_4108[0]), 
           .n6388(n6388), .n29039(n29039), .\saved_addr[0] (saved_addr[0]), 
           .sda_enable(sda_enable), .scl(scl), .n4_adj_4(n4_adj_5752), 
           .n29920(n29920), .n29919(n29919), .n29918(n29918), .n29917(n29917), 
           .n29916(n29916), .n29915(n29915), .n29914(n29914), .n4_adj_5(n4_adj_5753), 
           .n29647(n29647), .n38965(n38965), .n8(n8_adj_5860), .\state_7__N_4124[3] (state_7__N_4124[3]), 
           .n10(n10_adj_5833), .n6(n6_adj_5846), .n38852(n38852), .sda_out(sda_out), 
           .n25136(n25136), .n25119(n25119)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(390[10] 402[6])
    SB_LUT4 i13351_3_lut (.I0(current[10]), .I1(data_adj_5926[10]), .I2(n27270), 
            .I3(GND_net), .O(n29094));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n68930_bdd_4_lut (.I0(n68930), .I1(duty[20]), .I2(n250), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam n68930_bdd_4_lut.LUT_INIT = 16'haad8;
    pwm PWM (.pwm_setpoint({pwm_setpoint}), .GND_net(GND_net), .n39(n39), 
        .n3014(n3014), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .\pwm_counter[19] (pwm_counter[19]), 
        .reset(reset), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 i14007_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n22362), .I3(GND_net), .O(n29750));   // verilog/coms.v(130[12] 305[6])
    defparam i14007_3_lut.LUT_INIT = 16'hcaca;
    motorControl control (.GND_net(GND_net), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .VCC_net(VCC_net), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .n363(n363), .\Kp[2] (Kp[2]), 
            .\Kp[0] (Kp[0]), .\Kp[1] (Kp[1]), .\Kp[6] (Kp[6]), .\Kp[3] (Kp[3]), 
            .IntegralLimit({IntegralLimit}), .\PID_CONTROLLER.integral_23__N_3715 ({\PID_CONTROLLER.integral_23__N_3715 }), 
            .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Kp[11] (Kp[11]), .PWMLimit({PWMLimit}), 
            .\Ki[2] (Ki[2]), .\Kp[12] (Kp[12]), .\Ki[3] (Ki[3]), .deadband({deadband}), 
            .\Ki[4] (Ki[4]), .\Ki[11] (Ki[11]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .n29183(n29183), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .n29182(n29182), .n29181(n29181), .n29180(n29180), .n29179(n29179), 
            .n29178(n29178), .n29177(n29177), .n29176(n29176), .n29175(n29175), 
            .n29174(n29174), .n29173(n29173), .n29172(n29172), .n29171(n29171), 
            .n29170(n29170), .n29169(n29169), .n29168(n29168), .n29164(n29164), 
            .n29160(n29160), .n29159(n29159), .n29158(n29158), .n29157(n29157), 
            .n29156(n29156), .n29155(n29155), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
            .\Ki[12] (Ki[12]), .\Kp[13] (Kp[13]), .n29023(n29023), .\Kp[14] (Kp[14]), 
            .\Kp[15] (Kp[15]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), 
            .\Kp[10] (Kp[10]), .n35(n35), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
            .\Ki[15] (Ki[15]), .setpoint({setpoint}), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .n14(n14_adj_5843), .\motor_state[17] (motor_state[17]), .\motor_state[16] (motor_state[16]), 
            .\encoder1_position_scaled[0] (encoder1_position_scaled[0]), .n15(n15_adj_5731), 
            .n65364(n65364), .n15_adj_1(n15_adj_5725), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .\encoder1_position_scaled[1] (encoder1_position_scaled[1]), 
            .n65475(n65475), .\motor_state[13] (motor_state[13]), .\encoder1_position_scaled[2] (encoder1_position_scaled[2]), 
            .n65474(n65474), .\motor_state[12] (motor_state[12]), .\motor_state[11] (motor_state[11]), 
            .\motor_state[10] (motor_state[10]), .n38106(n38106), .\motor_state[8] (motor_state[8]), 
            .\motor_state[7] (motor_state[7]), .\motor_state[6] (motor_state[6]), 
            .\motor_state[5] (motor_state[5]), .\motor_state[4] (motor_state[4]), 
            .\motor_state[3] (motor_state[3]), .n25(n25)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 302[4])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (GND_net, clk16MHz, n111, state, 
            neopxl_color, \bit_ctr[1] , \bit_ctr[0] , n29244, VCC_net, 
            n5, n25, timer, n29205, \neo_pixel_transmitter.t0 , n29204, 
            n29203, n27429, n29202, n29201, n29200, n29199, n29198, 
            n29197, n29187, n29043, NEOPXL_c, n23, n39366, LED_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    output n111;
    output [1:0]state;
    input [23:0]neopxl_color;
    output \bit_ctr[1] ;
    output \bit_ctr[0] ;
    input n29244;
    input VCC_net;
    input n5;
    output n25;
    output [10:0]timer;
    input n29205;
    output [10:0]\neo_pixel_transmitter.t0 ;
    input n29204;
    input n29203;
    output n27429;
    input n29202;
    input n29201;
    input n29200;
    input n29199;
    input n29198;
    input n29197;
    input n29187;
    input n29043;
    output NEOPXL_c;
    output n23;
    output n39366;
    input LED_c;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done , n52751, start, n65560, \neo_pixel_transmitter.done_N_516 , 
        n61019, start_N_507, n7;
    wire [10:0]one_wire_N_479;
    
    wire n115, n41, n59124, n59074, n112, n68834;
    wire [5:0]color_bit_N_502;
    
    wire n68837;
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [31:0]n137;
    
    wire n6858, n68618, n59, n33;
    wire [10:0]n49;
    
    wire n68954, n28943, n36565, n68606, n52000, n51999, n51998, 
        n51997, n51996, n51995, n51994, n51993, n51992, n51991, 
        n1, n27423, n28420;
    wire [1:0]state_1__N_440;
    
    wire n27228, n28419, \neo_pixel_transmitter.done_N_524 , n27247, 
        n61025, n59076, n62599, n41_adj_5678, n53189, n58984, n65557, 
        n62791, n62792, n62795, n62794, n59160;
    wire [10:0]n13;
    
    wire n4, n51178, n51177, n51176, n51175, n7_adj_5682, n51174, 
        n6_adj_5683, n51173, n51172, n51171, n51170, n51169, n59184, 
        n48, n54_adj_5684, n39315, n53158, n68609, n68957, n67443, 
        n68657, n67735, n68621, n65552, n25093, n25094, n68654;
    
    SB_LUT4 i48770_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n52751), 
            .I2(start), .I3(GND_net), .O(n65560));   // verilog/neopixel.v(16[11:16])
    defparam i48770_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n61019), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n52751), 
            .I2(start), .I3(GND_net), .O(n111));   // verilog/neopixel.v(16[11:16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut (.I0(one_wire_N_479[10]), .I1(n115), .I2(GND_net), 
            .I3(GND_net), .O(n41));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n59124), .I1(n59074), .I2(n112), .I3(state[0]), 
            .O(n52751));   // verilog/neopixel.v(16[11:16])
    defparam i1_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 n68834_bdd_4_lut (.I0(n68834), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(color_bit_N_502[1]), .O(n68837));
    defparam n68834_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2093_2_lut_3_lut_4_lut (.I0(bit_ctr[2]), .I1(\bit_ctr[1] ), 
            .I2(\bit_ctr[0] ), .I3(bit_ctr[3]), .O(n137[3]));   // verilog/neopixel.v(68[23:32])
    defparam i2093_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_DFFE bit_ctr_i1 (.Q(\bit_ctr[1] ), .C(clk16MHz), .E(VCC_net), .D(n29244));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n5));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i2081_2_lut (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n6858));   // verilog/neopixel.v(68[23:32])
    defparam i2081_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 bit_ctr_0__bdd_4_lut_51777_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(\bit_ctr[1] ), .O(n68618));
    defparam bit_ctr_0__bdd_4_lut_51777_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n112), .I1(n59), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n33));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hdccd;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(state[1]), .I1(n33), .I2(n59074), .I3(start), 
            .O(n25));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'haaae;
    SB_DFF timer_1930__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n29205));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(\bit_ctr[1] ), .O(n68954));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n29204));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n29203));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr[2]), .C(clk16MHz), .E(n27429), .D(n137[2]), 
            .R(n28943));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr[3]), .C(clk16MHz), .E(n27429), .D(n137[3]), 
            .R(n28943));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i4 (.Q(bit_ctr[4]), .C(clk16MHz), .E(n27429), .D(n137[4]), 
            .R(n28943));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n29202));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n29201));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n29200));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n29199));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n29198));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n29197));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n29187));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i15_4_lut (.I0(n65560), .I1(n36565), .I2(state[1]), .I3(state[0]), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 bit_ctr_0__bdd_4_lut_51601_4_lut_4_lut (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n68606));   // verilog/neopixel.v(18[6:15])
    defparam bit_ctr_0__bdd_4_lut_51601_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 i51558_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 115[11])
    defparam i51558_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29043));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 timer_1930_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n52000), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1930_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n51999), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_11 (.CI(n51999), .I0(GND_net), .I1(timer[9]), 
            .CO(n52000));
    SB_LUT4 timer_1930_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n51998), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_10 (.CI(n51998), .I0(GND_net), .I1(timer[8]), 
            .CO(n51999));
    SB_LUT4 timer_1930_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n51997), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_9 (.CI(n51997), .I0(GND_net), .I1(timer[7]), 
            .CO(n51998));
    SB_LUT4 timer_1930_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n51996), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_8 (.CI(n51996), .I0(GND_net), .I1(timer[6]), 
            .CO(n51997));
    SB_LUT4 timer_1930_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n51995), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_7 (.CI(n51995), .I0(GND_net), .I1(timer[5]), 
            .CO(n51996));
    SB_LUT4 timer_1930_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n51994), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_6 (.CI(n51994), .I0(GND_net), .I1(timer[4]), 
            .CO(n51995));
    SB_LUT4 timer_1930_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n51993), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_5 (.CI(n51993), .I0(GND_net), .I1(timer[3]), 
            .CO(n51994));
    SB_LUT4 timer_1930_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n51992), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_4 (.CI(n51992), .I0(GND_net), .I1(timer[2]), 
            .CO(n51993));
    SB_LUT4 timer_1930_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n51991), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_3 (.CI(n51991), .I0(GND_net), .I1(timer[1]), 
            .CO(n51992));
    SB_LUT4 timer_1930_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1930_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1930_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n51991));
    SB_DFFESR bit_ctr_i0 (.Q(\bit_ctr[0] ), .C(clk16MHz), .E(n27423), 
            .D(n1), .R(n28420));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n27228), .D(state_1__N_440[0]), 
            .S(n28419));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n27247), .D(\neo_pixel_transmitter.done_N_524 ), 
            .R(n61025));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i42108_2_lut (.I0(state[1]), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n59076));
    defparam i42108_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut (.I0(n59124), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n59));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_adj_1774 (.I0(one_wire_N_479[3]), .I1(one_wire_N_479[2]), 
            .I2(GND_net), .I3(GND_net), .O(n112));
    defparam i1_2_lut_adj_1774.LUT_INIT = 16'heeee;
    SB_LUT4 i51571_4_lut (.I0(n62599), .I1(n112), .I2(one_wire_N_479[7]), 
            .I3(n59), .O(n61019));
    defparam i51571_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i20881_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(16[11:16])
    defparam i20881_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i52_3_lut (.I0(bit_ctr[2]), .I1(bit_ctr[3]), .I2(\bit_ctr[1] ), 
            .I3(GND_net), .O(n41_adj_5678));
    defparam i52_3_lut.LUT_INIT = 16'h2424;
    SB_LUT4 i3_4_lut (.I0(n53189), .I1(n41_adj_5678), .I2(\bit_ctr[1] ), 
            .I3(\bit_ctr[0] ), .O(n23));
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i42024_2_lut (.I0(n23), .I1(n39366), .I2(GND_net), .I3(GND_net), 
            .O(n58984));
    defparam i42024_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48943_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(one_wire_N_479[10]), 
            .I3(n115), .O(n65557));   // verilog/neopixel.v(34[12] 116[6])
    defparam i48943_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i13200_2_lut (.I0(n27429), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n28943));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45775_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n62791));
    defparam i45775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45776_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n62792));
    defparam i45776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45779_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n62795));
    defparam i45779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45778_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n62794));
    defparam i45778_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF timer_1930__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1930__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i42191_2_lut_3_lut (.I0(state[1]), .I1(start), .I2(n59074), 
            .I3(GND_net), .O(n59160));
    defparam i42191_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1775 (.I0(one_wire_N_479[2]), .I1(one_wire_N_479[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1775.LUT_INIT = 16'h8888;
    SB_LUT4 sub_67_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n51178), .O(one_wire_N_479[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_11_lut (.I0(one_wire_N_479[8]), .I1(timer[9]), 
            .I2(n13[9]), .I3(n51177), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_11 (.CI(n51177), .I0(timer[9]), .I1(n13[9]), 
            .CO(n51178));
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n51176), .O(one_wire_N_479[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n51176), .I0(timer[8]), .I1(n13[8]), 
            .CO(n51177));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n51175), .O(one_wire_N_479[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n51175), .I0(timer[7]), .I1(n13[7]), 
            .CO(n51176));
    SB_LUT4 sub_67_add_2_8_lut (.I0(one_wire_N_479[4]), .I1(timer[6]), .I2(n13[6]), 
            .I3(n51174), .O(n7_adj_5682)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_8 (.CI(n51174), .I0(timer[6]), .I1(n13[6]), 
            .CO(n51175));
    SB_LUT4 sub_67_add_2_7_lut (.I0(n115), .I1(timer[5]), .I2(n13[5]), 
            .I3(n51173), .O(n6_adj_5683)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_7 (.CI(n51173), .I0(timer[5]), .I1(n13[5]), 
            .CO(n51174));
    SB_LUT4 sub_67_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n13[4]), 
            .I3(n51172), .O(one_wire_N_479[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_6 (.CI(n51172), .I0(timer[4]), .I1(n13[4]), 
            .CO(n51173));
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n51171), .O(one_wire_N_479[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_5 (.CI(n51171), .I0(timer[3]), .I1(n13[3]), 
            .CO(n51172));
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n51170), .O(one_wire_N_479[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_4 (.CI(n51170), .I0(timer[2]), .I1(n13[2]), 
            .CO(n51171));
    SB_LUT4 sub_67_add_2_3_lut (.I0(n4), .I1(timer[1]), .I2(n13[1]), .I3(n51169), 
            .O(n59124)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_67_add_2_3 (.CI(n51169), .I0(timer[1]), .I1(n13[1]), 
            .CO(n51170));
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n51169));
    SB_LUT4 i1_2_lut_adj_1776 (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_502[1]));
    defparam i1_2_lut_adj_1776.LUT_INIT = 16'h6666;
    SB_LUT4 i42215_2_lut (.I0(n59124), .I1(n59160), .I2(GND_net), .I3(GND_net), 
            .O(n59184));
    defparam i42215_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i71_4_lut (.I0(n41), .I1(n59184), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[1]), .O(n48));
    defparam i71_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n112), .I1(\neo_pixel_transmitter.done_N_524 ), 
            .I2(n59124), .I3(state[0]), .O(n54_adj_5684));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'h5d55;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(state[0]), .I1(n54_adj_5684), .I2(n48), 
            .I3(n59160), .O(n27247));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'h50dc;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_524 ));   // verilog/neopixel.v(34[12] 116[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1779 (.I0(bit_ctr[3]), .I1(n39315), .I2(GND_net), 
            .I3(GND_net), .O(n53158));
    defparam i1_2_lut_adj_1779.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut (.I0(n65557), .I1(n59076), .I2(\neo_pixel_transmitter.done ), 
            .I3(n52751), .O(n28419));   // verilog/neopixel.v(34[12] 116[6])
    defparam i14_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i50427_3_lut (.I0(n68609), .I1(n68957), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n67443));
    defparam i50427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50719_3_lut (.I0(n67443), .I1(n68657), .I2(n53158), .I3(GND_net), 
            .O(n67735));   // verilog/neopixel.v(21[26:38])
    defparam i50719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49279_4_lut (.I0(n68837), .I1(n53158), .I2(n68621), .I3(color_bit_N_502[2]), 
            .O(n65552));
    defparam i49279_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23153_4_lut (.I0(n65552), .I1(n58984), .I2(n67735), .I3(n53189), 
            .O(state_1__N_440[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i23153_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 state_1__I_0_102_Mux_0_i1_4_lut (.I0(n25093), .I1(n25094), .I2(state[0]), 
            .I3(\bit_ctr[0] ), .O(n1));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_102_Mux_0_i1_4_lut.LUT_INIT = 16'hca35;
    SB_LUT4 i1_3_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n59074), .I3(n112), .O(n25094));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hbbbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1780 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n59074), .I3(n59124), .O(n25093));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_3_lut_4_lut_adj_1780.LUT_INIT = 16'hbbbf;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n41), .I3(\neo_pixel_transmitter.done_N_524 ), 
            .O(n61025));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_1781 (.I0(\neo_pixel_transmitter.done ), .I1(one_wire_N_479[10]), 
            .I2(n115), .I3(GND_net), .O(n36565));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_3_lut_adj_1781.LUT_INIT = 16'h4040;
    SB_LUT4 i2086_2_lut_3_lut (.I0(bit_ctr[2]), .I1(\bit_ctr[1] ), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n137[2]));   // verilog/neopixel.v(68[23:32])
    defparam i2086_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 bit_ctr_0__bdd_4_lut_51876_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(\bit_ctr[1] ), .O(n68834));
    defparam bit_ctr_0__bdd_4_lut_51876_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 n68606_bdd_4_lut_4_lut (.I0(color_bit_N_502[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n68606), .O(n68609));   // verilog/neopixel.v(18[6:15])
    defparam n68606_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 i1_4_lut_4_lut (.I0(n111), .I1(state[1]), .I2(n36565), .I3(state[0]), 
            .O(n27228));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'heee2;
    SB_LUT4 i1_2_lut_3_lut_adj_1782 (.I0(n111), .I1(state[1]), .I2(n27423), 
            .I3(GND_net), .O(n27429));
    defparam i1_2_lut_3_lut_adj_1782.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n58984), .I2(LED_c), .I3(state[1]), 
            .O(n27423));   // verilog/neopixel.v(35[4] 115[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 i12677_2_lut_4_lut (.I0(state[0]), .I1(n58984), .I2(LED_c), 
            .I3(state[1]), .O(n28420));   // verilog/neopixel.v(35[4] 115[11])
    defparam i12677_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23713_2_lut_3_lut (.I0(bit_ctr[3]), .I1(n39315), .I2(bit_ctr[4]), 
            .I3(GND_net), .O(n39366));
    defparam i23713_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1783 (.I0(bit_ctr[3]), .I1(n39315), .I2(bit_ctr[4]), 
            .I3(GND_net), .O(n53189));
    defparam i1_2_lut_3_lut_adj_1783.LUT_INIT = 16'h7878;
    SB_LUT4 i1_2_lut_3_lut_adj_1784 (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), 
            .I2(bit_ctr[2]), .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1784.LUT_INIT = 16'h1e1e;
    SB_LUT4 i23666_2_lut_3_lut (.I0(\bit_ctr[1] ), .I1(\bit_ctr[0] ), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n39315));
    defparam i23666_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i45592_2_lut_4_lut (.I0(n7_adj_5682), .I1(one_wire_N_479[10]), 
            .I2(n6_adj_5683), .I3(n59076), .O(n62599));   // verilog/neopixel.v(101[14:24])
    defparam i45592_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i42106_2_lut_4_lut (.I0(n7_adj_5682), .I1(one_wire_N_479[10]), 
            .I2(n6_adj_5683), .I3(one_wire_N_479[7]), .O(n59074));   // verilog/neopixel.v(101[14:24])
    defparam i42106_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n68954_bdd_4_lut (.I0(n68954), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_502[1]), .O(n68957));
    defparam n68954_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(color_bit_N_502[1]), .I1(n62794), 
            .I2(n62795), .I3(color_bit_N_502[2]), .O(n68654));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n68654_bdd_4_lut (.I0(n68654), .I1(n62792), .I2(n62791), .I3(color_bit_N_502[2]), 
            .O(n68657));
    defparam n68654_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n68618_bdd_4_lut (.I0(n68618), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(color_bit_N_502[1]), .O(n68621));
    defparam n68618_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2100_3_lut_4_lut (.I0(bit_ctr[2]), .I1(n6858), .I2(bit_ctr[3]), 
            .I3(bit_ctr[4]), .O(n137[4]));   // verilog/neopixel.v(68[23:32])
    defparam i2100_3_lut_4_lut.LUT_INIT = 16'h7f80;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (ENCODER0_B_N_keep, n1928, ENCODER0_A_N_keep, 
            n1883, GND_net, n1885, n1887, n1889, n1891, n1893, 
            n1895, n1897, n1899, n1901, n1903, \encoder0_position[20] , 
            \encoder0_position[19] , \encoder0_position[18] , \encoder0_position[17] , 
            \encoder0_position[16] , \encoder0_position[15] , \encoder0_position[14] , 
            \encoder0_position[13] , \encoder0_position[12] , \encoder0_position[11] , 
            \encoder0_position[10] , \encoder0_position[9] , \encoder0_position[8] , 
            \encoder0_position[7] , \encoder0_position[6] , \encoder0_position[5] , 
            \encoder0_position[4] , \encoder0_position[3] , \encoder0_position[2] , 
            \encoder0_position[1] , \encoder0_position[0] , VCC_net, \a_new[1] , 
            position_31__N_3827, b_prev, n29053, n1881) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1928;
    input ENCODER0_A_N_keep;
    output n1883;
    input GND_net;
    output n1885;
    output n1887;
    output n1889;
    output n1891;
    output n1893;
    output n1895;
    output n1897;
    output n1899;
    output n1901;
    output n1903;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    output \a_new[1] ;
    output position_31__N_3827;
    output b_prev;
    input n29053;
    output n1881;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3832, n52092, n52091, n52090, n52089, n52088, 
        n52087, n52086, n52085, n52084, n52083, n52082, n52081, 
        a_prev_N_3835, debounce_cnt, n52080, n52079, n52078, n52077, 
        n52076, n52075, n52074, n52073, n52072, n52071, n52070, 
        n52069, n52068, n52067, n52066, n52065, n52064, n52063, 
        n52062, n29055, a_prev, n29054, position_31__N_3830;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1928), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1928), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1935_add_4_33_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1883), .I3(n52092), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1935_add_4_32_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1885), .I3(n52091), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_32 (.CI(n52091), .I0(direction_N_3832), 
            .I1(n1885), .CO(n52092));
    SB_LUT4 position_1935_add_4_31_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1887), .I3(n52090), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_31 (.CI(n52090), .I0(direction_N_3832), 
            .I1(n1887), .CO(n52091));
    SB_LUT4 position_1935_add_4_30_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1889), .I3(n52089), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_30 (.CI(n52089), .I0(direction_N_3832), 
            .I1(n1889), .CO(n52090));
    SB_LUT4 position_1935_add_4_29_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1891), .I3(n52088), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_29 (.CI(n52088), .I0(direction_N_3832), 
            .I1(n1891), .CO(n52089));
    SB_LUT4 position_1935_add_4_28_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1893), .I3(n52087), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_28 (.CI(n52087), .I0(direction_N_3832), 
            .I1(n1893), .CO(n52088));
    SB_LUT4 position_1935_add_4_27_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1895), .I3(n52086), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_27 (.CI(n52086), .I0(direction_N_3832), 
            .I1(n1895), .CO(n52087));
    SB_LUT4 position_1935_add_4_26_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1897), .I3(n52085), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_26 (.CI(n52085), .I0(direction_N_3832), 
            .I1(n1897), .CO(n52086));
    SB_LUT4 position_1935_add_4_25_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1899), .I3(n52084), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_25 (.CI(n52084), .I0(direction_N_3832), 
            .I1(n1899), .CO(n52085));
    SB_LUT4 position_1935_add_4_24_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1901), .I3(n52083), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_24 (.CI(n52083), .I0(direction_N_3832), 
            .I1(n1901), .CO(n52084));
    SB_LUT4 position_1935_add_4_23_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1903), .I3(n52082), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_23 (.CI(n52082), .I0(direction_N_3832), 
            .I1(n1903), .CO(n52083));
    SB_LUT4 position_1935_add_4_22_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[20] ), .I3(n52081), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1928), .D(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_1935_add_4_22 (.CI(n52081), .I0(direction_N_3832), 
            .I1(\encoder0_position[20] ), .CO(n52082));
    SB_LUT4 position_1935_add_4_21_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[19] ), .I3(n52080), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_21 (.CI(n52080), .I0(direction_N_3832), 
            .I1(\encoder0_position[19] ), .CO(n52081));
    SB_LUT4 position_1935_add_4_20_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[18] ), .I3(n52079), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_20 (.CI(n52079), .I0(direction_N_3832), 
            .I1(\encoder0_position[18] ), .CO(n52080));
    SB_LUT4 position_1935_add_4_19_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[17] ), .I3(n52078), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_19 (.CI(n52078), .I0(direction_N_3832), 
            .I1(\encoder0_position[17] ), .CO(n52079));
    SB_LUT4 position_1935_add_4_18_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[16] ), .I3(n52077), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_18 (.CI(n52077), .I0(direction_N_3832), 
            .I1(\encoder0_position[16] ), .CO(n52078));
    SB_LUT4 position_1935_add_4_17_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[15] ), .I3(n52076), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_17 (.CI(n52076), .I0(direction_N_3832), 
            .I1(\encoder0_position[15] ), .CO(n52077));
    SB_LUT4 position_1935_add_4_16_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[14] ), .I3(n52075), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_16 (.CI(n52075), .I0(direction_N_3832), 
            .I1(\encoder0_position[14] ), .CO(n52076));
    SB_LUT4 position_1935_add_4_15_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[13] ), .I3(n52074), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_15 (.CI(n52074), .I0(direction_N_3832), 
            .I1(\encoder0_position[13] ), .CO(n52075));
    SB_LUT4 position_1935_add_4_14_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[12] ), .I3(n52073), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_14 (.CI(n52073), .I0(direction_N_3832), 
            .I1(\encoder0_position[12] ), .CO(n52074));
    SB_LUT4 position_1935_add_4_13_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[11] ), .I3(n52072), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_13 (.CI(n52072), .I0(direction_N_3832), 
            .I1(\encoder0_position[11] ), .CO(n52073));
    SB_LUT4 position_1935_add_4_12_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[10] ), .I3(n52071), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_12 (.CI(n52071), .I0(direction_N_3832), 
            .I1(\encoder0_position[10] ), .CO(n52072));
    SB_LUT4 position_1935_add_4_11_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[9] ), .I3(n52070), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_11 (.CI(n52070), .I0(direction_N_3832), 
            .I1(\encoder0_position[9] ), .CO(n52071));
    SB_LUT4 position_1935_add_4_10_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[8] ), .I3(n52069), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_10 (.CI(n52069), .I0(direction_N_3832), 
            .I1(\encoder0_position[8] ), .CO(n52070));
    SB_LUT4 position_1935_add_4_9_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[7] ), .I3(n52068), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_9 (.CI(n52068), .I0(direction_N_3832), 
            .I1(\encoder0_position[7] ), .CO(n52069));
    SB_LUT4 position_1935_add_4_8_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[6] ), .I3(n52067), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_8 (.CI(n52067), .I0(direction_N_3832), 
            .I1(\encoder0_position[6] ), .CO(n52068));
    SB_LUT4 position_1935_add_4_7_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[5] ), .I3(n52066), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_7 (.CI(n52066), .I0(direction_N_3832), 
            .I1(\encoder0_position[5] ), .CO(n52067));
    SB_LUT4 position_1935_add_4_6_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[4] ), .I3(n52065), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_6 (.CI(n52065), .I0(direction_N_3832), 
            .I1(\encoder0_position[4] ), .CO(n52066));
    SB_LUT4 position_1935_add_4_5_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[3] ), .I3(n52064), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_5 (.CI(n52064), .I0(direction_N_3832), 
            .I1(\encoder0_position[3] ), .CO(n52065));
    SB_LUT4 position_1935_add_4_4_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[2] ), .I3(n52063), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_4 (.CI(n52063), .I0(direction_N_3832), 
            .I1(\encoder0_position[2] ), .CO(n52064));
    SB_LUT4 position_1935_add_4_3_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[1] ), .I3(n52062), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_3 (.CI(n52062), .I0(direction_N_3832), 
            .I1(\encoder0_position[1] ), .CO(n52063));
    SB_LUT4 position_1935_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1935_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1935_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n52062));
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1928), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1928), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1935__i0 (.Q(\encoder0_position[0] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1928), .D(n29055));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1928), .D(n29054));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n1881), .C(n1928), .D(n29053));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1935__i1 (.Q(\encoder0_position[1] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i2 (.Q(\encoder0_position[2] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i3 (.Q(\encoder0_position[3] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i4 (.Q(\encoder0_position[4] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i5 (.Q(\encoder0_position[5] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i6 (.Q(\encoder0_position[6] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i7 (.Q(\encoder0_position[7] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i8 (.Q(\encoder0_position[8] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i9 (.Q(\encoder0_position[9] ), .C(n1928), .E(position_31__N_3827), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i10 (.Q(\encoder0_position[10] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i11 (.Q(\encoder0_position[11] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i12 (.Q(\encoder0_position[12] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i13 (.Q(\encoder0_position[13] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i14 (.Q(\encoder0_position[14] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i15 (.Q(\encoder0_position[15] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i16 (.Q(\encoder0_position[16] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i17 (.Q(\encoder0_position[17] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i18 (.Q(\encoder0_position[18] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i19 (.Q(\encoder0_position[19] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i20 (.Q(\encoder0_position[20] ), .C(n1928), 
            .E(position_31__N_3827), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i21 (.Q(n1903), .C(n1928), .E(position_31__N_3827), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i22 (.Q(n1901), .C(n1928), .E(position_31__N_3827), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i23 (.Q(n1899), .C(n1928), .E(position_31__N_3827), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i24 (.Q(n1897), .C(n1928), .E(position_31__N_3827), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i25 (.Q(n1895), .C(n1928), .E(position_31__N_3827), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i26 (.Q(n1893), .C(n1928), .E(position_31__N_3827), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i27 (.Q(n1891), .C(n1928), .E(position_31__N_3827), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i28 (.Q(n1889), .C(n1928), .E(position_31__N_3827), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i29 (.Q(n1887), .C(n1928), .E(position_31__N_3827), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i30 (.Q(n1885), .C(n1928), .E(position_31__N_3827), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1935__i31 (.Q(n1883), .C(n1928), .E(position_31__N_3827), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 i51432_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i51432_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 i13312_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29055));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13312_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13311_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(b_new[1]), 
            .I3(b_prev), .O(n29054));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13311_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3832));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3830));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3830), 
            .I3(\a_new[1] ), .O(position_31__N_3827));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (encoder1_position, GND_net, VCC_net, ENCODER1_B_N_keep, 
            n1928, ENCODER1_A_N_keep, \a_new[1] , position_31__N_3827, 
            n29051, n1933, b_prev) /* synthesis lattice_noprune=1 */ ;
    output [31:0]encoder1_position;
    input GND_net;
    input VCC_net;
    input ENCODER1_B_N_keep;
    input n1928;
    input ENCODER1_A_N_keep;
    output \a_new[1] ;
    output position_31__N_3827;
    input n29051;
    output n1933;
    output b_prev;
    
    wire [31:0]n133;
    
    wire direction_N_3832, n52154, n52153, n52152, n52151, n52150, 
        n52149, n52148, n52147, n52146, n52145, n52144, n52143, 
        n52142, n52141, n52140, n52139, n52138, n52137, n52136, 
        n52135, n52134, n52133, n52132, n52131, n52130, n52129, 
        n52128, n52127, n52126, n52125, n52124;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3835, debounce_cnt, n29050, n29049, a_prev, position_31__N_3830;
    
    SB_LUT4 position_1937_add_4_33_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[31]), .I3(n52154), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1937_add_4_32_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[30]), .I3(n52153), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_32 (.CI(n52153), .I0(direction_N_3832), 
            .I1(encoder1_position[30]), .CO(n52154));
    SB_LUT4 position_1937_add_4_31_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[29]), .I3(n52152), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_31 (.CI(n52152), .I0(direction_N_3832), 
            .I1(encoder1_position[29]), .CO(n52153));
    SB_LUT4 position_1937_add_4_30_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[28]), .I3(n52151), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_30 (.CI(n52151), .I0(direction_N_3832), 
            .I1(encoder1_position[28]), .CO(n52152));
    SB_LUT4 position_1937_add_4_29_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[27]), .I3(n52150), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_29 (.CI(n52150), .I0(direction_N_3832), 
            .I1(encoder1_position[27]), .CO(n52151));
    SB_LUT4 position_1937_add_4_28_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[26]), .I3(n52149), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_28 (.CI(n52149), .I0(direction_N_3832), 
            .I1(encoder1_position[26]), .CO(n52150));
    SB_LUT4 position_1937_add_4_27_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[25]), .I3(n52148), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_27 (.CI(n52148), .I0(direction_N_3832), 
            .I1(encoder1_position[25]), .CO(n52149));
    SB_LUT4 position_1937_add_4_26_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[24]), .I3(n52147), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_26 (.CI(n52147), .I0(direction_N_3832), 
            .I1(encoder1_position[24]), .CO(n52148));
    SB_LUT4 position_1937_add_4_25_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[23]), .I3(n52146), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_25 (.CI(n52146), .I0(direction_N_3832), 
            .I1(encoder1_position[23]), .CO(n52147));
    SB_LUT4 position_1937_add_4_24_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[22]), .I3(n52145), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_24 (.CI(n52145), .I0(direction_N_3832), 
            .I1(encoder1_position[22]), .CO(n52146));
    SB_LUT4 position_1937_add_4_23_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[21]), .I3(n52144), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_23 (.CI(n52144), .I0(direction_N_3832), 
            .I1(encoder1_position[21]), .CO(n52145));
    SB_LUT4 position_1937_add_4_22_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[20]), .I3(n52143), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_22 (.CI(n52143), .I0(direction_N_3832), 
            .I1(encoder1_position[20]), .CO(n52144));
    SB_LUT4 position_1937_add_4_21_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[19]), .I3(n52142), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_21 (.CI(n52142), .I0(direction_N_3832), 
            .I1(encoder1_position[19]), .CO(n52143));
    SB_LUT4 position_1937_add_4_20_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[18]), .I3(n52141), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_20 (.CI(n52141), .I0(direction_N_3832), 
            .I1(encoder1_position[18]), .CO(n52142));
    SB_LUT4 position_1937_add_4_19_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[17]), .I3(n52140), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_19 (.CI(n52140), .I0(direction_N_3832), 
            .I1(encoder1_position[17]), .CO(n52141));
    SB_LUT4 position_1937_add_4_18_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[16]), .I3(n52139), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_18 (.CI(n52139), .I0(direction_N_3832), 
            .I1(encoder1_position[16]), .CO(n52140));
    SB_LUT4 position_1937_add_4_17_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[15]), .I3(n52138), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_17 (.CI(n52138), .I0(direction_N_3832), 
            .I1(encoder1_position[15]), .CO(n52139));
    SB_LUT4 position_1937_add_4_16_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[14]), .I3(n52137), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_16 (.CI(n52137), .I0(direction_N_3832), 
            .I1(encoder1_position[14]), .CO(n52138));
    SB_LUT4 position_1937_add_4_15_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[13]), .I3(n52136), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_15 (.CI(n52136), .I0(direction_N_3832), 
            .I1(encoder1_position[13]), .CO(n52137));
    SB_LUT4 position_1937_add_4_14_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[12]), .I3(n52135), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_14 (.CI(n52135), .I0(direction_N_3832), 
            .I1(encoder1_position[12]), .CO(n52136));
    SB_LUT4 position_1937_add_4_13_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[11]), .I3(n52134), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_13 (.CI(n52134), .I0(direction_N_3832), 
            .I1(encoder1_position[11]), .CO(n52135));
    SB_LUT4 position_1937_add_4_12_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[10]), .I3(n52133), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_12 (.CI(n52133), .I0(direction_N_3832), 
            .I1(encoder1_position[10]), .CO(n52134));
    SB_LUT4 position_1937_add_4_11_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[9]), .I3(n52132), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_11 (.CI(n52132), .I0(direction_N_3832), 
            .I1(encoder1_position[9]), .CO(n52133));
    SB_LUT4 position_1937_add_4_10_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[8]), .I3(n52131), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_10 (.CI(n52131), .I0(direction_N_3832), 
            .I1(encoder1_position[8]), .CO(n52132));
    SB_LUT4 position_1937_add_4_9_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[7]), .I3(n52130), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_9 (.CI(n52130), .I0(direction_N_3832), 
            .I1(encoder1_position[7]), .CO(n52131));
    SB_LUT4 position_1937_add_4_8_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[6]), .I3(n52129), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_8 (.CI(n52129), .I0(direction_N_3832), 
            .I1(encoder1_position[6]), .CO(n52130));
    SB_LUT4 position_1937_add_4_7_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[5]), .I3(n52128), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_7 (.CI(n52128), .I0(direction_N_3832), 
            .I1(encoder1_position[5]), .CO(n52129));
    SB_LUT4 position_1937_add_4_6_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[4]), .I3(n52127), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_6 (.CI(n52127), .I0(direction_N_3832), 
            .I1(encoder1_position[4]), .CO(n52128));
    SB_LUT4 position_1937_add_4_5_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[3]), .I3(n52126), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_5 (.CI(n52126), .I0(direction_N_3832), 
            .I1(encoder1_position[3]), .CO(n52127));
    SB_LUT4 position_1937_add_4_4_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[2]), .I3(n52125), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_4 (.CI(n52125), .I0(direction_N_3832), 
            .I1(encoder1_position[2]), .CO(n52126));
    SB_LUT4 position_1937_add_4_3_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(encoder1_position[1]), .I3(n52124), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_3 (.CI(n52124), .I0(direction_N_3832), 
            .I1(encoder1_position[1]), .CO(n52125));
    SB_LUT4 position_1937_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1937_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1937_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n52124));
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1928), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1928), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1928), .D(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1928), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1928), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1937__i0 (.Q(encoder1_position[0]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF direction_40 (.Q(n1933), .C(n1928), .D(n29051));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1928), .D(n29050));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1928), .D(n29049));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1937__i1 (.Q(encoder1_position[1]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i2 (.Q(encoder1_position[2]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i3 (.Q(encoder1_position[3]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i4 (.Q(encoder1_position[4]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i5 (.Q(encoder1_position[5]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i6 (.Q(encoder1_position[6]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i7 (.Q(encoder1_position[7]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i8 (.Q(encoder1_position[8]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i9 (.Q(encoder1_position[9]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i10 (.Q(encoder1_position[10]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i11 (.Q(encoder1_position[11]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i12 (.Q(encoder1_position[12]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i13 (.Q(encoder1_position[13]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i14 (.Q(encoder1_position[14]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i15 (.Q(encoder1_position[15]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i16 (.Q(encoder1_position[16]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i17 (.Q(encoder1_position[17]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i18 (.Q(encoder1_position[18]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i19 (.Q(encoder1_position[19]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i20 (.Q(encoder1_position[20]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i21 (.Q(encoder1_position[21]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i22 (.Q(encoder1_position[22]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i23 (.Q(encoder1_position[23]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i24 (.Q(encoder1_position[24]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i25 (.Q(encoder1_position[25]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i26 (.Q(encoder1_position[26]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i27 (.Q(encoder1_position[27]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i28 (.Q(encoder1_position[28]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i29 (.Q(encoder1_position[29]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i30 (.Q(encoder1_position[30]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1937__i31 (.Q(encoder1_position[31]), .C(n1928), .E(position_31__N_3827), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 i51435_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i51435_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 i13307_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(b_new[1]), 
            .I3(b_prev), .O(n29050));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13307_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13306_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29049));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13306_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3832));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3830));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3830), 
            .I3(\a_new[1] ), .O(position_31__N_3827));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (GND_net, VCC_net, clk16MHz, n27270, \current[15] , 
            state_7__N_4317, n6, n5, n5_adj_23, n6_adj_24, n29103, 
            \current[1] , n29102, \current[2] , n29101, \current[3] , 
            n29100, \current[4] , n29099, \current[5] , n29098, \current[6] , 
            n29097, \current[7] , n29096, \current[8] , n29095, \current[9] , 
            n29094, \current[10] , n29093, \current[11] , n38922, 
            CS_c, n29032, \current[0] , n11, CS_CLK_c, n29904, \data[15] , 
            n29903, \data[12] , n29902, \data[11] , n29901, \data[10] , 
            n29900, \data[9] , n29899, \data[8] , n29898, \data[7] , 
            n29897, \data[6] , n29896, \data[5] , n29895, \data[4] , 
            n29894, \data[3] , n29893, \data[2] , n29892, \data[1] , 
            n29683, \data[0] , \duty[0] , \duty[1] , n4, n25112, 
            n25151, n25141, n25145, n25148, n6_adj_25, n5_adj_26) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input clk16MHz;
    output n27270;
    output \current[15] ;
    output state_7__N_4317;
    output n6;
    output n5;
    output n5_adj_23;
    output n6_adj_24;
    input n29103;
    output \current[1] ;
    input n29102;
    output \current[2] ;
    input n29101;
    output \current[3] ;
    input n29100;
    output \current[4] ;
    input n29099;
    output \current[5] ;
    input n29098;
    output \current[6] ;
    input n29097;
    output \current[7] ;
    input n29096;
    output \current[8] ;
    input n29095;
    output \current[9] ;
    input n29094;
    output \current[10] ;
    input n29093;
    output \current[11] ;
    output n38922;
    output CS_c;
    input n29032;
    output \current[0] ;
    output n11;
    output CS_CLK_c;
    input n29904;
    output \data[15] ;
    input n29903;
    output \data[12] ;
    input n29902;
    output \data[11] ;
    input n29901;
    output \data[10] ;
    input n29900;
    output \data[9] ;
    input n29899;
    output \data[8] ;
    input n29898;
    output \data[7] ;
    input n29897;
    output \data[6] ;
    input n29896;
    output \data[5] ;
    input n29895;
    output \data[4] ;
    input n29894;
    output \data[3] ;
    input n29893;
    output \data[2] ;
    input n29892;
    output \data[1] ;
    input n29683;
    output \data[0] ;
    input \duty[0] ;
    input \duty[1] ;
    output n4;
    output n25112;
    output n25151;
    output n25141;
    output n25145;
    output n25148;
    output n6_adj_25;
    output n5_adj_26;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n52167, n52166;
    wire [11:0]n1;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n52165, n52164, n52163, n52162, n52161, n52160, n52159, 
        n52158, n52157, n52156, n52155, clk_slow_N_4230, clk_slow_N_4231;
    wire [1:0]n2000;
    wire [7:0]n37;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n52030, n52029, n52028, n52027, n52026, n52025, n52024, 
        n65494, n6673;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n27404, n28948, n22322, delay_counter_15__N_4312, n9, clk_out, 
        n29037, n39297, n27275, n28432, n15;
    wire [7:0]n47;
    
    wire n9684, n6_adj_5676, n8, n12, n10;
    
    SB_LUT4 counter_1941_1942_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n52167), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1941_1942_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1941_1942_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n52166), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1941_1942_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1941_1942_add_4_3 (.CI(n52166), .I0(GND_net), .I1(counter[1]), 
            .CO(n52167));
    SB_LUT4 counter_1941_1942_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1941_1942_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1941_1942_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52166));
    SB_LUT4 delay_counter_1939_1940_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n52165), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1939_1940_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n52164), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_12 (.CI(n52164), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n52165));
    SB_LUT4 delay_counter_1939_1940_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n52163), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_11 (.CI(n52163), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n52164));
    SB_LUT4 delay_counter_1939_1940_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n52162), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_10 (.CI(n52162), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n52163));
    SB_LUT4 delay_counter_1939_1940_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n52161), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_9 (.CI(n52161), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n52162));
    SB_LUT4 delay_counter_1939_1940_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n52160), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_8 (.CI(n52160), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n52161));
    SB_LUT4 delay_counter_1939_1940_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n52159), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_7 (.CI(n52159), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n52160));
    SB_LUT4 delay_counter_1939_1940_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n52158), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_6 (.CI(n52158), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n52159));
    SB_LUT4 delay_counter_1939_1940_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n52157), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_5 (.CI(n52157), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n52158));
    SB_LUT4 delay_counter_1939_1940_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n52156), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_4 (.CI(n52156), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n52157));
    SB_LUT4 delay_counter_1939_1940_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n52155), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_3 (.CI(n52155), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n52156));
    SB_LUT4 delay_counter_1939_1940_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1939_1940_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1939_1940_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n52155));
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4230));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 i2057_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4231));
    defparam i2057_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4231), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4230));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27270), 
            .D(n2000[0]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_1932_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n52030), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_1932_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n52029), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1932_add_4_8 (.CI(n52029), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n52030));
    SB_LUT4 bit_counter_1932_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n52028), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1932_add_4_7 (.CI(n52028), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n52029));
    SB_LUT4 bit_counter_1932_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n52027), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1932_add_4_6 (.CI(n52027), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n52028));
    SB_LUT4 bit_counter_1932_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n52026), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1932_add_4_5 (.CI(n52026), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n52027));
    SB_LUT4 bit_counter_1932_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n52025), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1932_add_4_4 (.CI(n52025), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n52026));
    SB_LUT4 bit_counter_1932_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n52024), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1932_add_4_3 (.CI(n52024), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n52025));
    SB_LUT4 bit_counter_1932_add_4_2_lut (.I0(n6673), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n65494)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1932_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1932_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n52024));
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4317));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i11840_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27404));
    defparam i11840_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_341_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_341_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_341_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_341_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_332_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_23));   // verilog/tli4970.v(54[9:26])
    defparam equal_332_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_336_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_24));   // verilog/tli4970.v(54[9:26])
    defparam equal_336_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESR bit_counter_1932__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27404), 
            .D(n37[7]), .R(n28948));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1932__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27404), 
            .D(n37[6]), .R(n28948));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1932__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27404), 
            .D(n37[5]), .R(n28948));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1932__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27404), 
            .D(n37[4]), .R(n28948));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n29103));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n29102));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n29101));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n29100));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n29099));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n29098));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n29097));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n29096));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n29095));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n29094));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n29093));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i23276_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n38922));
    defparam i23276_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNE bit_counter_1932__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27404), 
            .D(n22322));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1939_1940__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n1[0]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1941_1942__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29037));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29032));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_272_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_272_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n27275), .D(n39297), 
            .S(n28432));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(delay_counter_15__N_4312), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n27275));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i12689_2_lut_4_lut (.I0(delay_counter_15__N_4312), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n28432));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12689_2_lut_4_lut.LUT_INIT = 16'h2202;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29904));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29903));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29902));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29901));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29900));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29899));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29898));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29897));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29896));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29895));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29894));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29893));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29892));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n29683));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1932__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27404), 
            .D(n47[1]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1932__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27404), 
            .D(n47[2]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1932__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27404), 
            .D(n47[3]));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n27275), .D(n9684), 
            .R(n28432));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNSR delay_counter_1939_1940__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n1[1]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n1[2]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n1[3]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n1[4]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n1[5]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n1[6]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n1[7]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n1[8]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n1[9]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n1[10]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1939_1940__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n1[11]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1941_1942__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1941_1942__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i1896_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n6673));   // verilog/tli4970.v(35[10] 68[6])
    defparam i1896_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_2025_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n9684));
    defparam mux_2025_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i51391_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n27270));
    defparam i51391_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2113_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2000[0]));
    defparam i2113_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18130_3_lut_4_lut (.I0(\duty[0] ), .I1(\current[0] ), .I2(\duty[1] ), 
            .I3(\current[1] ), .O(n4));   // verilog/tli4970.v(35[10] 68[6])
    defparam i18130_3_lut_4_lut.LUT_INIT = 16'h20f2;
    SB_LUT4 i51440_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n39297));
    defparam i51440_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(state[0]), 
            .I3(state[1]), .O(n25112));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_4_lut_adj_1767 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25151));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1767.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1768 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25141));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1768.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1769 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25145));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1769.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1770 (.I0(state[0]), .I1(state[1]), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25148));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1770.LUT_INIT = 16'hffbf;
    SB_LUT4 i13205_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n28948));   // verilog/tli4970.v(55[24:39])
    defparam i13205_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 bit_counter_1932_mux_6_i4_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state_7__N_4317), .I3(n37[3]), .O(n47[3]));
    defparam bit_counter_1932_mux_6_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_1932_mux_6_i3_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state_7__N_4317), .I3(n37[2]), .O(n47[2]));
    defparam bit_counter_1932_mux_6_i3_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 bit_counter_1932_mux_6_i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state_7__N_4317), .I3(n37[1]), .O(n47[1]));
    defparam bit_counter_1932_mux_6_i2_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 equal_343_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_25));   // verilog/tli4970.v(54[9:26])
    defparam equal_343_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_334_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_26));   // verilog/tli4970.v(54[9:26])
    defparam equal_334_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51574_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9));   // verilog/tli4970.v(35[10] 68[6])
    defparam i51574_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i13294_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n29037));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13294_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5676));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_adj_5676), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2058_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2058_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut_adj_1771 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(delay_counter[8]), .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut_adj_1771.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4312));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i6820_3_lut (.I0(state[0]), .I1(n65494), .I2(state[1]), .I3(GND_net), 
            .O(n22322));   // verilog/tli4970.v(55[24:39])
    defparam i6820_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_in_frame[5] , n3014, \data_out_frame[18] , clk16MHz, 
            n57886, n58004, n29483, VCC_net, \data_in_frame[15] , 
            n57892, n57893, n57885, n29480, n57884, \data_in_frame[4] , 
            \data_in_frame[2] , \data_in_frame[6] , n57894, n57883, 
            \data_out_frame[19] , n57882, n57881, n57880, n57879, 
            \data_out_frame[23] , GND_net, \data_in_frame[3] , n57878, 
            \data_out_frame[1][6] , n57996, \data_out_frame[1][7] , n57995, 
            n57877, \data_in_frame[8] , \data_out_frame[17] , \FRAME_MATCHER.i_31__N_2509 , 
            pwm_setpoint, n57876, n57875, \data_out_frame[20] , n57874, 
            n57873, n25488, n57872, n57871, \data_in_frame[14] , \data_in_frame[1] , 
            n29477, Kp_23__N_869, \data_out_frame[3][1] , n57994, n57870, 
            n57869, n58867, n58698, n53862, \data_out_frame[16] , 
            n57868, n57867, \data_out_frame[3][3] , n57993, \data_in_frame[2][5] , 
            n29474, \data_in_frame[9] , \data_in_frame[11] , \data_out_frame[3][4] , 
            n57992, \data_out_frame[3][6] , n57991, \data_out_frame[3][7] , 
            n57990, \data_in_frame[3][4] , n29471, \data_out_frame[4] , 
            n28927, n57989, n57895, \data_in_frame[5][6] , n29468, 
            n57988, n57987, \data_out_frame[21] , n57866, n57865, 
            n57864, n57863, n57862, n57861, n57860, n57859, \data_out_frame[22] , 
            n57858, n57857, n57856, n57855, n28782, n57854, n28780, 
            n57853, n57852, n57986, n29465, n57985, n62, n57984, 
            \data_out_frame[5] , n57983, n29462, n57982, n57981, n57980, 
            n29459, n57979, n57978, n57851, n29456, n57977, n29453, 
            n57976, n29450, \data_out_frame[6] , \encoder0_position_scaled[22] , 
            n57975, n29447, n57974, n29444, n28909, n57850, n57849, 
            n57848, n57847, n28772, n57896, \data_out_frame[24] , 
            n57846, n57845, n28768, n28767, n57844, n57843, n28764, 
            n57842, \data_out_frame[25] , n57841, n57840, n57839, 
            n57838, n57837, n57836, n57835, n57973, n29441, n57834, 
            neopxl_color, n22373, n58391, \data_in_frame[3][3] , \data_in_frame[5][3] , 
            n11, n12, \data_in_frame[20] , n29438, \data_in_frame[13] , 
            \data_in_frame[21] , \data_in_frame[23][2] , \data_in_frame[10] , 
            \data_out_frame[15] , \data_in_frame[23][6] , \data_in_frame[16] , 
            \data_in_frame[20][1] , n57972, \data_in_frame[3][0] , \data_in_frame[5][2] , 
            n57971, \data_in_frame[23][1] , \data_in_frame[23][7] , \data_in_frame[23][0] , 
            \data_in_frame[20][5] , reset, \data_in_frame[5][0] , n29435, 
            setpoint, \data_in_frame[20][6] , byte_transmit_counter, \data_in_frame[12] , 
            \data_in_frame[3][2] , n57970, \data_in_frame[16][5] , \data_in_frame[16][4] , 
            \byte_transmit_counter[0] , \data_out_frame[0][2] , n29432, 
            \data_out_frame[7] , \data_in_frame[17] , n29429, n57969, 
            \data_out_frame[14] , n29426, n57968, n29423, n57967, 
            rx_data, n7, \data_out_frame[13] , n29420, n29417, n29414, 
            n57966, n29411, n29408, n29405, n68861, n68855, \FRAME_MATCHER.state[3] , 
            n29402, n57965, \data_out_frame[12] , displacement, \encoder0_position_scaled[21] , 
            n29399, \data_in_frame[17][0] , PWMLimit, n29395, n57964, 
            n29392, \data_out_frame[11] , encoder1_position_scaled, n29389, 
            n29386, n27924, \data_in_frame[16][7] , n28009, n29383, 
            n29380, n68849, n29377, \data_out_frame[10] , n29374, 
            \encoder0_position_scaled[20] , n29371, n29368, n29365, 
            n29362, n29359, \data_out_frame[9] , n57963, n29356, n29353, 
            n29350, n29347, n29344, n29341, n29338, n29335, n29332, 
            n29329, n29326, n29323, n29320, n29317, n29314, n29311, 
            n29308, n29305, \data_out_frame[1][5] , n29302, n29299, 
            \data_out_frame[1][3] , n29296, \data_out_frame[1][1] , n57832, 
            \data_out_frame[1][0] , \data_out_frame[0][4] , \data_out_frame[0][3] , 
            n29107, n29110, n29113, n57504, n29165, n29184, n29188, 
            n29191, n29194, n29206, n29209, n57962, \data_out_frame[8][3] , 
            n57961, \data_out_frame[8][4] , n57960, \data_out_frame[8][5] , 
            n57959, \data_out_frame[8][6] , n57958, \data_out_frame[8][7] , 
            n57957, rx_data_ready, \FRAME_MATCHER.rx_data_ready_prev , 
            n68783, \encoder0_position_scaled[7] , \encoder0_position_scaled[6] , 
            \encoder0_position_scaled[5] , \encoder0_position_scaled[4] , 
            \encoder0_position_scaled[3] , \encoder0_position_scaled[15] , 
            n58003, n58002, n58001, n58000, n57999, n57998, n57997, 
            n57956, n57955, n26, n57954, n57953, n57952, n57951, 
            n57950, n57949, n57948, n57947, n57946, n57945, n57944, 
            n57943, n57942, n57941, n57940, n57939, n57938, n57937, 
            n57936, n57935, n57934, n57933, n57932, n57931, n57930, 
            n57929, n57928, n57927, n57926, n57925, n57924, n57923, 
            n57922, n57921, n57920, n57919, n57918, n57917, n57916, 
            n57915, n57914, n57913, n57912, n57911, n57898, n57910, 
            n57909, n57908, n57897, n28838, n28837, n57907, n57906, 
            n57904, n57905, n57833, n28831, n57903, n57902, n57901, 
            n28827, n57900, n28825, n57899, n57891, n57890, LED_c, 
            n29052, n22362, n58147, n27920, DE_c, n57889, n29018, 
            current_limit, n29017, control_mode, n29016, n58819, \Ki[0] , 
            n10, n38, n27972, n1510, n10_adj_6, n58707, n58653, 
            n2076, n57888, n29486, n27600, n363, n35, n29495, 
            n29498, n28969, n28972, n29501, n29504, n28976, n28979, 
            n29507, n29510, n57380, n29516, n57378, n28982, n57376, 
            n57374, n57372, n57370, n29593, n29599, n29602, n29605, 
            n29608, n29951, n29948, n29945, n29942, \Kp[0] , n28987, 
            n57356, n57354, n57350, n57346, n29704, n28993, \data_in_frame[2][3] , 
            n29000, deadband, IntegralLimit, \Kp[1] , \Kp[2] , \Kp[3] , 
            \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] , 
            \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , \Ki[6] , 
            \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , \Ki[12] , 
            \Ki[13] , \Ki[14] , \Ki[15] , n29778, n29777, n29776, 
            n29775, n29774, n29773, n29772, n29771, n29770, n29769, 
            n29768, n29767, n29765, n29763, n29762, n29761, n29760, 
            n29759, n29758, n29757, n29756, n29755, n29754, n29753, 
            n29752, n29751, n29750, n29749, n29748, n29747, n29745, 
            n29744, n29743, n29742, n29740, n29739, n29738, n29737, 
            n29736, n29735, n57887, n29009, n29013, n29020, n29024, 
            n29028, n7_adj_7, n29044, n27968, \encoder0_position_scaled[14] , 
            n53279, n28002, n53121, n58777, tx_active, n58922, n1130, 
            n58644, \encoder0_position_scaled[13] , n58225, n58436, 
            n58919, n58245, n25237, n25996, n58312, n58828, n58446, 
            n58680, n27997, n27994, n58835, n1191, n58845, n58276, 
            n58742, n58321, n25269, n58925, n58857, n58363, n58608, 
            n26180, \encoder0_position_scaled[19] , \encoder0_position_scaled[18] , 
            \encoder0_position_scaled[17] , \encoder0_position_scaled[16] , 
            \encoder0_position_scaled[12] , \current[15] , n30, n296, 
            \encoder0_position_scaled[11] , ID, \current[7] , \current[6] , 
            \current[5] , \current[4] , \current[3] , \current[2] , 
            \current[1] , \encoder0_position_scaled[10] , \current[0] , 
            \current[11] , \current[10] , \current[9] , \current[8] , 
            \encoder0_position_scaled[9] , \encoder0_position_scaled[8] , 
            \encoder0_position_scaled[23] , n21, n19, n20, n58143, 
            n58632, n68699, n58142, n53, n58141, n58185, n53988, 
            n68675, n68663, n58140, n58144, n58145, n58139, n60939, 
            n68639, n62904, n62902, n7_adj_8, n7_adj_9, n7_adj_10, 
            n1828, n209, n270, n68633, r_Clock_Count, n1, tx_o, 
            r_SM_Main, \r_Bit_Index[0] , n27, \tx_data[6] , \tx_data[3] , 
            \tx_data[2] , \tx_data[1] , n58968, n29040, n69042, n29653, 
            n27295, \o_Rx_DV_N_3488[12] , n4894, \o_Rx_DV_N_3488[24] , 
            n29, n23, n61278, n6, tx_enable, baudrate, r_Clock_Count_adj_22, 
            n25117, \o_Rx_DV_N_3488[8] , \r_SM_Main[2]_adj_19 , \o_Rx_DV_N_3488[7] , 
            r_Rx_Data, RX_N_2, \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , n4891, \r_Bit_Index[0]_adj_20 , 
            \r_SM_Main[1]_adj_21 , n58022, n27288, n58970, n61676, 
            n61604, n61658, n61640, n61586, n61622, n61550, n29912, 
            n29911, n29910, n29909, n29908, n29907, n29906, n29663, 
            n54370, n29667, n27292, n61568, n61280) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_in_frame[5] ;
    input n3014;
    output [7:0]\data_out_frame[18] ;
    input clk16MHz;
    input n57886;
    input n58004;
    input n29483;
    input VCC_net;
    output [7:0]\data_in_frame[15] ;
    input n57892;
    input n57893;
    input n57885;
    input n29480;
    input n57884;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[6] ;
    input n57894;
    input n57883;
    output [7:0]\data_out_frame[19] ;
    input n57882;
    input n57881;
    input n57880;
    input n57879;
    output [7:0]\data_out_frame[23] ;
    input GND_net;
    output [7:0]\data_in_frame[3] ;
    input n57878;
    output \data_out_frame[1][6] ;
    input n57996;
    output \data_out_frame[1][7] ;
    input n57995;
    input n57877;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_out_frame[17] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]pwm_setpoint;
    input n57876;
    input n57875;
    output [7:0]\data_out_frame[20] ;
    input n57874;
    input n57873;
    output n25488;
    input n57872;
    input n57871;
    output [7:0]\data_in_frame[14] ;
    output [7:0]\data_in_frame[1] ;
    input n29477;
    input Kp_23__N_869;
    output \data_out_frame[3][1] ;
    input n57994;
    input n57870;
    input n57869;
    input n58867;
    output n58698;
    output n53862;
    output [7:0]\data_out_frame[16] ;
    input n57868;
    input n57867;
    output \data_out_frame[3][3] ;
    input n57993;
    output \data_in_frame[2][5] ;
    input n29474;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[11] ;
    output \data_out_frame[3][4] ;
    input n57992;
    output \data_out_frame[3][6] ;
    input n57991;
    output \data_out_frame[3][7] ;
    input n57990;
    output \data_in_frame[3][4] ;
    input n29471;
    output [7:0]\data_out_frame[4] ;
    input n28927;
    input n57989;
    input n57895;
    output \data_in_frame[5][6] ;
    input n29468;
    input n57988;
    input n57987;
    output [7:0]\data_out_frame[21] ;
    input n57866;
    input n57865;
    input n57864;
    input n57863;
    input n57862;
    input n57861;
    input n57860;
    input n57859;
    output [7:0]\data_out_frame[22] ;
    input n57858;
    input n57857;
    input n57856;
    input n57855;
    input n28782;
    input n57854;
    input n28780;
    input n57853;
    input n57852;
    input n57986;
    input n29465;
    input n57985;
    output n62;
    input n57984;
    output [7:0]\data_out_frame[5] ;
    input n57983;
    input n29462;
    input n57982;
    input n57981;
    input n57980;
    input n29459;
    input n57979;
    input n57978;
    input n57851;
    input n29456;
    input n57977;
    input n29453;
    input n57976;
    input n29450;
    output [7:0]\data_out_frame[6] ;
    input \encoder0_position_scaled[22] ;
    input n57975;
    input n29447;
    input n57974;
    input n29444;
    input n28909;
    input n57850;
    input n57849;
    input n57848;
    input n57847;
    input n28772;
    input n57896;
    output [7:0]\data_out_frame[24] ;
    input n57846;
    input n57845;
    input n28768;
    input n28767;
    input n57844;
    input n57843;
    input n28764;
    input n57842;
    output [7:0]\data_out_frame[25] ;
    input n57841;
    input n57840;
    input n57839;
    input n57838;
    input n57837;
    input n57836;
    input n57835;
    input n57973;
    input n29441;
    input n57834;
    output [23:0]neopxl_color;
    output n22373;
    output n58391;
    output \data_in_frame[3][3] ;
    output \data_in_frame[5][3] ;
    input n11;
    input n12;
    output [7:0]\data_in_frame[20] ;
    input n29438;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[21] ;
    output \data_in_frame[23][2] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_out_frame[15] ;
    output \data_in_frame[23][6] ;
    output [7:0]\data_in_frame[16] ;
    output \data_in_frame[20][1] ;
    input n57972;
    output \data_in_frame[3][0] ;
    output \data_in_frame[5][2] ;
    input n57971;
    output \data_in_frame[23][1] ;
    output \data_in_frame[23][7] ;
    output \data_in_frame[23][0] ;
    output \data_in_frame[20][5] ;
    input reset;
    output \data_in_frame[5][0] ;
    input n29435;
    output [23:0]setpoint;
    output \data_in_frame[20][6] ;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_in_frame[12] ;
    output \data_in_frame[3][2] ;
    input n57970;
    output \data_in_frame[16][5] ;
    output \data_in_frame[16][4] ;
    output \byte_transmit_counter[0] ;
    output \data_out_frame[0][2] ;
    input n29432;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_in_frame[17] ;
    input n29429;
    input n57969;
    output [7:0]\data_out_frame[14] ;
    input n29426;
    input n57968;
    input n29423;
    input n57967;
    output [7:0]rx_data;
    output n7;
    output [7:0]\data_out_frame[13] ;
    input n29420;
    input n29417;
    input n29414;
    input n57966;
    input n29411;
    input n29408;
    input n29405;
    output n68861;
    output n68855;
    output \FRAME_MATCHER.state[3] ;
    input n29402;
    input n57965;
    output [7:0]\data_out_frame[12] ;
    input [23:0]displacement;
    input \encoder0_position_scaled[21] ;
    input n29399;
    output \data_in_frame[17][0] ;
    output [23:0]PWMLimit;
    input n29395;
    input n57964;
    input n29392;
    output [7:0]\data_out_frame[11] ;
    input [23:0]encoder1_position_scaled;
    input n29389;
    input n29386;
    output n27924;
    output \data_in_frame[16][7] ;
    output n28009;
    input n29383;
    input n29380;
    output n68849;
    input n29377;
    output [7:0]\data_out_frame[10] ;
    input n29374;
    input \encoder0_position_scaled[20] ;
    input n29371;
    input n29368;
    input n29365;
    input n29362;
    input n29359;
    output [7:0]\data_out_frame[9] ;
    input n57963;
    input n29356;
    input n29353;
    input n29350;
    input n29347;
    input n29344;
    input n29341;
    input n29338;
    input n29335;
    input n29332;
    input n29329;
    input n29326;
    input n29323;
    input n29320;
    input n29317;
    input n29314;
    input n29311;
    input n29308;
    input n29305;
    output \data_out_frame[1][5] ;
    input n29302;
    input n29299;
    output \data_out_frame[1][3] ;
    input n29296;
    output \data_out_frame[1][1] ;
    input n57832;
    output \data_out_frame[1][0] ;
    output \data_out_frame[0][4] ;
    output \data_out_frame[0][3] ;
    input n29107;
    input n29110;
    input n29113;
    input n57504;
    input n29165;
    input n29184;
    input n29188;
    input n29191;
    input n29194;
    input n29206;
    input n29209;
    input n57962;
    output \data_out_frame[8][3] ;
    input n57961;
    output \data_out_frame[8][4] ;
    input n57960;
    output \data_out_frame[8][5] ;
    input n57959;
    output \data_out_frame[8][6] ;
    input n57958;
    output \data_out_frame[8][7] ;
    input n57957;
    output rx_data_ready;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output n68783;
    input \encoder0_position_scaled[7] ;
    input \encoder0_position_scaled[6] ;
    input \encoder0_position_scaled[5] ;
    input \encoder0_position_scaled[4] ;
    input \encoder0_position_scaled[3] ;
    input \encoder0_position_scaled[15] ;
    input n58003;
    input n58002;
    input n58001;
    input n58000;
    input n57999;
    input n57998;
    input n57997;
    input n57956;
    input n57955;
    input n26;
    input n57954;
    input n57953;
    input n57952;
    input n57951;
    input n57950;
    input n57949;
    input n57948;
    input n57947;
    input n57946;
    input n57945;
    input n57944;
    input n57943;
    input n57942;
    input n57941;
    input n57940;
    input n57939;
    input n57938;
    input n57937;
    input n57936;
    input n57935;
    input n57934;
    input n57933;
    input n57932;
    input n57931;
    input n57930;
    input n57929;
    input n57928;
    input n57927;
    input n57926;
    input n57925;
    input n57924;
    input n57923;
    input n57922;
    input n57921;
    input n57920;
    input n57919;
    input n57918;
    input n57917;
    input n57916;
    input n57915;
    input n57914;
    input n57913;
    input n57912;
    input n57911;
    input n57898;
    input n57910;
    input n57909;
    input n57908;
    input n57897;
    input n28838;
    input n28837;
    input n57907;
    input n57906;
    input n57904;
    input n57905;
    input n57833;
    input n28831;
    input n57903;
    input n57902;
    input n57901;
    input n28827;
    input n57900;
    input n28825;
    input n57899;
    input n57891;
    input n57890;
    output LED_c;
    input n29052;
    output n22362;
    output n58147;
    output n27920;
    output DE_c;
    input n57889;
    input n29018;
    output [15:0]current_limit;
    input n29017;
    output [7:0]control_mode;
    input n29016;
    output n58819;
    output \Ki[0] ;
    output n10;
    output n38;
    output n27972;
    input n1510;
    input n10_adj_6;
    input n58707;
    input n58653;
    input n2076;
    input n57888;
    input n29486;
    output n27600;
    input n363;
    output n35;
    input n29495;
    input n29498;
    input n28969;
    input n28972;
    input n29501;
    input n29504;
    input n28976;
    input n28979;
    input n29507;
    input n29510;
    input n57380;
    input n29516;
    input n57378;
    input n28982;
    input n57376;
    input n57374;
    input n57372;
    input n57370;
    input n29593;
    input n29599;
    input n29602;
    input n29605;
    input n29608;
    input n29951;
    input n29948;
    input n29945;
    input n29942;
    output \Kp[0] ;
    input n28987;
    input n57356;
    input n57354;
    input n57350;
    input n57346;
    input n29704;
    input n28993;
    output \data_in_frame[2][3] ;
    input n29000;
    output [23:0]deadband;
    output [23:0]IntegralLimit;
    output \Kp[1] ;
    output \Kp[2] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output \Kp[5] ;
    output \Kp[6] ;
    output \Kp[7] ;
    output \Kp[8] ;
    output \Kp[9] ;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    output \Kp[13] ;
    output \Kp[14] ;
    output \Kp[15] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    output \Ki[14] ;
    output \Ki[15] ;
    input n29778;
    input n29777;
    input n29776;
    input n29775;
    input n29774;
    input n29773;
    input n29772;
    input n29771;
    input n29770;
    input n29769;
    input n29768;
    input n29767;
    input n29765;
    input n29763;
    input n29762;
    input n29761;
    input n29760;
    input n29759;
    input n29758;
    input n29757;
    input n29756;
    input n29755;
    input n29754;
    input n29753;
    input n29752;
    input n29751;
    input n29750;
    input n29749;
    input n29748;
    input n29747;
    input n29745;
    input n29744;
    input n29743;
    input n29742;
    input n29740;
    input n29739;
    input n29738;
    input n29737;
    input n29736;
    input n29735;
    input n57887;
    input n29009;
    input n29013;
    input n29020;
    input n29024;
    input n29028;
    output n7_adj_7;
    input n29044;
    output n27968;
    input \encoder0_position_scaled[14] ;
    input n53279;
    output n28002;
    output n53121;
    output n58777;
    output tx_active;
    input n58922;
    output n1130;
    output n58644;
    input \encoder0_position_scaled[13] ;
    input n58225;
    input n58436;
    output n58919;
    input n58245;
    input n25237;
    output n25996;
    input n58312;
    output n58828;
    output n58446;
    input n58680;
    output n27997;
    output n27994;
    output n58835;
    output n1191;
    output n58845;
    input n58276;
    input n58742;
    input n58321;
    input n25269;
    input n58925;
    input n58857;
    output n58363;
    input n58608;
    output n26180;
    input \encoder0_position_scaled[19] ;
    input \encoder0_position_scaled[18] ;
    input \encoder0_position_scaled[17] ;
    input \encoder0_position_scaled[16] ;
    input \encoder0_position_scaled[12] ;
    input \current[15] ;
    input n30;
    output n296;
    input \encoder0_position_scaled[11] ;
    input [7:0]ID;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \encoder0_position_scaled[10] ;
    input \current[0] ;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input \encoder0_position_scaled[9] ;
    input \encoder0_position_scaled[8] ;
    input \encoder0_position_scaled[23] ;
    input n21;
    input n19;
    input n20;
    output n58143;
    output n58632;
    output n68699;
    output n58142;
    input n53;
    output n58141;
    input n58185;
    input n53988;
    output n68675;
    output n68663;
    output n58140;
    output n58144;
    output n58145;
    output n58139;
    output n60939;
    output n68639;
    input n62904;
    input n62902;
    output n7_adj_8;
    output n7_adj_9;
    output n7_adj_10;
    input n1828;
    input n209;
    output n270;
    output n68633;
    output [8:0]r_Clock_Count;
    output n1;
    output tx_o;
    output [2:0]r_SM_Main;
    output \r_Bit_Index[0] ;
    output n27;
    input \tx_data[6] ;
    input \tx_data[3] ;
    input \tx_data[2] ;
    input \tx_data[1] ;
    output n58968;
    input n29040;
    input n69042;
    input n29653;
    output n27295;
    output \o_Rx_DV_N_3488[12] ;
    input n4894;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    output n61278;
    output n6;
    output tx_enable;
    input [31:0]baudrate;
    output [7:0]r_Clock_Count_adj_22;
    output n25117;
    output \o_Rx_DV_N_3488[8] ;
    output \r_SM_Main[2]_adj_19 ;
    output \o_Rx_DV_N_3488[7] ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    input n4891;
    output \r_Bit_Index[0]_adj_20 ;
    output \r_SM_Main[1]_adj_21 ;
    input n58022;
    output n27288;
    output n58970;
    output n61676;
    output n61604;
    output n61658;
    output n61640;
    output n61586;
    output n61622;
    output n61550;
    input n29912;
    input n29911;
    input n29910;
    input n29909;
    input n29908;
    input n29907;
    input n29906;
    input n29663;
    input n54370;
    input n29667;
    output n27292;
    output n61568;
    output n61280;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n58730, n58409, n26031, n2, n2_adj_5283, n2_adj_5284, n2_adj_5285, 
        n2_adj_5286, n2_adj_5287, n6_c, Kp_23__N_875, n25908, n58173, 
        n2_adj_5288, n2_adj_5289, n2_adj_5290, n2_adj_5291, n2_adj_5292, 
        n2_adj_5293, n53191, n25947, n58539, n25963, n2_adj_5294, 
        n2_adj_5295, n58327, n10_c, n2_adj_5296, n2_adj_5297, n26388, 
        n25497, n3;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5298, n58620, n25871, n6_adj_5299, n25426, n2_adj_5300, 
        n2_adj_5301, n2_adj_5302, n2_adj_5303;
    wire [7:0]\data_in_frame[5]_c ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58267, n2_adj_5304, n2_adj_5305, n25280, n58468, n10_adj_5306, 
        n58677;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n58300, Kp_23__N_993, n7_c, n4, n58873, n58285, n25405, 
        Kp_23__N_872, n25476, n25511, n2_adj_5307, n2_adj_5308, n2_adj_5309, 
        n2_adj_5310, n58340, n25503, n58565, n25479, n25923, n58182, 
        n2_adj_5311, n2_adj_5312, n2_adj_5313, n2_adj_5314, n58337, 
        n58534, n25319, n58162, n25466, n2_adj_5315;
    wire [7:0]\data_in_frame[2]_c ;   // verilog/coms.v(99[12:25])
    
    wire n25448, n58282, n58330, n58674, n62210, n2_adj_5316, n26297, 
        n58822, n58179, n58279, n58545, n2_adj_5317, n2_adj_5318, 
        Kp_23__N_748, n2_adj_5319, n2_adj_5320, n2_adj_5321, n2_adj_5322, 
        n2_adj_5323, n58455, n2_adj_5324, n25936, n2_adj_5325, n2_adj_5326, 
        n2_adj_5327, n2_adj_5328, n2_adj_5329, n2_adj_5330, n2_adj_5331, 
        n2_adj_5332, n2_adj_5333, n2_adj_5334, n2_adj_5335, n2_adj_5336, 
        n2_adj_5337, n2_adj_5338, n2_adj_5339, n2_adj_5340, n2_adj_5341, 
        n58548, n2_adj_5342, n2_adj_5343, n2_adj_5344;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n39291, n65543, n2_adj_5345, n2_adj_5346, n2_adj_5347, n2_adj_5348, 
        n2_adj_5349, n2_adj_5350, n2_adj_5351, n2_adj_5352, n58352, 
        n2_adj_5353, n2_adj_5354, n2_adj_5355, n2_adj_5356, n2_adj_5357, 
        n2_adj_5358, n2_adj_5359, n2_adj_5360, n2_adj_5361, n2_adj_5362, 
        n2_adj_5363, n2_adj_5364, n2_adj_5365, n2_adj_5366, n2_adj_5367, 
        n2_adj_5368, n2_adj_5369, n2_adj_5370, n2_adj_5371, n2_adj_5372, 
        n2_adj_5373, n2_adj_5374, n2_adj_5375, n2_adj_5376, n2_adj_5377, 
        n2_adj_5378, n2_adj_5379, n2_adj_5380, n2_adj_5381, n58659, 
        n29764, n3_adj_5382;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n58017, n3_adj_5383, n58016, n3_adj_5384, n58015, n62300, 
        n2_adj_5385, n3_adj_5386, n58018, n58219, n62306, n58692, 
        n60869, n60943, n29766, n3_adj_5387, n58014, n58359, n53274, 
        n14, n60269, n62641, n20_c, n53770, n62639, n25859, n62494, 
        n25569, n53463, n33, n25549, n7_adj_5388, n32797;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    
    wire n58765, n8, n23480, n60337, n2_adj_5389, n3_adj_5390, n58009, 
        n58554, n58801;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n60508, n24730, n53067, n10_adj_5391, n2_adj_5392, n60682, 
        n62116, n25649, n62118, n53135, n60506, n58374, n6_adj_5393, 
        n60137, n58465, Kp_23__N_1080, n3_adj_5394, n58007, n2_adj_5395, 
        n60685, n26043, n53398, n62124;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    
    wire n10_adj_5396, n58427, n62126, Kp_23__N_974, n62314, n3_adj_5397, 
        n58021, n3_adj_5398;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n58008, n58780, n62434, Kp_23__N_1551, n54291, n62128, 
        n2_adj_5399, n58739, n62130;
    wire [7:0]\data_in_frame[20]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58514, n58891, n60934, n3_adj_5400, n58011, n2_adj_5401, 
        n62322, n62328, n58297, n58200, n58717, n62332, n2_adj_5402, 
        n3_adj_5403, n58012, n58934, n58158, n58810, n62338, n58472, 
        n54148, n58596, n62344, n53903, n58727, n58897, n62350, 
        n3_adj_5404, n58019, n60820, n62160, n23529, n53904, n2_adj_5405, 
        n62376, n58430, n54226, n62392, n59916, n62388, n25604, 
        n60174, n58394, n62134, n3_adj_5406, n58013, n58388, n58724, 
        n58876, n54203, n60227, n58542, n58248, n53374, n3_adj_5407, 
        n58006, n58711, n60149, n3_adj_5408, n58010, n58383, n62146, 
        n24756, n58452, n3_adj_5409, n58020, n2209, Kp_23__N_1748, 
        n69245, n62140, n30_c;
    wire [23:0]n4793;
    
    wire n27308, n2_adj_5410, n58854, n58303, n12_adj_5411, n13, 
        n54274, n1_c, n57823, n62154, n53063, n26158, n25944, 
        n62236, n58768, n58910, n58798, Kp_23__N_1389, n62248, n1_adj_5412, 
        n57825, n1_adj_5413, n57824, n25726, n62246, n58928, Kp_23__N_654, 
        n58324, n62252, n58946, n58459, n58813, n62258, n58879, 
        n62264, n54180, n62272, n58349, n60010, n58759, n62278, 
        n25343, n54184, n58816, n62284, n1_adj_5414, n57826, n53879, 
        n54154;
    wire [7:0]\data_in_frame[16]_c ;   // verilog/coms.v(99[12:25])
    
    wire n1_adj_5415;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n57821, \FRAME_MATCHER.i_31__N_2513 , n1_adj_5416, n57822, 
        n53171, n60815, n53071, n62170, n53772, n62398, n24742, 
        n65539, n2_adj_5417, n62876, n62877, n62404, n62875, n58668, 
        n58885, n62410, n53102, n58913, n54173, n1_adj_5418, n57827, 
        n62456, n58870, n58787, n58671, n54284, n58574, n25437, 
        n2_adj_5419, n58588, n59932, n25544, n2_adj_5420, n25363, 
        Kp_23__N_669, n62448, n53187, n60197, n25525, n62220, n2_adj_5421, 
        n2_adj_5422, n51254, n57819, n26055, n53703, n25538, n2_adj_5423, 
        n62150, n58194, n62222, n58346, n53096, n62360, n25596, 
        n51253, n2_adj_5424, n58825, n62182, n51252, n58851, n62188, 
        n62192, n58424, n62198, n58958, n58551, n58931, n62204, 
        n60751, n2_adj_5425, n51251, n2_adj_5426, n2_adj_5427, n44, 
        n58701, n10_adj_5428, Kp_23__N_878, n42, n2_adj_5429, n58571, 
        n60574, n43;
    wire [7:0]\data_in_frame[17]_c ;   // verilog/coms.v(99[12:25])
    
    wire n41, n40, n58955, n2_adj_5430, n39, n50, n45, n25154, 
        n4452, n2_adj_5431, n2_adj_5432, \FRAME_MATCHER.i_31__N_2514 , 
        n6_adj_5433, n25757, n6_adj_5434, n2_adj_5435, n57446, Kp_23__N_1271, 
        n2_adj_5437, n24758, n2_adj_5438, n2_adj_5439, n2_adj_5440, 
        n11_adj_5441, n12_adj_5442, n68858, n2_adj_5443, n2_adj_5444, 
        n2_adj_5445, n53130, n2_adj_5446, n58695, n6_adj_5447, n60436, 
        n12_adj_5448, n51250, n58228, n28, n2_adj_5449, n51249, 
        n26_c, n27_c, n58270, n25, n9, n65440, n11_adj_5450, n12_adj_5451, 
        n68852, n9_adj_5452, n65441, n69037, \FRAME_MATCHER.i_31__N_2507 , 
        n51248, n58552, n58656, n26617, \FRAME_MATCHER.i_31__N_2508 , 
        n2189, n2190, n57820, tx_transmit_N_3416, n20741, \FRAME_MATCHER.i_31__N_2511 , 
        n57202, \FRAME_MATCHER.i_31__N_2512 , n2201, n27160, n2_adj_5453, 
        n2_adj_5454, n25729, n2_adj_5455, n2_adj_5456, n57444, n4_adj_5457, 
        n5, n68846, n53179, n6_adj_5458, n60509, n58433, n58906, 
        n58484, n54307, n22, n58900, n58421, n58665, n26424, n24, 
        n58804, n58254, n58943, n23_c, n25_adj_5459, n54144, n25462, 
        n54138, n53925, n58499, n2_adj_5460, n27700, n27913, n52061, 
        n65372, n27698, n52060, n65373, n58864, n57424, n2_adj_5461, 
        n58400, n27696, n52059, n65374, n2_adj_5462, n57442, n2_adj_5463, 
        n12_adj_5464, n58599, n58531, n2_adj_5465, n27694, n52058, 
        n65379, n29398, n58291, n12_adj_5466, n27692, n52057, n65382, 
        n2_adj_5467, n27690, n52056, n65386, n2_adj_5468, n27688, 
        n52055, n65387, n25441, n27686, n52054, n65393, n27684, 
        n52053, n65394, n27682, n52052, n65395, n27680, n52051, 
        n65398, n2_adj_5469, n27678, n52050, n65399, n38036, n27676, 
        n52049, n65400, n6_adj_5470, n29864, n10_adj_5471, n27674, 
        n52048, n65401, n2_adj_5472, n58520, n57300, n27672, n52047, 
        n65428, n6_adj_5473, n27670, n52046, n65451, n27668, n52045, 
        n65465, n57302, n54156, n2_adj_5474, n27666, n52044, n65476;
    wire [7:0]\data_in_frame[21]_c ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5475, n27664, n52043, n65479, n7_adj_5476, n25370, 
        n26225, n8_adj_5477, n27662, n52042, n65480, n27660, n52041, 
        n65481, n65442, n1_adj_5478, n2_adj_5479, n27658, n52040, 
        n65482, n27656, n52039, n65487, n38022, n4_adj_5480, n5_adj_5481, 
        n68840, n65444, n65443, n68843, n68828, n68831, n68822, 
        n2_adj_5482, n68825, n27654, n52038, n65489, n27652, n52037, 
        n65491, n27650, n52036, n65495, n2_adj_5483, n2_adj_5484, 
        n68816, n2_adj_5485, n34, n54235, n58582, n8_adj_5486, n27648, 
        n52035, n65499, n27646, n52034, n65500, n27644, n52033, 
        n65501, n2_adj_5487, n58294, n12_adj_5488, n8_adj_5489, n2_adj_5490, 
        n27642, n52032, n65503, n27640, n52031, n65506, n2_adj_5491, 
        n6_adj_5492;
    wire [31:0]n133;
    
    wire n161, n58794, n58315, n54146, n58207, n10_adj_5493, n58527, 
        n68374, n58961, n43_adj_5494, n14_adj_5495, n2_adj_5496, n25645, 
        n58937, n58791, n25845, n13_adj_5497, n53247, n68380, n58212, 
        n2_adj_5498, n2_adj_5499, n2_adj_5500, n10_adj_5501, n58882, 
        n2_adj_5502, n2_adj_5503, n60532, n6_adj_5504, n58848, n15, 
        n2_adj_5505, n2_adj_5506, n2_adj_5507, n68819, n58288, n14_adj_5508, 
        n2_adj_5509, n2_adj_5510, n2_adj_5511, n11_adj_5512, n54197, 
        n58380, n2_adj_5513, n2_adj_5514, n2_adj_5515, n29293, n29290, 
        n29287, n29284, n29281, n2_adj_5516, n2_adj_5517, n29278, 
        n54150, n6_adj_5518, n29275, n8_adj_5519, n27926, n29272, 
        n29269, n29266, n29263, n29260, n2_adj_5520, n29087, n2_adj_5521, 
        n2_adj_5522, n57510, n57494, n68810, n68813, n2_adj_5523, 
        n68804, n68807, n68798, n29212, n57514, n57520, n29221, 
        n29231, n68801, n29224, n29227, n2_adj_5524, n2_adj_5525, 
        n2_adj_5526, n2_adj_5527, n2_adj_5528, n27592, n2_adj_5529, 
        n62873, n62874, n68780, n62872, n3579, n58121, n10_adj_5530, 
        n58133, n10_adj_5531, n58118, n68750, n53055, n60075, n53790, 
        n6_adj_5532, n53666, n58478, n2_adj_5534, n2_adj_5535, n29086;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n68753, n28540, n62621, n29085, n29084, n29083, n29082, 
        n29081, n29080, n2_adj_5536, n29079;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n29078, n68744, n26862, n24_adj_5537, n28536, n29077, n68747, 
        n29076, n29075, n29074, n29073, n29072, n29071;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n29070, n29069, n29068, n27612, n29067, n29066, n29065, 
        n1_adj_5538;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n29064, n29063;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n5_adj_5539, n29062, n29061, n29060, n29059, n29058, n29057, 
        n29056, n11_adj_5540, n12_adj_5541, n69014, n29041, n58418, 
        n58146, n53119, n58736, n10_adj_5542, n26494, n28471, n2_adj_5543, 
        n32799, n6_adj_5544, n29019, n58903, n53169, n58940, n6_adj_5545, 
        n58714, n1_adj_5546, n58916, n42_adj_5547, n58784, n53283, 
        n54293, n40_adj_5548, n41_adj_5549, n58462, n54278, n39_adj_5550, 
        n58689, n38_c, n60272, n58778, n43_adj_5551, n48, n29012, 
        n47, n8_adj_5552, n27918, n58197, n58626, n25656, n58318, 
        n58306, n58397, n58511, n58398, n25814, n23340, n54259, 
        n58370, n58561, n1699, n58774, n58502, n26202, n53164, 
        n58491, n25797, n6_adj_5556, n1673, n58475, n58629, n16, 
        n58166, n58635, n58683, n58579, n17, n58231, n60061, n54182, 
        n1513, n14_adj_5557, n24670, n25666, n15_adj_5558, n59852, 
        n58495, n25830, n16_adj_5559, n27916, n771, n25082, n62488, 
        n26431, n58733, n17_adj_5560, n58771, n25992, n58443, n14_adj_5561, 
        n58647, n13_adj_5562, n60254, n22_adj_5563, n54243, n26199, 
        n20_adj_5564, n2107, n58686, n26288, n21_c, n19_c, n58602, 
        n58807, n63004, n63005, n63002, n63001, n62845, n62846, 
        n62864, n9_adj_5565, n65490, n62994, n62863, n62851, n62852, 
        n68732, n2_adj_5566, n62837, n62836, n62857, n62858, n25800, 
        n62813, n2217, n62812, n62900, n27707, n62901, n62899, 
        n68693, n65478, n67527, n68615, n65546, n67533, n62866, 
        n62867, n62888, n54224, n14_adj_5567, n62889, n62887, n58568, 
        n58377, n10_adj_5568, n68735, n65559, n67535, n62918, n62917, 
        n58412, n65591, n69005, n67569, n31, n57608, n57330, n29537, 
        n57450, n57430, n29546, n57436, n29552, n29555, n57448, 
        n29561, n29564, n29567, n29570, n29577, n57482, n29584, 
        n29587, n57292, n57304, n57288, n29939, n29936, n28999, 
        n29933, n29930, n29927, n29924, n29921, n8_adj_5569, n29614, 
        n29617, n29620, n33_adj_5570, n57414, n29630, n29633, n29638, 
        n29641, n29644, n29648, n29655, n29658, n57420, n29671, 
        n29674, n29677, n29855, n29854, n29853, n29852, n29851, 
        n29850, n29849, n29848, n29847, n29846, n29845, n29844, 
        n29843, n29842, n29841, n29840, n29839, n29838, n29837, 
        n29836, n29835, n29834, n29832, n29831, n29830, n29829, 
        n29828, n29827, n29826, n29825, n29824, n29823, n29822, 
        n29821, n29820, n29819, n29818, n29817, n29816, n29815, 
        n29814, n29813, n29812, n29811, n29810, n29809, n29808, 
        n29807, n29806, n29805, n29804, n29803, n29802, n29801, 
        n29800, n29799, n29798, n29797, n29796, n29795, n29794, 
        n29793, n29792, n29791, n29790, n29789, n29788, n29787, 
        n29786, n29785, n29784, n29783, n29782, n29781, n29780, 
        n29779, n29746, n29741, n29734;
    wire [15:0]current_limit_c;   // verilog/TinyFPGA_B.v(251[22:35])
    
    wire n29733, n29732, n29731, n29730, n29729, n29728, n29727, 
        n29726, n29725, n29724, n29723, n29722, n29721, n29720, 
        n29719, n29718, n29717, n2_adj_5571, n29716, n29715, n29714, 
        n29713, n29712, n53880, n22_adj_5572, n60594, n16_adj_5573, 
        n24_adj_5574, n20_adj_5575, n58222, n10_adj_5576, n8_adj_5578, 
        n28986, n29580, n28985, n2095, n2092, n2098, n60080, n58894, 
        n6_adj_5579, n7_adj_5580, n54324, n58641, n10_adj_5581, n54253, 
        n53721, n8_adj_5582, n12_adj_5583, n23344, n58623, n8_adj_5584, 
        n6_adj_5585, n5_adj_5586, n58605, n39337, n58273, n58949, 
        n58662, n58614, n53285, n40_adj_5587, n54237, n10_adj_5588, 
        n53999, n58440, n26088, n58638, n25673, n26235, n58704, 
        n12_adj_5589, n24827, n58838, n10_adj_5590, n25763, n58650, 
        n58242, n8_adj_5591, n4_adj_5592, n28_adj_5593, n58449, n58189, 
        n26_adj_5594, n27_adj_5595, n25_adj_5596, n25663, n6_adj_5597, 
        n60866, n60941, n10_adj_5598, n14_adj_5599, n10_adj_5600, 
        n58343, n10_adj_5601, n7_adj_5602, n5_adj_5603, n25456, n26100, 
        n1312, n26085, n25639, n10_adj_5604, n25335, n14_adj_5605, 
        n58585, n58216, n25259, n15_adj_5606, n14_adj_5607, n22_adj_5608, 
        n34_adj_5609, n23_adj_5610, n38_adj_5611, n58562, n58258, 
        n36, n37, n58617, n35_adj_5612, n12_adj_5613, n60872, n10_adj_5614, 
        n58151, n25377, n25301, n6_adj_5615, n6_adj_5616, n58611, 
        n26330, n7_adj_5617, n60003, n20750, n22366, n3303, n62469, 
        n60217, n2096, n25001, n26612, n60942, n25090, n10_adj_5619, 
        n14_adj_5620, n25127, n20_adj_5621, n25029, n19_adj_5622, 
        n62651, n25157, n18, n25096, n20_adj_5623, n15_adj_5624, 
        n10_adj_5625, n16_adj_5626, n17_adj_5627, n14_adj_5628, n15_adj_5629, 
        n16_adj_5630, n17_adj_5631, n38817, n4_adj_5632, n4_adj_5633, 
        n6_adj_5634, n27598, n62894, n62895, n62893, n69002, n68996, 
        n10_adj_5638, n68711;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n68708, n12_adj_5639, n68984, n10_adj_5640, n68681, n7_adj_5641, 
        n58108, n10_adj_5642, n68978, n68669, n7_adj_5643, n68696, 
        n11_adj_5644, n68972, n68690, n7_adj_5645, n9_adj_5646, n23_adj_5647, 
        n26_adj_5648, n29_c, n32809, n68678, n22_adj_5649, n68672, 
        n32, n58092, n68666, n68660, n68636, n68630, n68612, n27_adj_5653, 
        n57758, n61290;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n59805;
    
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[7] [2]), .I1(n58730), .I2(n58409), 
            .I3(\data_in_frame[5] [1]), .O(n26031));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2), .S(n57886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5283), .S(n58004));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29483));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5284), .S(n57892));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5285), .S(n57893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5286), .S(n57885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29480));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5287), .S(n57884));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[4] [3]), .I3(n6_c), .O(Kp_23__N_875));   // verilog/coms.v(76[16:42])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1109 (.I0(\data_in_frame[4] [6]), .I1(n25908), 
            .I2(\data_in_frame[6] [6]), .I3(\data_in_frame[7] [0]), .O(n58173));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5288), .S(n57894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5289), .S(n57883));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5290), .S(n57882));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5291), .S(n57881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5292), .S(n57880));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5293), .S(n57879));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n53191), .I1(\data_out_frame[23] [3]), .I2(n25947), 
            .I3(GND_net), .O(n58539));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i14_2_lut (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n25963));   // verilog/coms.v(99[12:25])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5294), .S(n57878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5295), .S(n57996));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1110 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [4]), 
            .I2(\data_in_frame[7] [5]), .I3(n58327), .O(n10_c));
    defparam i4_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5296), .S(n57995));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5297), .S(n57877));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[8] [2]), .I1(n26388), .I2(n25497), 
            .I3(GND_net), .O(n3));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5298));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut (.I0(n58173), .I1(n58620), .I2(GND_net), .I3(GND_net), 
            .O(n25871));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1111 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8] [5]), 
            .I2(\data_in_frame[6] [3]), .I3(n6_adj_5299), .O(n25426));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5300), .S(n57876));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5301), .S(n57875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5302), .S(n57874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5303), .S(n57873));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1112 (.I0(\data_in_frame[5]_c [7]), .I1(\data_in_frame[3]_c [7]), 
            .I2(n25488), .I3(\data_in_frame[6] [1]), .O(n58267));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5304), .S(n57872));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5305), .S(n57871));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(n25280), .I1(n58468), .I2(n10_adj_5306), 
            .I3(\data_in_frame[14] [2]), .O(n58677));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58300));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29477));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), .I2(GND_net), 
            .I3(GND_net), .O(n7_c));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1114 (.I0(n25497), .I1(Kp_23__N_869), .I2(\data_in_frame[6] [2]), 
            .I3(\data_in_frame[8] [3]), .O(n4));   // verilog/coms.v(239[9:81])
    defparam i3_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1115 (.I0(\data_in_frame[0] [0]), .I1(n58873), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n58285));
    defparam i2_3_lut_adj_1115.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25488));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(n25405), .I1(n58285), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1118 (.I0(n25476), .I1(Kp_23__N_872), .I2(Kp_23__N_869), 
            .I3(\data_in_frame[8] [4]), .O(n25511));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25476));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5307));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5308), .S(n57994));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5309), .S(n57870));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5310), .S(n57869));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1120 (.I0(\data_in_frame[6] [0]), .I1(n58867), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(n58340));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1120.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut (.I0(n58698), .I1(n53862), .I2(n58340), .I3(n25503), 
            .O(n58565));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1121 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[5]_c [5]), 
            .I2(n25479), .I3(n25923), .O(n58182));
    defparam i3_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5312), .S(n57868));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5313), .S(n57867));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5314), .S(n57993));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1122 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58337));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[5]_c [5]), .I1(n58534), 
            .I2(GND_net), .I3(GND_net), .O(n25319));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1124 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58162));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25466));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5315));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_in_frame[2]_c [7]), .I1(n25448), 
            .I2(GND_net), .I3(GND_net), .O(n58282));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2]_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58330));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1128 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3]_c [7]), .I3(GND_net), .O(n58873));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[2] [1]), .I1(n25908), .I2(\data_in_frame[4] [3]), 
            .I3(GND_net), .O(n58674));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[2][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n62210));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29474));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1130 (.I0(n58330), .I1(n58282), .I2(n62210), 
            .I3(\data_in_frame[2]_c [6]), .O(n58730));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[9] [2]), .I1(n26297), .I2(\data_in_frame[11] [4]), 
            .I3(\data_in_frame[14] [7]), .O(n58822));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58179));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58279));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58545));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5317), .S(n57992));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5318), .S(n57991));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1134 (.I0(\data_in_frame[0] [7]), .I1(n58545), 
            .I2(n58279), .I3(n58179), .O(Kp_23__N_748));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5319), .S(n57990));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1135 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3][4] ), .I3(GND_net), .O(n25479));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29471));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5321), .S(n28927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5322), .S(n57989));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5323), .S(n57895));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_in_frame[5][6] ), .I1(n25479), 
            .I2(GND_net), .I3(GND_net), .O(n58455));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29468));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5324), .S(n57988));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1137 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2]_c [2]), .I3(GND_net), .O(n25936));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5325), .S(n57987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5326), .S(n57866));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5327), .S(n57865));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5328), .S(n57864));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5329), .S(n57863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5330), .S(n57862));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5331), .S(n57861));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5332), .S(n57860));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5333), .S(n57859));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5334), .S(n57858));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5335), .S(n57857));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5336), .S(n57856));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5337), .S(n57855));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5338), .S(n28782));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5339), .S(n57854));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5340), .S(n28780));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5341), .S(n57853));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[4] [4]), .I1(n25936), 
            .I2(GND_net), .I3(GND_net), .O(n58548));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5342), .S(n57852));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5343), .S(n57986));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29465));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5344), .S(n57985));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48874_2_lut_3_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n39291), 
            .I2(n62), .I3(GND_net), .O(n65543));
    defparam i48874_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5345), .S(n57984));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5346), .S(n57983));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29462));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5347), .S(n57982));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5348), .S(n57981));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5349), .S(n57980));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29459));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5350), .S(n57979));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5351), .S(n57978));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5352), .S(n57851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29456));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[2] [0]), .I1(Kp_23__N_748), 
            .I2(GND_net), .I3(GND_net), .O(n58352));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5353), .S(n57977));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29453));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5354), .S(n57976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29450));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[22] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5356), .S(n57975));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29447));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5357), .S(n57974));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29444));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5358), .S(n28909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5359), .S(n57850));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5360), .S(n57849));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5361), .S(n57848));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5362), .S(n57847));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5363), .S(n28772));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5364), .S(n57896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5365), .S(n57846));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5366), .S(n57845));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5367), .S(n28768));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5368), .S(n28767));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5369), .S(n57844));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5370), .S(n57843));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5371), .S(n28764));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5372), .S(n57842));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5373), .S(n57841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5374), .S(n57840));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5375), .S(n57839));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5376), .S(n57838));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5377), .S(n57837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5378), .S(n57836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5379), .S(n57835));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5380), .S(n57973));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29441));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5381), .S(n57834));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58659));
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25503));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i18978_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5]_c [7]), 
            .I2(n22373), .I3(GND_net), .O(n29764));
    defparam i18978_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5382), .S(n58017));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1142 (.I0(\data_in_frame[5]_c [7]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3]_c [5]), .I3(GND_net), .O(n58391));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1142.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5383), .S(n58016));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5384), .S(n58015));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1143 (.I0(n25405), .I1(n58659), .I2(\data_in_frame[3]_c [5]), 
            .I3(\data_in_frame[3][3] ), .O(n62300));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5386), .S(n58018));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1144 (.I0(n58352), .I1(n58219), .I2(n62300), 
            .I3(n58548), .O(n62306));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1145 (.I0(n58692), .I1(n58730), .I2(n58674), 
            .I3(n58873), .O(n60869));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1146 (.I0(\data_in_frame[5][3] ), .I1(n25319), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[4] [0]), .O(n60943));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i19034_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5]_c [5]), 
            .I2(n22373), .I3(GND_net), .O(n29766));
    defparam i19034_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5387), .S(n58014));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1147 (.I0(n60943), .I1(n60869), .I2(n58359), 
            .I3(n62306), .O(n53862));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1148 (.I0(n53274), .I1(n58182), .I2(\data_in_frame[8] [0]), 
            .I3(n58565), .O(n14));
    defparam i3_4_lut_adj_1148.LUT_INIT = 16'h1248;
    SB_LUT4 i45634_4_lut (.I0(n25511), .I1(n60269), .I2(n11), .I3(n12), 
            .O(n62641));
    defparam i45634_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i9_4_lut (.I0(n62641), .I1(n4), .I2(n14), .I3(n7_c), .O(n20_c));
    defparam i9_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i45632_4_lut (.I0(n25426), .I1(n25871), .I2(n3), .I3(n53770), 
            .O(n62639));
    defparam i45632_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45490_2_lut (.I0(n25859), .I1(n26031), .I2(GND_net), .I3(GND_net), 
            .O(n62494));
    defparam i45490_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(n25569), .I1(n53463), .I2(n62639), .I3(n20_c), 
            .O(n33));
    defparam i2_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1_4_lut_adj_1149 (.I0(n25549), .I1(n33), .I2(n62494), .I3(n7_adj_5388), 
            .O(n32797));
    defparam i1_4_lut_adj_1149.LUT_INIT = 16'h0008;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[22] [4]), .I1(\data_in_frame[18] [2]), 
            .I2(n58765), .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1150 (.I0(n23480), .I1(n8), .I2(\data_in_frame[20] [2]), 
            .I3(\data_in_frame[20] [3]), .O(n60337));
    defparam i4_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5390), .S(n58009));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1151 (.I0(n58554), .I1(n58801), .I2(\data_in_frame[23] [4]), 
            .I3(GND_net), .O(n60508));
    defparam i2_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29438));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1152 (.I0(n24730), .I1(\data_in_frame[18] [1]), 
            .I2(n53067), .I3(\data_in_frame[20] [4]), .O(n10_adj_5391));
    defparam i4_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1153 (.I0(n60508), .I1(n60682), .I2(n60337), 
            .I3(n60269), .O(n62116));
    defparam i1_4_lut_adj_1153.LUT_INIT = 16'h0008;
    SB_LUT4 i1_4_lut_adj_1154 (.I0(\data_in_frame[21] [1]), .I1(n62116), 
            .I2(\data_in_frame[23][2] ), .I3(n25649), .O(n62118));
    defparam i1_4_lut_adj_1154.LUT_INIT = 16'h4884;
    SB_LUT4 i2_4_lut_adj_1155 (.I0(n53135), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[23] [3]), .I3(n58801), .O(n60506));   // verilog/coms.v(99[12:25])
    defparam i2_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1156 (.I0(\data_in_frame[22] [1]), .I1(\data_in_frame[21] [7]), 
            .I2(n58374), .I3(n6_adj_5393), .O(n60137));
    defparam i4_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1157 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n58465), .I3(n25280), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5394), .S(n58007));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[20] [3]), .I1(n10_adj_5391), .I2(\data_in_frame[22] [5]), 
            .I3(GND_net), .O(n60685));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1158 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n26043), .I3(\data_in_frame[10] [0]), .O(n53398));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1159 (.I0(n60685), .I1(n60137), .I2(n60506), 
            .I3(n62118), .O(n62124));
    defparam i1_4_lut_adj_1159.LUT_INIT = 16'h0400;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[22] [0]), .I3(\data_in_frame[21] [6]), .O(n10_adj_5396));
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1161 (.I0(\data_in_frame[23] [5]), .I1(n62124), 
            .I2(n58427), .I3(n58554), .O(n62126));
    defparam i1_4_lut_adj_1161.LUT_INIT = 16'h8448;
    SB_LUT4 i1_3_lut_4_lut (.I0(n4), .I1(n3), .I2(Kp_23__N_974), .I3(n26297), 
            .O(n62314));   // verilog/coms.v(77[16:43])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5397), .S(n58021));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5398), .S(n58008));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1162 (.I0(n58780), .I1(\data_in_frame[20] [2]), 
            .I2(\data_in_frame[19] [7]), .I3(\data_in_frame[22] [3]), .O(n62434));
    defparam i1_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1163 (.I0(n62126), .I1(Kp_23__N_1551), .I2(n10_adj_5396), 
            .I3(n54291), .O(n62128));
    defparam i1_4_lut_adj_1163.LUT_INIT = 16'h2882;
    SB_LUT4 select_776_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1164 (.I0(n58427), .I1(n62128), .I2(n58739), 
            .I3(\data_in_frame[23][6] ), .O(n62130));
    defparam i1_4_lut_adj_1164.LUT_INIT = 16'h4884;
    SB_LUT4 i2_3_lut_adj_1165 (.I0(\data_in_frame[20]_c [0]), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n58374));
    defparam i2_3_lut_adj_1165.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1166 (.I0(n58514), .I1(n58891), .I2(n58765), 
            .I3(n62434), .O(n60934));
    defparam i1_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5400), .S(n58011));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1167 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[20][1] ), .I3(GND_net), .O(n62322));
    defparam i1_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1168 (.I0(\data_in_frame[20] [2]), .I1(n58374), 
            .I2(n62322), .I3(\data_in_frame[20] [3]), .O(n62328));
    defparam i1_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1169 (.I0(n58297), .I1(n62328), .I2(n58200), 
            .I3(n58717), .O(n62332));
    defparam i1_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5402), .S(n57972));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5403), .S(n58012));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[0] [6]), .I1(n25448), .I2(\data_in_frame[3][0] ), 
            .I3(\data_in_frame[5][2] ), .O(n58692));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1170 (.I0(n58934), .I1(n58158), .I2(n58810), 
            .I3(n62332), .O(n62338));
    defparam i1_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1171 (.I0(n58472), .I1(n54148), .I2(n58596), 
            .I3(n62338), .O(n62344));
    defparam i1_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1172 (.I0(n53903), .I1(n58727), .I2(n58897), 
            .I3(n62344), .O(n62350));
    defparam i1_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5404), .S(n58019));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1173 (.I0(n60820), .I1(n62160), .I2(n23529), 
            .I3(n62350), .O(n53904));
    defparam i1_4_lut_adj_1173.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5405), .S(n57971));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1174 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[21] [7]), 
            .I2(n58801), .I3(GND_net), .O(n62376));
    defparam i1_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1175 (.I0(n58427), .I1(n58430), .I2(n62376), 
            .I3(n58554), .O(n54226));
    defparam i1_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1176 (.I0(n58514), .I1(\data_in_frame[18] [1]), 
            .I2(\data_in_frame[22] [2]), .I3(n58780), .O(n62392));
    defparam i1_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1177 (.I0(n24730), .I1(n59916), .I2(\data_in_frame[19] [6]), 
            .I3(\data_in_frame[20]_c [0]), .O(n62388));
    defparam i1_4_lut_adj_1177.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1178 (.I0(n53903), .I1(n54291), .I2(n59916), 
            .I3(\data_in_frame[19] [5]), .O(n60820));
    defparam i1_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1179 (.I0(n58739), .I1(n60820), .I2(\data_in_frame[21] [6]), 
            .I3(GND_net), .O(n58430));
    defparam i1_3_lut_adj_1179.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1180 (.I0(n4), .I1(n3), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n25604));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1181 (.I0(n54226), .I1(n53904), .I2(n53135), 
            .I3(\data_in_frame[23][1] ), .O(n60174));
    defparam i1_4_lut_adj_1181.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1182 (.I0(\data_in_frame[19] [4]), .I1(n53903), 
            .I2(n58394), .I3(GND_net), .O(n54291));
    defparam i1_3_lut_adj_1182.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1183 (.I0(n60934), .I1(\data_in_frame[23][7] ), 
            .I2(n62130), .I3(n58430), .O(n62134));
    defparam i1_4_lut_adj_1183.LUT_INIT = 16'h2080;
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5406), .S(n58013));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1184 (.I0(n58388), .I1(n58724), .I2(n58876), 
            .I3(n58465), .O(n54203));
    defparam i2_3_lut_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1185 (.I0(n54226), .I1(n25649), .I2(\data_in_frame[23][0] ), 
            .I3(n53904), .O(n60227));
    defparam i1_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1186 (.I0(n58388), .I1(n58724), .I2(n58542), 
            .I3(\data_in_frame[11] [7]), .O(n58248));
    defparam i1_3_lut_4_lut_adj_1186.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1187 (.I0(n58388), .I1(n58724), .I2(Kp_23__N_1080), 
            .I3(GND_net), .O(n53374));
    defparam i1_2_lut_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5407), .S(n58006));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1188 (.I0(n62388), .I1(n62392), .I2(n58891), 
            .I3(n58711), .O(n60149));
    defparam i1_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5408), .S(n58010));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1189 (.I0(n58727), .I1(n58383), .I2(\data_in_frame[20][5] ), 
            .I3(\data_in_frame[22] [7]), .O(n62146));
    defparam i1_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1190 (.I0(n24756), .I1(n54291), .I2(\data_in_frame[21] [5]), 
            .I3(n58452), .O(n58739));
    defparam i1_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n3014), .D(n3_adj_5409), .S(n58020));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2209), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i1_rep_228_2_lut (.I0(n25649), .I1(n53904), .I2(GND_net), 
            .I3(GND_net), .O(n69245));
    defparam i1_rep_228_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1191 (.I0(n60149), .I1(n60227), .I2(n62134), 
            .I3(n60174), .O(n62140));
    defparam i1_4_lut_adj_1191.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1192 (.I0(n62140), .I1(n54226), .I2(n69245), 
            .I3(n62146), .O(n30_c));
    defparam i1_4_lut_adj_1192.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1193 (.I0(\data_in_frame[0] [6]), .I1(n25448), 
            .I2(\data_in_frame[3][0] ), .I3(\data_in_frame[5][0] ), .O(n58409));
    defparam i1_2_lut_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29435));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27308), 
            .D(n4793[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut (.I0(n58854), .I1(n58303), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_5411));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[16] [2]), 
            .I2(\data_in_frame[18] [4]), .I3(\data_in_frame[20][6] ), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n13), .I1(n54274), .I2(n12_adj_5411), .I3(n58677), 
            .O(n25649));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n3014), .D(n1_c), .S(n57823));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1194 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [5]), 
            .I2(n58780), .I3(GND_net), .O(n62154));
    defparam i1_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1195 (.I0(n53063), .I1(n26158), .I2(n25944), 
            .I3(n62154), .O(n62160));
    defparam i1_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1196 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[14] [0]), .I3(\data_in_frame[15] [6]), .O(n62236));
    defparam i1_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1197 (.I0(n58768), .I1(n58910), .I2(n58798), 
            .I3(Kp_23__N_1389), .O(n62248));
    defparam i1_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n3014), .D(n1_adj_5412), .S(n57825));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n3014), .D(n1_adj_5413), .S(n57824));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1198 (.I0(n62236), .I1(n25726), .I2(\data_in_frame[13] [5]), 
            .I3(\data_in_frame[12] [6]), .O(n62246));
    defparam i1_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1199 (.I0(\data_in_frame[1] [1]), .I1(n58337), 
            .I2(\data_in_frame[3][2] ), .I3(\data_in_frame[7] [4]), .O(n58928));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1200 (.I0(n62246), .I1(n62248), .I2(Kp_23__N_654), 
            .I3(n58324), .O(n62252));
    defparam i1_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1201 (.I0(n58946), .I1(n58459), .I2(n58813), 
            .I3(n62252), .O(n62258));
    defparam i1_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1202 (.I0(n58468), .I1(n58822), .I2(n58879), 
            .I3(n62258), .O(n62264));
    defparam i1_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1203 (.I0(n54180), .I1(n25944), .I2(\data_in_frame[16] [6]), 
            .I3(n62264), .O(n62272));
    defparam i1_4_lut_adj_1203.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1204 (.I0(n58349), .I1(n60010), .I2(n58759), 
            .I3(n62272), .O(n62278));
    defparam i1_4_lut_adj_1204.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1205 (.I0(n25343), .I1(n54184), .I2(n58816), 
            .I3(n62278), .O(n62284));
    defparam i1_4_lut_adj_1205.LUT_INIT = 16'h9669;
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n3014), .D(n1_adj_5414), .S(n57826));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5355), .S(n57970));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1206 (.I0(n53879), .I1(n54154), .I2(\data_in_frame[16]_c [0]), 
            .I3(n62284), .O(n53063));
    defparam i1_4_lut_adj_1206.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[16][5] ), .I1(\data_in_frame[16][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n25726));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n3014), .D(n1_adj_5415), .S(n57821));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17063_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n30_c), .I3(n32797), .O(n27308));   // verilog/coms.v(118[11:12])
    defparam i17063_4_lut.LUT_INIT = 16'he420;
    SB_LUT4 i2_3_lut_4_lut_adj_1208 (.I0(n53463), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[12] [1]), .I3(\data_in_frame[9] [7]), .O(n58876));
    defparam i2_3_lut_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n3014), .D(n1_adj_5416), .S(n57822));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1209 (.I0(n53171), .I1(n53063), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n60815));
    defparam i1_3_lut_adj_1209.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1210 (.I0(n53071), .I1(n25726), .I2(\data_in_frame[18] [3]), 
            .I3(GND_net), .O(n62170));
    defparam i1_3_lut_adj_1210.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1211 (.I0(n58383), .I1(n53772), .I2(\data_in_frame[18] [3]), 
            .I3(GND_net), .O(n62398));
    defparam i1_3_lut_adj_1211.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1212 (.I0(n62398), .I1(n62160), .I2(n62170), 
            .I3(n60815), .O(n58891));
    defparam i1_4_lut_adj_1212.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_in_frame[20][1] ), .I1(n24742), 
            .I2(GND_net), .I3(GND_net), .O(n58514));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58768));
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i49265_2_lut (.I0(\byte_transmit_counter[0] ), .I1(\data_out_frame[0][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65539));
    defparam i49265_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 data_in_frame_14__7__I_0_4037_2_lut (.I0(\data_in_frame[14] [7]), 
            .I1(\data_in_frame[14] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_654));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_14__7__I_0_4037_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[15] [4]), 
            .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29432));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i45860_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62876));
    defparam i45860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45861_4_lut (.I0(n62876), .I1(n65539), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n62877));
    defparam i45861_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i1_4_lut_adj_1216 (.I0(Kp_23__N_654), .I1(n58768), .I2(\data_in_frame[15] [1]), 
            .I3(\data_in_frame[17] [2]), .O(n62404));
    defparam i1_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i45859_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62875));
    defparam i45859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1217 (.I0(n25604), .I1(n58668), .I2(n58885), 
            .I3(n62404), .O(n62410));
    defparam i1_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1218 (.I0(n53102), .I1(n58913), .I2(n54173), 
            .I3(n62410), .O(n58394));
    defparam i1_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n3014), .D(n1_adj_5418), .S(n57827));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_in_frame[17] [1]), .I1(n58394), 
            .I2(GND_net), .I3(GND_net), .O(n53879));
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(n23529), .I1(\data_in_frame[21] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58427));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n62456));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1222 (.I0(n53463), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[11] [5]), .I3(GND_net), .O(n58879));
    defparam i1_2_lut_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1223 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n58465));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1224 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n58870));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1224.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29429));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1225 (.I0(n58885), .I1(n58787), .I2(n58671), 
            .I3(n62456), .O(n54184));
    defparam i1_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1226 (.I0(\data_in_frame[10] [5]), .I1(n4), 
            .I2(n25426), .I3(GND_net), .O(n58885));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1226.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1227 (.I0(n54284), .I1(n54184), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n53171));
    defparam i1_3_lut_adj_1227.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_adj_1228 (.I0(\data_in_frame[15] [3]), .I1(n58574), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n59916));
    defparam i1_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1229 (.I0(\data_in_frame[15] [5]), .I1(n54148), 
            .I2(n54284), .I3(GND_net), .O(n25343));
    defparam i2_3_lut_adj_1229.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1230 (.I0(\data_in_frame[10] [5]), .I1(n4), 
            .I2(n25511), .I3(\data_in_frame[12] [4]), .O(n25437));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [2]), .I3(\data_in_frame[18] [4]), .O(n58780));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1231 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[15] [3]), 
            .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1231.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1232 (.I0(n58588), .I1(n59932), .I2(n58822), 
            .I3(n25544), .O(n58913));
    defparam i1_4_lut_adj_1232.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1233 (.I0(n25604), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58946));
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h6666;
    SB_LUT4 equal_1927_i7_2_lut (.I0(Kp_23__N_974), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5388));   // verilog/coms.v(239[9:81])
    defparam equal_1927_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5420));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1234 (.I0(n25363), .I1(Kp_23__N_669), .I2(\data_in_frame[10] [7]), 
            .I3(GND_net), .O(n62448));
    defparam i1_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1235 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[19] [0]), .I3(GND_net), .O(n58303));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1236 (.I0(n58946), .I1(n53187), .I2(n60197), 
            .I3(n62448), .O(n58574));
    defparam i1_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1237 (.I0(n58816), .I1(n58574), .I2(n25525), 
            .I3(\data_in_frame[13] [5]), .O(n62220));
    defparam i1_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1238 (.I0(n62220), .I1(n54148), .I2(n58913), 
            .I3(\data_in_frame[17] [3]), .O(n53903));
    defparam i1_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5421));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(n25343), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58711));
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_LUT4 add_1083_9_lut (.I0(n57819), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n51254), .O(n57827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(Kp_23__N_1551), .I1(n53903), .I2(GND_net), 
            .I3(GND_net), .O(n54154));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_in_frame[16]_c [1]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58910));
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(n26055), .I1(n53703), .I2(GND_net), 
            .I3(GND_net), .O(n54173));
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25538));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5423), .S(n57969));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1244 (.I0(n25511), .I1(n25859), .I2(n25426), 
            .I3(GND_net), .O(n58459));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1245 (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[22] [6]), .I3(n58472), .O(n60682));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1246 (.I0(\data_in_frame[10] [7]), .I1(n62150), 
            .I2(\data_in_frame[11] [1]), .I3(n53374), .O(n58194));
    defparam i1_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1247 (.I0(\data_in_frame[1] [1]), .I1(n58337), 
            .I2(\data_in_frame[3][2] ), .I3(\data_in_frame[5] [4]), .O(n58534));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n62222));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1249 (.I0(n58346), .I1(n53096), .I2(n25538), 
            .I3(n62222), .O(n53102));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n62360));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1251 (.I0(n58588), .I1(n53102), .I2(n25596), 
            .I3(n62360), .O(n59932));
    defparam i1_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[13] [1]), .I1(n53187), 
            .I2(GND_net), .I3(GND_net), .O(n58787));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 add_1083_8_lut (.I0(n57819), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n51253), .O(n57822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1083_8 (.CI(n51253), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n51254));
    SB_LUT4 data_in_frame_12__7__I_0_4035_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_669));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_12__7__I_0_4035_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58798));
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5424));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25363));
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(n58825), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[12] [1]), .O(n62182));
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 add_1083_7_lut (.I0(n57819), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n51252), .O(n57821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1256 (.I0(n62182), .I1(n58798), .I2(Kp_23__N_669), 
            .I3(n58851), .O(n62188));
    defparam i1_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1257 (.I0(n25437), .I1(n62188), .I2(n58870), 
            .I3(GND_net), .O(n62192));
    defparam i1_3_lut_adj_1257.LUT_INIT = 16'h9696;
    SB_CARRY add_1083_7 (.CI(n51252), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n51253));
    SB_DFFE data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29426));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1258 (.I0(n53463), .I1(n58424), .I2(n58388), 
            .I3(n62192), .O(n62198));
    defparam i1_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1259 (.I0(n58958), .I1(n62198), .I2(n58551), 
            .I3(n58931), .O(n62204));
    defparam i1_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1260 (.I0(n53374), .I1(n58194), .I2(n54173), 
            .I3(n62204), .O(n53096));
    defparam i1_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1261 (.I0(n53096), .I1(n25363), .I2(\data_in_frame[15] [7]), 
            .I3(n25596), .O(n60751));
    defparam i3_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5425), .S(n57968));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1083_6_lut (.I0(n57819), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n51251), .O(n57826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_6_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29423));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1083_6 (.CI(n51251), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n51252));
    SB_LUT4 i1_4_lut_adj_1262 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [6]), 
            .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5426));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1262.LUT_INIT = 16'ha088;
    SB_LUT4 select_776_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5427));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_adj_1263 (.I0(\data_in_frame[16]_c [0]), .I1(n58787), 
            .I2(n59932), .I3(n60751), .O(n58897));
    defparam i2_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1264 (.I0(n58701), .I1(n58870), .I2(\data_in_frame[8] [7]), 
            .I3(n25503), .O(n10_adj_5428));
    defparam i4_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1265 (.I0(Kp_23__N_878), .I1(n10_adj_5428), .I2(n58620), 
            .I3(GND_net), .O(n25525));
    defparam i5_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1266 (.I0(Kp_23__N_993), .I1(n25525), .I2(n25859), 
            .I3(GND_net), .O(n58813));
    defparam i2_3_lut_adj_1266.LUT_INIT = 16'h9696;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(\FRAME_MATCHER.i [12]), .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5429), .S(n57967));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1267 (.I0(\data_in_frame[9] [4]), .I1(n58346), 
            .I2(n58571), .I3(n58813), .O(n60574));
    defparam i3_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1268 (.I0(n58910), .I1(\data_in_frame[16] [2]), 
            .I2(n60574), .I3(\data_in_frame[9] [3]), .O(n24742));
    defparam i3_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [20]), .I3(\FRAME_MATCHER.i [27]), .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_in_frame[18] [3]), .I1(n24742), 
            .I2(GND_net), .I3(GND_net), .O(n53067));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1270 (.I0(\data_in_frame[15] [5]), .I1(n58897), 
            .I2(\data_in_frame[13] [7]), .I3(\data_in_frame[17]_c [7]), 
            .O(n24730));
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [26]), .O(n41));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1271 (.I0(n58565), .I1(n58955), .I2(\data_in_frame[14] [1]), 
            .I3(GND_net), .O(n58934));
    defparam i2_3_lut_adj_1271.LUT_INIT = 16'h6969;
    SB_LUT4 select_776_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5430));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [18]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n25154));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23341_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25154), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i23341_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 select_776_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i472_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2209));   // verilog/coms.v(148[4] 304[11])
    defparam i472_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1272 (.I0(n58571), .I1(\data_in_frame[13] [7]), 
            .I2(n58810), .I3(n6_adj_5433), .O(n58854));
    defparam i4_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(n25757), .I1(n25944), .I2(\data_in_frame[16][5] ), 
            .I3(GND_net), .O(n53071));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[20]_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58717));
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1275 (.I0(n53071), .I1(n54274), .I2(n58383), 
            .I3(n6_adj_5434), .O(n53135));
    defparam i4_4_lut_adj_1275.LUT_INIT = 16'h9669;
    SB_LUT4 select_776_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51348_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[2]_c [7]), 
            .I2(n7), .I3(GND_net), .O(n57446));   // verilog/coms.v(94[13:20])
    defparam i51348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1271));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n24758), .I1(\data_in_frame[14] [0]), 
            .I2(n25544), .I3(Kp_23__N_1271), .O(n10_adj_5306));
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58324));
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29420));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29417));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29414));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51926 (.I0(byte_transmit_counter[1]), 
            .I1(n11_adj_5441), .I2(n12_adj_5442), .I3(byte_transmit_counter[2]), 
            .O(n68858));
    defparam byte_transmit_counter_1__bdd_4_lut_51926.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5443), .S(n57966));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29411));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1278 (.I0(n53772), .I1(\data_in_frame[20] [4]), 
            .I2(\data_in_frame[20][5] ), .I3(GND_net), .O(n58472));
    defparam i2_3_lut_adj_1278.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(\data_in_frame[16] [6]), .I1(n53130), 
            .I2(GND_net), .I3(GND_net), .O(n58158));
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58825));
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1281 (.I0(\data_in_frame[11] [7]), .I1(n53398), 
            .I2(GND_net), .I3(GND_net), .O(n58958));
    defparam i1_2_lut_adj_1281.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1282 (.I0(n58695), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[8] [0]), .I3(n6_adj_5447), .O(n60436));
    defparam i4_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29408));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1283 (.I0(n60436), .I1(\data_in_frame[6] [3]), 
            .I2(n58248), .I3(n58285), .O(n12_adj_5448));
    defparam i5_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 add_1083_5_lut (.I0(n57819), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n51250), .O(n57824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut (.I0(\data_in_frame[8] [3]), .I1(n12_adj_5448), .I2(\data_in_frame[12] [0]), 
            .I3(\data_in_frame[8] [4]), .O(n58955));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n58228), .I1(\data_in_frame[9] [5]), .I2(\data_in_frame[11] [6]), 
            .I3(n53862), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_1083_5 (.CI(n51250), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n51251));
    SB_DFFE data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29405));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1083_4_lut (.I0(n57819), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n51249), .O(n57825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10_4_lut (.I0(n58955), .I1(n58173), .I2(n58409), .I3(\data_in_frame[9] [0]), 
            .O(n26_c));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(n58958), .I1(n58542), .I2(n58928), .I3(n58340), 
            .O(n27_c));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1284 (.I0(\data_in_frame[5][3] ), .I1(n58876), 
            .I2(n58270), .I3(\data_in_frame[7] [1]), .O(n25));
    defparam i9_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_CARRY add_1083_4 (.CI(n51249), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n51250));
    SB_LUT4 i15_4_lut_adj_1285 (.I0(n25), .I1(n27_c), .I2(n26_c), .I3(n28), 
            .O(n24758));
    defparam i15_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 n68858_bdd_4_lut (.I0(n68858), .I1(n9), .I2(n65440), .I3(byte_transmit_counter[2]), 
            .O(n68861));
    defparam n68858_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51797 (.I0(byte_transmit_counter[1]), 
            .I1(n11_adj_5450), .I2(n12_adj_5451), .I3(byte_transmit_counter[2]), 
            .O(n68852));
    defparam byte_transmit_counter_1__bdd_4_lut_51797.LUT_INIT = 16'he4aa;
    SB_LUT4 n68852_bdd_4_lut (.I0(n68852), .I1(n9_adj_5452), .I2(n65441), 
            .I3(byte_transmit_counter[2]), .O(n68855));
    defparam n68852_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n69037), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 add_1083_3_lut (.I0(n57819), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n51248), .O(n57823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1083_3 (.CI(n51248), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n51249));
    SB_LUT4 i3_4_lut_adj_1286 (.I0(n58552), .I1(n58656), .I2(\data_in_frame[12] [2]), 
            .I3(n54203), .O(n25757));
    defparam i3_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n26617), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2189), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2190), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 add_1083_2_lut (.I0(n57819), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n57820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1083_2_lut.LUT_INIT = 16'h8228;
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20741), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n57202), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_in_frame[14] [2]), .I1(n24758), 
            .I2(GND_net), .I3(GND_net), .O(n26158));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2201), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n27160), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 select_776_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29402));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5454), .S(n57965));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1083_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3416), .CO(n51248));
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_in_frame[16][4] ), .I1(n58349), 
            .I2(GND_net), .I3(GND_net), .O(n25729));
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1289 (.I0(\data_in_frame[10] [3]), .I1(n58695), 
            .I2(n58455), .I3(n58267), .O(n26055));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51347_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[2]_c [6]), 
            .I2(n7), .I3(GND_net), .O(n57444));   // verilog/coms.v(94[13:20])
    defparam i51347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(n53770), .I1(Kp_23__N_1080), .I2(GND_net), 
            .I3(GND_net), .O(n58542));
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51792 (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5457), .I2(n5), .I3(byte_transmit_counter[2]), 
            .O(n68846));
    defparam byte_transmit_counter_1__bdd_4_lut_51792.LUT_INIT = 16'he4aa;
    SB_LUT4 select_776_Select_223_i3_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n58539), .I3(\data_out_frame[25] [6]), 
            .O(n3_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_776_Select_222_i3_4_lut (.I0(n53179), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5458), .I3(n60509), .O(n3_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_776_Select_221_i3_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n58433), .I3(\data_out_frame[25] [4]), 
            .O(n3_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_221_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i8_4_lut (.I0(n58906), .I1(n58484), .I2(n54307), .I3(\data_out_frame[25] [3]), 
            .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1291 (.I0(n58900), .I1(n58421), .I2(n58665), 
            .I3(n26424), .O(n24));
    defparam i10_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1292 (.I0(n58804), .I1(\data_out_frame[23] [0]), 
            .I2(n58254), .I3(n58943), .O(n23_c));
    defparam i9_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(\data_out_frame[20] [5]), .I1(n22), .I2(\data_out_frame[25] [2]), 
            .I3(GND_net), .O(n25_adj_5459));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_220_i3_4_lut (.I0(n25_adj_5459), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n23_c), .I3(n24), .O(n3_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(Kp_23__N_993), .I1(n53463), .I2(GND_net), 
            .I3(GND_net), .O(n54144));
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5297));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5296));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_776_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5295));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_776_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5294));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1294 (.I0(n25462), .I1(n53274), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n54138));
    defparam i1_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[21] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_219_i3_3_lut (.I0(n53925), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58499), .I3(GND_net), .O(n3_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_219_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 select_776_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_33_lut  (.I0(n65372), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n52061), .O(n27700)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_32_lut  (.I0(n65373), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n52060), .O(n27698)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1295 (.I0(n58864), .I1(n54138), .I2(n54144), 
            .I3(n62314), .O(n58724));
    defparam i1_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1296 (.I0(\data_in_frame[9] [0]), .I1(n25511), 
            .I2(n25859), .I3(GND_net), .O(n58388));
    defparam i2_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i51343_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[2]_c [4]), 
            .I2(n7), .I3(GND_net), .O(n57424));   // verilog/coms.v(94[13:20])
    defparam i51343_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_32  (.CI(n52060), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n52061));
    SB_LUT4 select_776_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5461));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_in_frame[14] [3]), .I1(n58248), 
            .I2(GND_net), .I3(GND_net), .O(n58656));
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1298 (.I0(\data_in_frame[14] [5]), .I1(n26055), 
            .I2(n58400), .I3(\data_in_frame[12] [4]), .O(n53130));
    defparam i3_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_31_lut  (.I0(n65374), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n52059), .O(n27696)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_776_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(n25604), .I1(\data_in_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58424));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i51346_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[2]_c [2]), 
            .I2(n7), .I3(GND_net), .O(n57442));   // verilog/coms.v(94[13:20])
    defparam i51346_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29399));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_31  (.CI(n52059), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n52060));
    SB_LUT4 select_776_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5463));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(n25549), .I1(n25569), .I2(GND_net), 
            .I3(GND_net), .O(n26043));
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1301 (.I0(n54138), .I1(n58534), .I2(\data_in_frame[10] [2]), 
            .I3(\data_in_frame[7] [6]), .O(n12_adj_5464));
    defparam i5_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(\data_in_frame[7] [7]), .I1(n12_adj_5464), 
            .I2(n58565), .I3(n25923), .O(n53703));
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1303 (.I0(n53703), .I1(\data_in_frame[14] [4]), 
            .I2(n53398), .I3(GND_net), .O(n58599));
    defparam i2_3_lut_adj_1303.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1304 (.I0(\data_in_frame[17][0] ), .I1(n54180), 
            .I2(\data_in_frame[14] [6]), .I3(GND_net), .O(n58531));
    defparam i2_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5465));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_30_lut  (.I0(n65379), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n52058), .O(n27694)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_30  (.CI(n52058), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n52059));
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n29398), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1305 (.I0(n58531), .I1(n58599), .I2(\data_in_frame[16][5] ), 
            .I3(n58291), .O(n12_adj_5466));
    defparam i5_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29395));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1306 (.I0(n53130), .I1(n12_adj_5466), .I2(n58656), 
            .I3(n54203), .O(n60010));
    defparam i6_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_29_lut  (.I0(n65382), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n52057), .O(n27692)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5467), .S(n57964));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_29  (.CI(n52057), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n52058));
    SB_LUT4 i1_2_lut_adj_1307 (.I0(n60010), .I1(\data_in_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58596));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h9999;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_28_lut  (.I0(n65386), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n52056), .O(n27690)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_776_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_28  (.CI(n52056), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n52057));
    SB_DFFE data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29392));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_27_lut  (.I0(n65387), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n52055), .O(n27688)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_in_frame[1] [5]), .I1(n58182), 
            .I2(GND_net), .I3(GND_net), .O(n25441));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_27  (.CI(n52055), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n52056));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_26_lut  (.I0(n65393), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n52054), .O(n27686)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i3_4_lut_adj_1309 (.I0(\data_in_frame[8] [0]), .I1(n58391), 
            .I2(n25963), .I3(n25441), .O(n25462));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_26  (.CI(n52054), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n52055));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_25_lut  (.I0(n65394), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n52053), .O(n27684)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_25  (.CI(n52053), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n52054));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_24_lut  (.I0(n65395), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n52052), .O(n27682)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_24  (.CI(n52052), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n52053));
    SB_LUT4 i3_4_lut_adj_1310 (.I0(n53770), .I1(n26388), .I2(n25462), 
            .I3(\data_in_frame[10] [1]), .O(n58551));
    defparam i3_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_23_lut  (.I0(n65398), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n52051), .O(n27680)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[9] [7]), .I1(n58551), 
            .I2(GND_net), .I3(GND_net), .O(n58552));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_23  (.CI(n52051), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n52052));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_22_lut  (.I0(n65399), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n52050), .O(n27678)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_22  (.CI(n52050), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n52051));
    SB_DFFE data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29389));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29386));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22376_4_lut (.I0(n27924), .I1(n65543), .I2(rx_data[5]), .I3(\data_in_frame[23] [5]), 
            .O(n38036));   // verilog/coms.v(94[13:20])
    defparam i22376_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_21_lut  (.I0(n65400), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n52049), .O(n27676)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_21  (.CI(n52049), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n52050));
    SB_LUT4 i2_3_lut_adj_1312 (.I0(n25437), .I1(\data_in_frame[15] [0]), 
            .I2(\data_in_frame[12] [6]), .I3(GND_net), .O(n58668));
    defparam i2_3_lut_adj_1312.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1313 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [5]), 
            .I2(n58291), .I3(n6_adj_5470), .O(n24756));
    defparam i4_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i22377_3_lut (.I0(n38036), .I1(\data_in_frame[23] [5]), .I2(reset), 
            .I3(GND_net), .O(n29864));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1314 (.I0(n25944), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[17] [1]), .I3(n58531), .O(n10_adj_5471));
    defparam i4_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_20_lut  (.I0(n65401), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n52048), .O(n27674)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_20  (.CI(n52048), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n52049));
    SB_LUT4 select_776_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_adj_1315 (.I0(\data_in_frame[16][7] ), .I1(n10_adj_5471), 
            .I2(\data_in_frame[19] [2]), .I3(GND_net), .O(n58520));
    defparam i5_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[23] [4]), .I1(n27924), .I2(n28009), 
            .I3(rx_data[4]), .O(n57300));   // verilog/coms.v(94[13:20])
    defparam i13_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_19_lut  (.I0(n65428), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n52047), .O(n27672)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_19  (.CI(n52047), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n52048));
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_in_frame[21] [2]), .I1(n54274), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5473));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_18_lut  (.I0(n65451), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n52046), .O(n27670)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_18  (.CI(n52046), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n52047));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_17_lut  (.I0(n65465), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n52045), .O(n27668)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13_4_lut_adj_1317 (.I0(\data_in_frame[23] [3]), .I1(n27924), 
            .I2(n28009), .I3(rx_data[3]), .O(n57302));   // verilog/coms.v(94[13:20])
    defparam i13_4_lut_adj_1317.LUT_INIT = 16'h3a0a;
    SB_LUT4 i4_4_lut_adj_1318 (.I0(n25729), .I1(n54156), .I2(n58303), 
            .I3(n6_adj_5473), .O(n58801));
    defparam i4_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5474));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_17  (.CI(n52045), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n52046));
    SB_DFFE data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29383));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_16_lut  (.I0(n65476), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n52044), .O(n27666)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i3_4_lut_adj_1319 (.I0(\data_in_frame[21]_c [3]), .I1(n54156), 
            .I2(n58520), .I3(n24756), .O(n58554));
    defparam i3_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_16  (.CI(n52044), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n52045));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_15_lut  (.I0(n65479), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n52043), .O(n27664)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(n58270), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5476));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1321 (.I0(n25370), .I1(n7_adj_5476), .I2(n26225), 
            .I3(n8_adj_5477), .O(n53463));
    defparam i5_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29380));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_15  (.CI(n52043), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n52044));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_14_lut  (.I0(n65480), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n52042), .O(n27662)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_14  (.CI(n52042), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n52043));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_13_lut  (.I0(n65481), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n52041), .O(n27660)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 n68846_bdd_4_lut (.I0(n68846), .I1(n65442), .I2(n1_adj_5478), 
            .I3(byte_transmit_counter[2]), .O(n68849));
    defparam n68846_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_776_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5479));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_13  (.CI(n52041), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n52042));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_12_lut  (.I0(n65482), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n52040), .O(n27658)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_12  (.CI(n52040), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n52041));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_11_lut  (.I0(n65487), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n52039), .O(n27656)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(n38022), .I1(n39291), .I2(GND_net), 
            .I3(GND_net), .O(n27924));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'hbbbb;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_11  (.CI(n52039), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n52040));
    SB_DFFE data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29377));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51787 (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5480), .I2(n5_adj_5481), .I3(byte_transmit_counter[2]), 
            .O(n68840));
    defparam byte_transmit_counter_1__bdd_4_lut_51787.LUT_INIT = 16'he4aa;
    SB_LUT4 n68840_bdd_4_lut (.I0(n68840), .I1(n65444), .I2(n65443), .I3(byte_transmit_counter[2]), 
            .O(n68843));
    defparam n68840_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51881 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n68828));
    defparam byte_transmit_counter_0__bdd_4_lut_51881.LUT_INIT = 16'he4aa;
    SB_LUT4 n68828_bdd_4_lut (.I0(n68828), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n68831));
    defparam n68828_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51772 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n68822));
    defparam byte_transmit_counter_0__bdd_4_lut_51772.LUT_INIT = 16'he4aa;
    SB_LUT4 select_776_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5482));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n68822_bdd_4_lut (.I0(n68822), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n68825));
    defparam n68822_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_10_lut  (.I0(n65489), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n52038), .O(n27654)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_10  (.CI(n52038), .I0(n27913), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n52039));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_9_lut  (.I0(n65491), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n52037), .O(n27652)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_9  (.CI(n52037), .I0(n27913), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n52038));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_8_lut  (.I0(n65495), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n52036), .O(n27650)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_776_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5484));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_8  (.CI(n52036), .I0(n27913), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n52037));
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58200));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51767 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n68816));
    defparam byte_transmit_counter_0__bdd_4_lut_51767.LUT_INIT = 16'he4aa;
    SB_LUT4 select_776_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_adj_1324 (.I0(n34), .I1(n54235), .I2(n58582), .I3(GND_net), 
            .O(n8_adj_5486));
    defparam i3_3_lut_adj_1324.LUT_INIT = 16'h6969;
    SB_LUT4 select_776_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5486), .I3(\data_out_frame[25] [0]), 
            .O(n3_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_7_lut  (.I0(n65499), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n52035), .O(n27648)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_7  (.CI(n52035), .I0(n27913), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n52036));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_6_lut  (.I0(n65500), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n52034), .O(n27646)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1325 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58671));
    defparam i1_2_lut_adj_1325.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_6  (.CI(n52034), .I0(n27913), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n52035));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_5_lut  (.I0(n65501), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n52033), .O(n27644)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_776_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5487));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1326 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58851));
    defparam i1_2_lut_adj_1326.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17]_c [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_5  (.CI(n52033), .I0(n27913), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n52034));
    SB_DFFE data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29374));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[20] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1327 (.I0(n58294), .I1(n58671), .I2(\data_in_frame[10] [7]), 
            .I3(n25511), .O(n12_adj_5488));
    defparam i5_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1328 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[13] [3]), 
            .I2(n12_adj_5488), .I3(n8_adj_5489), .O(n54284));
    defparam i1_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_4_lut  (.I0(n65503), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n52032), .O(n27642)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_4  (.CI(n52032), .I0(n27913), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n52033));
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_3_lut  (.I0(n65506), .I1(n27913), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n52031), .O(n27640)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 select_776_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_3  (.CI(n52031), .I0(n27913), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n52032));
    SB_LUT4 i2_4_lut_adj_1329 (.I0(n54284), .I1(Kp_23__N_1389), .I2(n6_adj_5492), 
            .I3(n58297), .O(n58765));
    defparam i2_4_lut_adj_1329.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1330 (.I0(n58692), .I1(n58327), .I2(n58928), 
            .I3(n26225), .O(n25549));
    defparam i1_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1934_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1934_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1331 (.I0(\data_in_frame[11] [6]), .I1(n25549), 
            .I2(GND_net), .I3(GND_net), .O(n58931));
    defparam i1_2_lut_adj_1331.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29371));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1332 (.I0(n58794), .I1(n58315), .I2(n54146), 
            .I3(n58207), .O(n10_adj_5493));
    defparam i4_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1333 (.I0(\data_out_frame[18] [7]), .I1(n58527), 
            .I2(n68374), .I3(\data_out_frame[19] [1]), .O(n58900));
    defparam i3_4_lut_adj_1333.LUT_INIT = 16'h9669;
    SB_CARRY \FRAME_MATCHER.i_1934_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n52031));
    SB_LUT4 i6_4_lut_adj_1334 (.I0(n58961), .I1(n58207), .I2(n58900), 
            .I3(n43_adj_5494), .O(n14_adj_5495));
    defparam i6_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5496));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25280));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_in_frame[6] [5]), .I1(Kp_23__N_875), 
            .I2(GND_net), .I3(GND_net), .O(n58228));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1337 (.I0(n25645), .I1(n58937), .I2(n58791), 
            .I3(n25845), .O(n13_adj_5497));
    defparam i5_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i51364_4_lut (.I0(n53247), .I1(n13_adj_5497), .I2(n25845), 
            .I3(n14_adj_5495), .O(n68380));
    defparam i51364_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29368));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1338 (.I0(\data_out_frame[22] [7]), .I1(n58212), 
            .I2(\data_out_frame[16] [1]), .I3(n68380), .O(n58665));
    defparam i3_4_lut_adj_1338.LUT_INIT = 16'h9669;
    SB_LUT4 select_776_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29365));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1339 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[10] [1]), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1339.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29362));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29359));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1340 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58294));
    defparam i1_2_lut_adj_1340.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1341 (.I0(n25871), .I1(\data_in_frame[8] [6]), 
            .I2(\data_in_frame[13] [5]), .I3(\data_in_frame[13] [4]), .O(n10_adj_5501));   // verilog/coms.v(88[17:63])
    defparam i4_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1342 (.I0(\data_in_frame[15] [6]), .I1(n10_adj_5501), 
            .I2(\data_in_frame[11] [2]), .I3(GND_net), .O(n58882));   // verilog/coms.v(88[17:63])
    defparam i5_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58212));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5503), .S(n57963));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1344 (.I0(n60532), .I1(\data_out_frame[23] [3]), 
            .I2(n58212), .I3(n6_adj_5504), .O(n60509));
    defparam i4_4_lut_adj_1344.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29356));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1345 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[23] [1]), 
            .I2(n58665), .I3(n58848), .O(n15));
    defparam i6_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29353));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29350));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5507));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n68816_bdd_4_lut (.I0(n68816), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n68819));
    defparam n68816_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29347));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i8_4_lut_adj_1346 (.I0(n15), .I1(n58288), .I2(n14_adj_5508), 
            .I3(\data_out_frame[21] [1]), .O(n58433));
    defparam i8_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29344));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29341));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5509));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29338));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29335));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1347 (.I0(\data_out_frame[16] [4]), .I1(n53247), 
            .I2(GND_net), .I3(GND_net), .O(n58421));
    defparam i1_2_lut_adj_1347.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29332));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1348 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [2]), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1348.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29329));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29326));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29323));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29320));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29317));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29314));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29311));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1349 (.I0(n11_adj_5512), .I1(n54197), .I2(n58380), 
            .I3(GND_net), .O(n53925));
    defparam i6_4_lut_adj_1349.LUT_INIT = 16'h6969;
    SB_LUT4 select_776_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27308), 
            .D(n4793[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29308));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29305));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29302));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29299));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5515));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29296));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29293));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29290));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29287));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29284));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29281));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5516));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5517), .S(n57832));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29278));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_217_i3_4_lut (.I0(n54150), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5518), .I3(n58433), .O(n3_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_217_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29275));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1350 (.I0(n8_adj_5519), .I1(n38022), .I2(GND_net), 
            .I3(GND_net), .O(n27926));
    defparam i1_2_lut_adj_1350.LUT_INIT = 16'heeee;
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29272));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29269));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29266));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29263));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29260));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3]_c [7]), .C(clk16MHz), 
           .D(n29087));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5521));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_776_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n57510));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n57494));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n29107));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n29110));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n29113));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n57504));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n29165));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n29184));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5][0] ), .C(clk16MHz), 
           .D(n29188));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n29191));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5][2] ), .C(clk16MHz), 
           .D(n29194));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1351 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [2]), 
            .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5284));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1351.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51762 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[1]), .O(n68810));
    defparam byte_transmit_counter_0__bdd_4_lut_51762.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5][3] ), .C(clk16MHz), 
           .D(n29206));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n29209));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n68810_bdd_4_lut (.I0(n68810), .I1(\data_out_frame[21] [0]), 
            .I2(\data_out_frame[20] [0]), .I3(byte_transmit_counter[1]), 
            .O(n68813));
    defparam n68810_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_776_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51757 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(byte_transmit_counter[1]), .O(n68804));
    defparam byte_transmit_counter_0__bdd_4_lut_51757.LUT_INIT = 16'he4aa;
    SB_LUT4 n68804_bdd_4_lut (.I0(n68804), .I1(\data_out_frame[21] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(byte_transmit_counter[1]), 
            .O(n68807));
    defparam n68804_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51752 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(byte_transmit_counter[1]), .O(n68798));
    defparam byte_transmit_counter_0__bdd_4_lut_51752.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5]_c [5]), .C(clk16MHz), 
           .D(n29212));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5][6] ), .C(clk16MHz), 
           .D(n57514));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5]_c [7]), .C(clk16MHz), 
           .D(n57520));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27308), 
            .D(n4793[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27308), 
            .D(n4793[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27308), 
            .D(n4793[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27308), 
            .D(n4793[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n29221));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29231));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n68798_bdd_4_lut (.I0(n68798), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(byte_transmit_counter[1]), 
            .O(n68801));
    defparam n68798_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27308), 
            .D(n4793[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27308), 
            .D(n4793[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27308), 
            .D(n4793[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27308), 
            .D(n4793[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27308), 
            .D(n4793[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27308), 
            .D(n4793[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27308), 
            .D(n4793[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27308), 
            .D(n4793[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27308), 
            .D(n4793[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27308), 
            .D(n4793[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27308), 
            .D(n4793[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27308), 
            .D(n4793[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27308), 
            .D(n4793[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27308), 
            .D(n4793[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27308), 
            .D(n4793[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27308), 
            .D(n4793[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27308), 
            .D(n4793[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27308), 
            .D(n4793[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n29224));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29227));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5524), .S(n57962));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n39291), 
            .I2(reset), .I3(n62), .O(n28009));
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h0400;
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8][3] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5525), .S(n57961));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8][4] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5526), .S(n57960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8][5] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5527), .S(n57959));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8][6] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5528), .S(n57958));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11852_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27592));   // verilog/coms.v(109[34:55])
    defparam i11852_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8][7] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5529), .S(n57957));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i45857_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62873));
    defparam i45857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_2_lut_adj_1352 (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut_adj_1352.LUT_INIT = 16'h2222;
    SB_LUT4 i45858_4_lut (.I0(n62873), .I1(n27592), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n62874));
    defparam i45858_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51737 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n68780));
    defparam byte_transmit_counter_0__bdd_4_lut_51737.LUT_INIT = 16'he4aa;
    SB_LUT4 i45856_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62872));
    defparam i45856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n68780_bdd_4_lut (.I0(n68780), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n68783));
    defparam n68780_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1353 (.I0(n3579), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(reset), .O(n58121));
    defparam i1_2_lut_3_lut_4_lut_adj_1353.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1354 (.I0(n3579), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_5530), 
            .O(n58133));
    defparam i1_2_lut_3_lut_4_lut_adj_1354.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1355 (.I0(n3579), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_5531), 
            .O(n58118));
    defparam i1_2_lut_3_lut_4_lut_adj_1355.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1356 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2]_c [7]), 
            .I2(n25448), .I3(\data_in_frame[5][3] ), .O(n58327));
    defparam i1_2_lut_3_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1357 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [1]), 
            .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5283));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1357.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51732 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n68750));
    defparam byte_transmit_counter_0__bdd_4_lut_51732.LUT_INIT = 16'he4aa;
    SB_LUT4 select_776_Select_71_i2_4_lut (.I0(\data_out_frame[8][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_70_i2_4_lut (.I0(\data_out_frame[8][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_69_i2_4_lut (.I0(\data_out_frame[8][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5527));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_68_i2_4_lut (.I0(\data_out_frame[8][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n53055), .I1(n60075), .I2(\data_out_frame[20] [4]), 
            .I3(n53790), .O(n6_adj_5532));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_776_Select_67_i2_4_lut (.I0(\data_out_frame[8][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1358 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(n53666), .I3(\data_out_frame[18] [3]), .O(n58478));
    defparam i1_2_lut_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5523), .S(n58003));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5522), .S(n58002));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5521), .S(n58001));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5520), .S(n58000));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5516), .S(n57999));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5515), .S(n57998));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5514), .S(n57997));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5513), .S(n57956));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5511), .S(n57955));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5510), .S(n26));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5509), .S(n57954));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5507), .S(n57953));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5506), .S(n57952));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5505), .S(n57951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5502), .S(n57950));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5500), .S(n57949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5499), .S(n57948));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5498), .S(n57947));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5496), .S(n57946));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5491), .S(n57945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5490), .S(n57944));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5487), .S(n57943));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5485), .S(n57942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5484), .S(n57941));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5483), .S(n57940));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5482), .S(n57939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5479), .S(n57938));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5475), .S(n57937));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5474), .S(n57936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5472), .S(n57935));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5469), .S(n57934));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5468), .S(n57933));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5465), .S(n57932));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5463), .S(n57931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5462), .S(n57930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5461), .S(n57929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5460), .S(n57928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5456), .S(n57927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5455), .S(n57926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5453), .S(n57925));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5449), .S(n57924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5446), .S(n57923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5445), .S(n57922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5444), .S(n57921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5440), .S(n57920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5439), .S(n57919));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5438), .S(n57918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5437), .S(n57917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5435), .S(n57916));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5432), .S(n57915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5431), .S(n57914));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5430), .S(n57913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5427), .S(n57912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5426), .S(n57911));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5424), .S(n57898));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5422), .S(n57910));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5421), .S(n57909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5420), .S(n57908));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5419), .S(n57897));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5417), .S(n28838));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5410), .S(n28837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5401), .S(n57907));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5399), .S(n57906));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5395), .S(n57904));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5392), .S(n57905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5389), .S(n57833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5385), .S(n28831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5320), .S(n57903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5316), .S(n57902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5315), .S(n57901));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5311), .S(n28827));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5307), .S(n57900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5298), .S(n28825));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5534), .S(n57899));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5535), .S(n57891));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n29086));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n68750_bdd_4_lut (.I0(n68750), .I1(\data_out_frame[21] [4]), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n68753));
    defparam n68750_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12797_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28540));   // verilog/coms.v(130[12] 305[6])
    defparam i12797_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i45614_3_lut_4_lut (.I0(n25370), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [0]), .I3(Kp_23__N_748), .O(n62621));
    defparam i45614_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1359 (.I0(Kp_23__N_974), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[9] [1]), .I3(n58934), .O(n58759));
    defparam i1_2_lut_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n29085));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n29084));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n29083));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n29082));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n29081));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n29080));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5536), .S(n57890));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n29079));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n29078));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51707 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n68744));
    defparam byte_transmit_counter_0__bdd_4_lut_51707.LUT_INIT = 16'he4aa;
    SB_LUT4 i12793_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n26862), .I3(n24_adj_5537), .O(n28536));   // verilog/coms.v(130[12] 305[6])
    defparam i12793_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n29077));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n68744_bdd_4_lut (.I0(n68744), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n68747));
    defparam n68744_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n29076));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n29075));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n29074));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n29073));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n29072));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n29071));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n29070));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n29069));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n29068));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1934__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n27612), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n29067));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n29066));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n29065));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n3014), .D(n1_adj_5538), .S(n28540));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n29064));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n29063));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n3014), .D(n5_adj_5539), 
            .S(n28536));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n29062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n29061));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n29060));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n29059));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n29058));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n29057));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n29056));   // verilog/coms.v(130[12] 305[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29052));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n11_adj_5540), .I2(n12_adj_5541), .I3(byte_transmit_counter[2]), 
            .O(n69014));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_3_lut_adj_1360 (.I0(\data_out_frame[22] [5]), .I1(n6_adj_5532), 
            .I2(\data_out_frame[22] [4]), .I3(GND_net), .O(n34));
    defparam i3_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1361 (.I0(n25544), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[9] [1]), .O(n6_adj_5492));
    defparam i2_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29041));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_776_Select_216_i3_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n58418), .I3(n34), .O(n3_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_216_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i2_2_lut_3_lut_3_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(reset), 
            .I3(GND_net), .O(n22362));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58499));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1363 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n58146), .O(n58147));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1363.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1364 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n38022), .O(n27920));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1364.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_1365 (.I0(\data_out_frame[21] [1]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58484));
    defparam i1_2_lut_adj_1365.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1366 (.I0(n58484), .I1(n53119), .I2(n60532), 
            .I3(n58736), .O(n10_adj_5542));
    defparam i4_4_lut_adj_1366.LUT_INIT = 16'h9669;
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n3014), .D(n26494), 
            .S(n28471));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1367 (.I0(\data_out_frame[16] [2]), .I1(n58961), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n58794));
    defparam i2_3_lut_adj_1367.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5543), .S(n57889));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1368 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[22] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58943));
    defparam i1_2_lut_adj_1368.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(n32799), .O(n6_adj_5544));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29019), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12728_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28471));   // verilog/coms.v(130[12] 305[6])
    defparam i12728_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4_4_lut_adj_1369 (.I0(n58903), .I1(n53169), .I2(n58940), 
            .I3(n6_adj_5545), .O(n58380));
    defparam i4_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(\data_out_frame[23] [0]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58582));
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[24] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58714));
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h6666;
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29018));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(clk16MHz), .E(n3014), .D(n1_adj_5546), .S(n57820));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29017));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29016));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17_4_lut_adj_1372 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[23] [5]), 
            .I2(\data_out_frame[24] [3]), .I3(n58916), .O(n42_adj_5547));
    defparam i17_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1373 (.I0(n58784), .I1(\data_out_frame[23] [2]), 
            .I2(n53283), .I3(n54293), .O(n40_adj_5548));
    defparam i15_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1374 (.I0(n58714), .I1(n54197), .I2(\data_out_frame[23] [6]), 
            .I3(\data_out_frame[24] [5]), .O(n41_adj_5549));
    defparam i16_4_lut_adj_1374.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut_adj_1375 (.I0(n58462), .I1(n58582), .I2(\data_out_frame[23] [3]), 
            .I3(n54278), .O(n39_adj_5550));
    defparam i14_4_lut_adj_1375.LUT_INIT = 16'h9669;
    SB_LUT4 i13_3_lut (.I0(\data_out_frame[20] [1]), .I1(n58689), .I2(\data_out_frame[24] [4]), 
            .I3(GND_net), .O(n38_c));
    defparam i13_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i18_4_lut_adj_1376 (.I0(n58380), .I1(n60272), .I2(n58778), 
            .I3(n58819), .O(n43_adj_5551));
    defparam i18_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n39_adj_5550), .I1(n41_adj_5549), .I2(n40_adj_5548), 
            .I3(n42_adj_5547), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29012), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22_4_lut (.I0(n43_adj_5551), .I1(\data_out_frame[21] [5]), 
            .I2(n38_c), .I3(n53191), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1377 (.I0(n47), .I1(n8_adj_5552), .I2(n58499), 
            .I3(n48), .O(n54150));
    defparam i4_4_lut_adj_1377.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1378 (.I0(n54150), .I1(\data_out_frame[25] [0]), 
            .I2(n25947), .I3(GND_net), .O(n58418));
    defparam i2_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1379 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n58118), .O(n27918));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1379.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1380 (.I0(n58197), .I1(n58626), .I2(\data_out_frame[7] [1]), 
            .I3(n25656), .O(n10));   // verilog/coms.v(74[16:62])
    defparam i2_2_lut_3_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1381 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[8][6] ), .O(n38));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i51353_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[5]_c [7]), 
            .I2(n27972), .I3(GND_net), .O(n57520));   // verilog/coms.v(94[13:20])
    defparam i51353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51352_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[5][6] ), .I2(n27972), 
            .I3(GND_net), .O(n57514));   // verilog/coms.v(94[13:20])
    defparam i51352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1382 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[5] [6]), .O(n58626));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1383 (.I0(\data_out_frame[24] [4]), .I1(n53790), 
            .I2(n58318), .I3(GND_net), .O(n58306));
    defparam i1_3_lut_adj_1383.LUT_INIT = 16'h6969;
    SB_LUT4 select_776_Select_213_i3_4_lut (.I0(n58306), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58397), .I3(\data_out_frame[24] [3]), .O(n3_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_213_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13469_3_lut (.I0(\data_in_frame[5]_c [5]), .I1(rx_data[5]), 
            .I2(n27972), .I3(GND_net), .O(n29212));   // verilog/coms.v(130[12] 305[6])
    defparam i13469_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1384 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(\data_out_frame[14] [4]), .I3(n58254), .O(n58511));
    defparam i2_2_lut_3_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_212_i3_4_lut (.I0(n58398), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\data_out_frame[24] [2]), .I3(\data_out_frame[24] [3]), 
            .O(n3_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_212_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_adj_1385 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58462));
    defparam i1_2_lut_adj_1385.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1386 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(\data_out_frame[14] [4]), .I3(n25814), .O(n58207));
    defparam i2_2_lut_3_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_211_i3_4_lut (.I0(n23340), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58462), .I3(n54259), .O(n3_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_211_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_4_lut_adj_1387 (.I0(\data_in_frame[3]_c [5]), .I1(n58162), 
            .I2(\data_in_frame[1] [5]), .I3(n58267), .O(n25497));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n58017));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 select_776_Select_210_i3_4_lut (.I0(n53283), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_6), .I3(\data_out_frame[24] [0]), .O(n3_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_210_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i2_3_lut_adj_1388 (.I0(n58370), .I1(n58561), .I2(n1699), .I3(GND_net), 
            .O(n58804));
    defparam i2_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1389 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n58016));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1389.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1390 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n58015));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1390.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1391 (.I0(n53055), .I1(n60075), .I2(GND_net), 
            .I3(GND_net), .O(n54307));
    defparam i1_2_lut_adj_1391.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1392 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n58018));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1392.LUT_INIT = 16'h5100;
    SB_LUT4 i3_4_lut_adj_1393 (.I0(\data_out_frame[20] [2]), .I1(n58774), 
            .I2(n58502), .I3(n26202), .O(n53790));
    defparam i3_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1394 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n58014));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1394.LUT_INIT = 16'h5100;
    SB_LUT4 i3_4_lut_adj_1395 (.I0(n53164), .I1(n58491), .I2(n25797), 
            .I3(n58707), .O(n58774));
    defparam i3_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1396 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n58009));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1396.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1397 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n58007));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1397.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1398 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n58021));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1398.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1399 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n58008));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1399.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1400 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n58011));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1400.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1401 (.I0(n54146), .I1(n53119), .I2(GND_net), 
            .I3(GND_net), .O(n58937));
    defparam i1_2_lut_adj_1401.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25797));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1403 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n58012));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1403.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58315));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1405 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[12] [1]), .I3(n6_adj_5556), .O(n1673));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1406 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n58019));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1406.LUT_INIT = 16'h5100;
    SB_LUT4 i6_4_lut_adj_1407 (.I0(n58475), .I1(n1673), .I2(n58653), .I3(n58629), 
            .O(n16));
    defparam i6_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1408 (.I0(n58166), .I1(n58635), .I2(n58683), 
            .I3(n58579), .O(n17));
    defparam i7_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1409 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n58013));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1409.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1410 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n58006));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1410.LUT_INIT = 16'h5100;
    SB_LUT4 i9_4_lut_adj_1411 (.I0(n17), .I1(n58231), .I2(n16), .I3(\data_out_frame[10] [7]), 
            .O(n60061));
    defparam i9_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1412 (.I0(n54182), .I1(n1513), .I2(n1673), .I3(GND_net), 
            .O(n14_adj_5557));
    defparam i5_3_lut_adj_1412.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1413 (.I0(n60061), .I1(\data_out_frame[14] [1]), 
            .I2(n24670), .I3(n25666), .O(n15_adj_5558));
    defparam i6_4_lut_adj_1413.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1414 (.I0(n15_adj_5558), .I1(n1510), .I2(n14_adj_5557), 
            .I3(\data_out_frame[13] [7]), .O(n53247));
    defparam i8_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1415 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26202));
    defparam i1_2_lut_adj_1415.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1416 (.I0(n53247), .I1(n58254), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n59852));
    defparam i2_3_lut_adj_1416.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1417 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [3]), 
            .I2(n58495), .I3(n25830), .O(n16_adj_5559));
    defparam i6_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1418 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n58010));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1418.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1419 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n58020));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1419.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1420 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n58118), .O(n27916));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1420.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1421 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25082), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n62488));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1421.LUT_INIT = 16'hfff4;
    SB_LUT4 i7_4_lut_adj_1422 (.I0(\data_out_frame[17] [4]), .I1(n26431), 
            .I2(n58733), .I3(\data_out_frame[17] [2]), .O(n17_adj_5560));
    defparam i7_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1423 (.I0(n58771), .I1(n25992), .I2(n58443), 
            .I3(\data_out_frame[14] [3]), .O(n14_adj_5561));   // verilog/coms.v(78[16:43])
    defparam i6_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1424 (.I0(n25797), .I1(n58647), .I2(n25814), 
            .I3(\data_out_frame[16] [5]), .O(n13_adj_5562));   // verilog/coms.v(78[16:43])
    defparam i5_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1425 (.I0(n17_adj_5560), .I1(n68374), .I2(n16_adj_5559), 
            .I3(\data_out_frame[17] [1]), .O(n60254));
    defparam i9_4_lut_adj_1425.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1426 (.I0(\data_out_frame[19] [4]), .I1(n58315), 
            .I2(n58848), .I3(\data_out_frame[14] [4]), .O(n22_adj_5563));
    defparam i9_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n54243), .I1(n26199), .I2(n2076), .I3(GND_net), 
            .O(n20_adj_5564));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1427 (.I0(n58937), .I1(n2107), .I2(n58686), .I3(n26288), 
            .O(n21_c));
    defparam i8_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1428 (.I0(n60254), .I1(\data_out_frame[19] [3]), 
            .I2(n13_adj_5562), .I3(n14_adj_5561), .O(n19_c));
    defparam i6_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1429 (.I0(n19_c), .I1(n21_c), .I2(n20_adj_5564), 
            .I3(n22_adj_5563), .O(n58602));
    defparam i12_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1430 (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[19] [5]), 
            .I2(n58602), .I3(n59852), .O(n58807));
    defparam i3_4_lut_adj_1430.LUT_INIT = 16'h9669;
    SB_LUT4 i45988_3_lut (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[9] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63004));
    defparam i45988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45989_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63005));
    defparam i45989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45986_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63002));
    defparam i45986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45985_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63001));
    defparam i45985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45829_3_lut (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62845));
    defparam i45829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45830_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62846));
    defparam i45830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45848_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62864));
    defparam i45848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n69014_bdd_4_lut (.I0(n69014), .I1(n9_adj_5565), .I2(n65490), 
            .I3(byte_transmit_counter[2]), .O(n62994));
    defparam n69014_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i45847_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62863));
    defparam i45847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45835_3_lut (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62851));
    defparam i45835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45836_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62852));
    defparam i45836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51697 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n68732));
    defparam byte_transmit_counter_0__bdd_4_lut_51697.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5566), .S(n57888));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i45821_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62837));
    defparam i45821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45820_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62836));
    defparam i45820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45841_3_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[9] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62857));
    defparam i45841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45842_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62858));
    defparam i45842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1431 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25800));
    defparam i1_2_lut_adj_1431.LUT_INIT = 16'h6666;
    SB_LUT4 i45797_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62813));
    defparam i45797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1432 (.I0(n2217), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [4]), .I3(GND_net), .O(n58791));
    defparam i2_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_LUT4 i45796_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62812));
    defparam i45796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45884_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62900));
    defparam i45884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45885_4_lut (.I0(n62900), .I1(n27707), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n62901));
    defparam i45885_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i45883_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62899));
    defparam i45883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48733_2_lut (.I0(n68693), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65478));
    defparam i48733_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n29486));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50511_3_lut (.I0(n68831), .I1(n68813), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67527));
    defparam i50511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11860_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27600));   // verilog/coms.v(109[34:55])
    defparam i11860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_2_lut (.I0(PWMLimit[17]), .I1(n363), .I2(GND_net), .I3(GND_net), 
            .O(n35));
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48950_2_lut (.I0(n68615), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65546));
    defparam i48950_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50517_3_lut (.I0(n68825), .I1(n68807), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67533));
    defparam i50517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45850_3_lut (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[9] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62866));
    defparam i45850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45851_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62867));
    defparam i45851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11965_2_lut (.I0(byte_transmit_counter[1]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n27707));   // verilog/coms.v(109[34:55])
    defparam i11965_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i45872_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62888));
    defparam i45872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1433 (.I0(n54197), .I1(n54224), .I2(n58807), 
            .I3(n25800), .O(n14_adj_5567));
    defparam i6_4_lut_adj_1433.LUT_INIT = 16'h9669;
    SB_LUT4 i45873_4_lut (.I0(n62888), .I1(n27707), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][5] ), .O(n62889));
    defparam i45873_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i45871_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62887));
    defparam i45871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1434 (.I0(n58568), .I1(n14_adj_5567), .I2(n6_adj_5532), 
            .I3(\data_out_frame[20] [5]), .O(n58916));
    defparam i7_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1435 (.I0(n53169), .I1(n58791), .I2(n58377), 
            .I3(\data_out_frame[20] [0]), .O(n10_adj_5568));
    defparam i4_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i49278_2_lut (.I0(n68735), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65559));
    defparam i49278_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50519_3_lut (.I0(n68819), .I1(n68801), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67535));
    defparam i50519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45902_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62918));
    defparam i45902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45901_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62917));
    defparam i45901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1436 (.I0(n58412), .I1(\data_out_frame[21] [7]), 
            .I2(n58916), .I3(GND_net), .O(n58397));
    defparam i2_3_lut_adj_1436.LUT_INIT = 16'h9696;
    SB_LUT4 i48869_2_lut (.I0(n68747), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65591));
    defparam i48869_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50553_3_lut (.I0(n69005), .I1(n68753), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n67569));
    defparam i50553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n57819));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16]_c [0]), .C(clk16MHz), 
           .D(n31));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16]_c [1]), .C(clk16MHz), 
           .D(n57608));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n29495));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n29498));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n28969));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n28972));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16][4] ), .C(clk16MHz), 
           .D(n29501));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16][5] ), .C(clk16MHz), 
           .D(n29504));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n28976));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n28979));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n29507));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16][7] ), .C(clk16MHz), 
           .D(n29510));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17][0] ), .C(clk16MHz), 
           .D(n57380));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n29516));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n57378));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
           .D(n28982));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n57376));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n57374));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n57372));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n57370));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17]_c [7]), .C(clk16MHz), 
           .D(n57330));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n29537));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n57450));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n57430));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29546));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n57436));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29552));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n29555));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n57448));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29561));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29564));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29567));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29570));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n29577));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n57482));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29584));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29587));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20]_c [0]), .C(clk16MHz), 
           .D(n57292));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20][1] ), .C(clk16MHz), 
           .D(n29593));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n57304));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29599));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29602));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20][5] ), .C(clk16MHz), 
           .D(n29605));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20][6] ), .C(clk16MHz), 
           .D(n29608));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20]_c [7]), .C(clk16MHz), 
           .D(n57288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29948));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n28999), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29933));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29921));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i42088_3_lut (.I0(reset), .I1(n8_adj_5569), .I2(n58133), .I3(GND_net), 
            .O(n27972));
    defparam i42088_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29614));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29617));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29620));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n28987));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21]_c [3]), .C(clk16MHz), 
           .D(n33_adj_5570));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n57414));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29630));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29633));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29638));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29641));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
           .D(n29644));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29648));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29655));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29658));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n57420));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29671));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29674));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29677));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23][0] ), .C(clk16MHz), 
           .D(n57356));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23][1] ), .C(clk16MHz), 
           .D(n57354));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23][2] ), .C(clk16MHz), 
           .D(n57350));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n57302));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n57300));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29864));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23][6] ), .C(clk16MHz), 
           .D(n57346));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23][7] ), .C(clk16MHz), 
           .D(n29704));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2]_c [2]), .C(clk16MHz), 
           .D(n57442));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2][3] ), .C(clk16MHz), 
           .D(n28993));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2]_c [4]), .C(clk16MHz), 
           .D(n57424));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2][5] ), .C(clk16MHz), 
           .D(n29000));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2]_c [6]), .C(clk16MHz), 
           .D(n57444));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29855), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29854), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29853), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29852), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29851), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29850), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29849), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29848), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29847), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29846), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29845), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29844), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29843), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29842), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29841), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29840), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29839), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29838), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29837), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29836), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29835), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29834), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2]_c [7]), .C(clk16MHz), 
           .D(n57446));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29832), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29831), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29830), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29829), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29828), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29827), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29826), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29825), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29824), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29823), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29822), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29821), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29820), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29819), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29818), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29817), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29816), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29815), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29814), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29813), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29812), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29811), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29810), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29809), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29808), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29807), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29806), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29805), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29804), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29803), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29802), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29801), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29800), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29799), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29798), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29797), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29796), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29795), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29794), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29793), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29792), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29791), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29790), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29789), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29788), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29787), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29786), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29785), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29784), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29783), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29782), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29781), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29780), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29779), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29778));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29777));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29776));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29775));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29774));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29773));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29772));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29771));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29770));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29769));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29768));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29767));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29766));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29765));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29764));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29763));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29762));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29761));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29760));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29759));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29758));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29757));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29756));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29755));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29754));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29753));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29752));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n29751));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n29750));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n29749));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n29748));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n29747));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n29746));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n29745));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n29744));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n29743));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29742));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29741));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29740));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29739));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29738));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29737));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29736));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29735));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit_c[15]), .C(clk16MHz), 
           .D(n29734));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29733), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n29732), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n29731), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n29730), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n29729), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n29728), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n29727), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n29726), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n29725), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n29724), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n29723), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n29722), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n29721), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n29720), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n29719), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n29718), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n29717), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n3014), .D(n2_adj_5571), .S(n57887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n29716), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n29715), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n29714), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n29713), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n29712), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
           .D(n29009));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n29013));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
           .D(n29020));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
           .D(n29024));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1437 (.I0(n54293), .I1(n58412), .I2(n58774), 
            .I3(n53880), .O(n22_adj_5572));
    defparam i9_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i4_3_lut_4_lut (.I0(n53055), .I1(\data_out_frame[23] [1]), .I2(\data_out_frame[24] [7]), 
            .I3(n25645), .O(n11_adj_5512));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1438 (.I0(n60594), .I1(n22_adj_5572), .I2(n16_adj_5573), 
            .I3(n58807), .O(n24_adj_5574));
    defparam i11_4_lut_adj_1438.LUT_INIT = 16'h9669;
    SB_LUT4 n68732_bdd_4_lut (.I0(n68732), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n68735));
    defparam n68732_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1439 (.I0(\data_out_frame[21] [6]), .I1(n24_adj_5574), 
            .I2(n20_adj_5575), .I3(n54307), .O(n54259));
    defparam i12_4_lut_adj_1439.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3][4] ), .C(clk16MHz), 
           .D(n29028));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1440 (.I0(n58222), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(n58647), .O(n10_adj_5576));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i51349_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[4] [1]), .I2(n7_adj_7), 
            .I3(GND_net), .O(n57494));   // verilog/coms.v(94[13:20])
    defparam i51349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42090_3_lut (.I0(reset), .I1(n8_adj_5578), .I2(n58133), .I3(GND_net), 
            .O(n7_adj_7));
    defparam i42090_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i51351_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[4] [0]), .I2(n7_adj_7), 
            .I3(GND_net), .O(n57510));   // verilog/coms.v(94[13:20])
    defparam i51351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1441 (.I0(\data_out_frame[15] [5]), .I1(n10_adj_5576), 
            .I2(\data_out_frame[18] [0]), .I3(GND_net), .O(n53880));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1442 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n53880), .I3(GND_net), .O(n60272));
    defparam i2_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n28986), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1934__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n27640), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n27642), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n27644), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n27646), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n27648), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n27650), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n27652), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n27654), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n27656), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n27658), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n27660), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n27662), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n27664), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n27666), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n27668), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n27670), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n27672), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n27674), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n27676), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n27678), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n27680), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n27682), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n27684), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n27686), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n27688), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n27690), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n27692), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n27694), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n27696), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n27698), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1934__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n27700), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i13313_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n29056));   // verilog/coms.v(130[12] 305[6])
    defparam i13313_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13298_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29041));   // verilog/coms.v(130[12] 305[6])
    defparam i13298_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3]_c [5]), .C(clk16MHz), 
           .D(n29580));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(reset), 
            .I2(n32797), .I3(GND_net), .O(n22373));
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
           .D(n29044));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13344_3_lut (.I0(\data_in_frame[3]_c [7]), .I1(rx_data[7]), 
            .I2(n27968), .I3(GND_net), .O(n29087));   // verilog/coms.v(130[12] 305[6])
    defparam i13344_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13314_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n29057));   // verilog/coms.v(130[12] 305[6])
    defparam i13314_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13315_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n29058));   // verilog/coms.v(130[12] 305[6])
    defparam i13315_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13316_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n29059));   // verilog/coms.v(130[12] 305[6])
    defparam i13316_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13317_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n29060));   // verilog/coms.v(130[12] 305[6])
    defparam i13317_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n28985), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13318_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n29061));   // verilog/coms.v(130[12] 305[6])
    defparam i13318_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13319_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n29062));   // verilog/coms.v(130[12] 305[6])
    defparam i13319_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13320_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n29063));   // verilog/coms.v(130[12] 305[6])
    defparam i13320_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13321_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n29064));   // verilog/coms.v(130[12] 305[6])
    defparam i13321_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13322_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n29065));   // verilog/coms.v(130[12] 305[6])
    defparam i13322_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13323_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n29066));   // verilog/coms.v(130[12] 305[6])
    defparam i13323_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13324_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n29067));   // verilog/coms.v(130[12] 305[6])
    defparam i13324_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13325_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n29068));   // verilog/coms.v(130[12] 305[6])
    defparam i13325_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13326_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n29069));   // verilog/coms.v(130[12] 305[6])
    defparam i13326_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_776_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[14] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1443 (.I0(n2095), .I1(n2092), .I2(n2098), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n60080));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1443.LUT_INIT = 16'h8000;
    SB_LUT4 i13327_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n29070));   // verilog/coms.v(130[12] 305[6])
    defparam i13327_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13328_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n29071));   // verilog/coms.v(130[12] 305[6])
    defparam i13328_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13329_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n29072));   // verilog/coms.v(130[12] 305[6])
    defparam i13329_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13330_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n29073));   // verilog/coms.v(130[12] 305[6])
    defparam i13330_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13331_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n29074));   // verilog/coms.v(130[12] 305[6])
    defparam i13331_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13332_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n29075));   // verilog/coms.v(130[12] 305[6])
    defparam i13332_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13333_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n29076));   // verilog/coms.v(130[12] 305[6])
    defparam i13333_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13334_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n29077));   // verilog/coms.v(130[12] 305[6])
    defparam i13334_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1444 (.I0(\data_out_frame[21] [7]), .I1(n26288), 
            .I2(GND_net), .I3(GND_net), .O(n58894));
    defparam i1_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1445 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[22] [0]), 
            .I2(n53279), .I3(GND_net), .O(n53283));
    defparam i2_3_lut_adj_1445.LUT_INIT = 16'h9696;
    SB_LUT4 i1319_2_lut (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2107));   // verilog/coms.v(74[16:27])
    defparam i1319_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(\data_out_frame[22] [2]), .I1(n53279), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5579));
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'h6666;
    SB_LUT4 i13335_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n29078));   // verilog/coms.v(130[12] 305[6])
    defparam i13335_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1447 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(n2107), .I3(n6_adj_5579), .O(n58568));
    defparam i4_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1448 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58784));
    defparam i1_2_lut_adj_1448.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1449 (.I0(\data_out_frame[19] [5]), .I1(n58784), 
            .I2(n58377), .I3(n54293), .O(n7_adj_5580));
    defparam i2_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1450 (.I0(n7_adj_5580), .I1(n53283), .I2(n54324), 
            .I3(n58894), .O(n23340));
    defparam i4_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1451 (.I0(\data_in_frame[3]_c [5]), .I1(n58162), 
            .I2(n58565), .I3(n58455), .O(n53274));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut_adj_1451.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1452 (.I0(n54224), .I1(n58568), .I2(\data_out_frame[22] [3]), 
            .I3(GND_net), .O(n58318));
    defparam i2_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1453 (.I0(\data_out_frame[17] [7]), .I1(n58707), 
            .I2(GND_net), .I3(GND_net), .O(n58222));
    defparam i1_2_lut_adj_1453.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58686));
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1455 (.I0(n58641), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[13] [7]), .I3(n58686), .O(n10_adj_5581));
    defparam i4_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1456 (.I0(\data_out_frame[15] [7]), .I1(n58641), 
            .I2(n58222), .I3(n54253), .O(n53164));
    defparam i3_4_lut_adj_1456.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1457 (.I0(n53164), .I1(\data_out_frame[18] [1]), 
            .I2(n60075), .I3(GND_net), .O(n60594));
    defparam i2_3_lut_adj_1457.LUT_INIT = 16'h6969;
    SB_LUT4 i51341_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[20]_c [7]), 
            .I2(n28002), .I3(GND_net), .O(n57288));   // verilog/coms.v(94[13:20])
    defparam i51341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1458 (.I0(n54278), .I1(n53721), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n25947));
    defparam i2_3_lut_adj_1458.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1459 (.I0(\data_out_frame[20] [3]), .I1(n60594), 
            .I2(GND_net), .I3(GND_net), .O(n54197));
    defparam i1_2_lut_adj_1459.LUT_INIT = 16'h9999;
    SB_LUT4 i13336_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n29079));   // verilog/coms.v(130[12] 305[6])
    defparam i13336_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1460 (.I0(n54259), .I1(n58397), .I2(GND_net), 
            .I3(GND_net), .O(n58398));
    defparam i1_2_lut_adj_1460.LUT_INIT = 16'h6666;
    SB_LUT4 i13337_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n29080));   // verilog/coms.v(130[12] 305[6])
    defparam i13337_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(n58689), .I1(n58398), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5582));
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1462 (.I0(\data_out_frame[22] [4]), .I1(n58318), 
            .I2(\data_out_frame[25] [7]), .I3(n23340), .O(n12_adj_5583));
    defparam i5_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_209_i3_4_lut (.I0(n23344), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5583), .I3(n8_adj_5582), .O(n3_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13338_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n29081));   // verilog/coms.v(130[12] 305[6])
    defparam i13338_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13339_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n29082));   // verilog/coms.v(130[12] 305[6])
    defparam i13339_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_3_lut_adj_1463 (.I0(rx_data[2]), .I1(\data_in_frame[20] [2]), 
            .I2(n28002), .I3(GND_net), .O(n57304));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1463.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1464 (.I0(\data_out_frame[15] [1]), .I1(n53121), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[17] [2]), 
            .O(n58623));
    defparam i3_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i13340_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n29083));   // verilog/coms.v(130[12] 305[6])
    defparam i13340_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_5584));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i42104_3_lut (.I0(reset), .I1(n8_adj_5578), .I2(n38022), .I3(GND_net), 
            .O(n28002));
    defparam i42104_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1465 (.I0(\data_out_frame[19] [3]), .I1(n58623), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5585));
    defparam i1_2_lut_adj_1465.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1466 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n25154), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_5586));
    defparam i1_3_lut_4_lut_adj_1466.LUT_INIT = 16'hfefc;
    SB_LUT4 i51342_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[20]_c [0]), 
            .I2(n28002), .I3(GND_net), .O(n57292));   // verilog/coms.v(94[13:20])
    defparam i51342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1467 (.I0(\data_out_frame[21] [4]), .I1(n26199), 
            .I2(n26431), .I3(n6_adj_5585), .O(n53721));
    defparam i4_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1468 (.I0(n53721), .I1(n54324), .I2(\data_out_frame[21] [5]), 
            .I3(GND_net), .O(n58777));
    defparam i2_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 i13341_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n29084));   // verilog/coms.v(130[12] 305[6])
    defparam i13341_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58605));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1470 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3545[0]), .I3(n39337), .O(n25082));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1470.LUT_INIT = 16'ha8aa;
    SB_LUT4 i3_4_lut_adj_1471 (.I0(n58273), .I1(n58949), .I2(n58922), 
            .I3(n58662), .O(n25666));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i51544_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n39337), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i51544_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i2_3_lut_4_lut_adj_1472 (.I0(\data_in_frame[0] [7]), .I1(n25466), 
            .I2(n58614), .I3(n58659), .O(n8_adj_5477));
    defparam i2_3_lut_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\data_out_frame[17] [0]), .I1(n58207), 
            .I2(GND_net), .I3(GND_net), .O(n26431));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 i13342_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n29085));   // verilog/coms.v(130[12] 305[6])
    defparam i13342_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13343_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n29086));   // verilog/coms.v(130[12] 305[6])
    defparam i13343_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1474 (.I0(\data_out_frame[16] [0]), .I1(n25830), 
            .I2(GND_net), .I3(GND_net), .O(n58771));
    defparam i1_2_lut_adj_1474.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1475 (.I0(\data_out_frame[15] [5]), .I1(n53285), 
            .I2(GND_net), .I3(GND_net), .O(n58495));
    defparam i1_2_lut_adj_1475.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1476 (.I0(\data_out_frame[19] [0]), .I1(n40_adj_5587), 
            .I2(n54253), .I3(n54237), .O(n10_adj_5588));
    defparam i4_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1477 (.I0(n68374), .I1(n10_adj_5588), .I2(n53999), 
            .I3(n2076), .O(n58440));
    defparam i5_4_lut_adj_1477.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58273));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1479 (.I0(n26088), .I1(n58638), .I2(n58273), 
            .I3(\data_out_frame[11] [7]), .O(n24670));   // verilog/coms.v(74[16:62])
    defparam i3_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1480 (.I0(\data_out_frame[12] [1]), .I1(n24670), 
            .I2(GND_net), .I3(GND_net), .O(n58443));
    defparam i1_2_lut_adj_1480.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1481 (.I0(\data_out_frame[16] [3]), .I1(n25673), 
            .I2(\data_out_frame[16] [7]), .I3(\data_out_frame[16] [5]), 
            .O(n40_adj_5587));
    defparam i3_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1482 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25673));
    defparam i1_2_lut_adj_1482.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1483 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25992));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1483.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n58635));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1485 (.I0(n26235), .I1(n58704), .I2(\data_out_frame[13] [4]), 
            .I3(\data_out_frame[7] [1]), .O(n12_adj_5589));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1486 (.I0(n24827), .I1(n12_adj_5589), .I2(n58838), 
            .I3(n38), .O(n53285));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1487 (.I0(n1130), .I1(\data_out_frame[6] [6]), 
            .I2(n58644), .I3(n25656), .O(n10_adj_5590));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1488 (.I0(n25763), .I1(n10_adj_5590), .I2(\data_out_frame[9] [2]), 
            .I3(GND_net), .O(n58561));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1488.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[13] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(\data_out_frame[15] [6]), .I1(n53285), 
            .I2(GND_net), .I3(GND_net), .O(n58491));
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26235));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1491 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58838));
    defparam i1_2_lut_adj_1491.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1492 (.I0(n58650), .I1(n58242), .I2(n58838), 
            .I3(GND_net), .O(n8_adj_5591));
    defparam i3_3_lut_adj_1492.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1493 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[7] [3]), .I3(n4_adj_5592), .O(n28_adj_5593));
    defparam i12_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1494 (.I0(n58449), .I1(\data_out_frame[7] [4]), 
            .I2(n58189), .I3(\data_out_frame[6] [7]), .O(n26_adj_5594));
    defparam i10_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1495 (.I0(n58626), .I1(n58225), .I2(n58436), 
            .I3(\data_out_frame[6] [4]), .O(n27_adj_5595));
    defparam i11_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1496 (.I0(n58919), .I1(n58245), .I2(n25237), 
            .I3(\data_out_frame[7] [1]), .O(n25_adj_5596));
    defparam i9_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i19233_3_lut (.I0(n27968), .I1(rx_data[5]), .I2(\data_in_frame[3]_c [5]), 
            .I3(GND_net), .O(n29580));   // verilog/coms.v(94[13:20])
    defparam i19233_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1497 (.I0(n25996), .I1(n25663), .I2(n8_adj_5591), 
            .I3(\data_out_frame[9] [1]), .O(n6_adj_5597));
    defparam i1_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1498 (.I0(n25_adj_5596), .I1(n27_adj_5595), .I2(n26_adj_5594), 
            .I3(n28_adj_5593), .O(n60866));
    defparam i15_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1499 (.I0(n60866), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[7] [5]), .I3(n6_adj_5597), .O(n60941));
    defparam i4_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1500 (.I0(n60941), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [7]), .I3(\data_out_frame[10] [0]), 
            .O(n10_adj_5598));
    defparam i4_4_lut_adj_1500.LUT_INIT = 16'h9669;
    SB_LUT4 i13242_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16]_c [0]), 
            .I3(deadband[0]), .O(n28985));   // verilog/coms.v(148[4] 304[11])
    defparam i13242_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1501 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[11] [5]), .I3(n58166), .O(n14_adj_5599));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1502 (.I0(n58312), .I1(n14_adj_5599), .I2(n10_adj_5600), 
            .I3(\data_out_frame[11] [1]), .O(n54182));   // verilog/coms.v(88[17:63])
    defparam i7_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1503 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[8][4] ), 
            .I2(n58579), .I3(n25237), .O(n58828));
    defparam i3_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 i13243_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n28986));   // verilog/coms.v(148[4] 304[11])
    defparam i13243_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1504 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[8][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n58446));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1504.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1505 (.I0(\data_out_frame[6] [3]), .I1(n58343), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n25996));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1505.LUT_INIT = 16'h9696;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_776_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5571));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1506 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[10] [3]), .I3(n58683), .O(n10_adj_5600));   // verilog/coms.v(88[17:63])
    defparam i2_2_lut_3_lut_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1507 (.I0(n58680), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[13] [3]), .I3(n58704), .O(n10_adj_5601));
    defparam i4_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1508 (.I0(\data_out_frame[9] [1]), .I1(n10_adj_5601), 
            .I2(\data_out_frame[11] [2]), .I3(GND_net), .O(n25830));
    defparam i5_3_lut_adj_1508.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_1509 (.I0(\data_in_frame[17]_c [7]), .I1(n27920), 
            .I2(n27997), .I3(rx_data[7]), .O(n57330));
    defparam i13_4_lut_adj_1509.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13969_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n29712));   // verilog/coms.v(148[4] 304[11])
    defparam i13969_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1510 (.I0(reset), .I1(n38022), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n7_adj_5602), .O(n27994));
    defparam i2_3_lut_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1511 (.I0(n60532), .I1(n54278), .I2(\data_out_frame[23] [4]), 
            .I3(\data_out_frame[23] [6]), .O(n5_adj_5603));
    defparam i1_2_lut_4_lut_adj_1511.LUT_INIT = 16'h9669;
    SB_LUT4 i19758_3_lut (.I0(current_limit_c[15]), .I1(\data_in_frame[20]_c [7]), 
            .I2(n22362), .I3(GND_net), .O(n29734));
    defparam i19758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1512 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25663));
    defparam i1_2_lut_adj_1512.LUT_INIT = 16'h6666;
    SB_LUT4 i19759_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20]_c [0]), 
            .I2(n22362), .I3(GND_net), .O(n29741));
    defparam i19759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19583_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21]_c [3]), 
            .I2(n22362), .I3(GND_net), .O(n29746));
    defparam i19583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1513 (.I0(\data_out_frame[15] [5]), .I1(n53285), 
            .I2(\data_out_frame[16] [0]), .I3(n25830), .O(n54253));
    defparam i1_2_lut_4_lut_adj_1513.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58189));
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1515 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(n58189), .I3(n25456), .O(n58644));
    defparam i3_4_lut_adj_1515.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1516 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[10] [2]), .O(n58835));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i13970_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n29713));   // verilog/coms.v(148[4] 304[11])
    defparam i13970_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(\data_out_frame[7] [1]), .I1(n25656), 
            .I2(GND_net), .I3(GND_net), .O(n26100));
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1518 (.I0(n24827), .I1(n26100), .I2(n25663), 
            .I3(n1312), .O(n58475));
    defparam i3_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1519 (.I0(\data_out_frame[11] [6]), .I1(n26085), 
            .I2(n25639), .I3(\data_out_frame[14] [0]), .O(n58370));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1520 (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[6] [0]), .I3(n1191), .O(n58231));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i48823_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65506));   // verilog/coms.v(158[12:15])
    defparam i48823_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58662));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i48817_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65503));   // verilog/coms.v(158[12:15])
    defparam i48817_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1522 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58845));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1522.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1523 (.I0(\data_out_frame[13] [0]), .I1(n58845), 
            .I2(n58343), .I3(\data_out_frame[4] [2]), .O(n10_adj_5604));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1523.LUT_INIT = 16'h6996;
    SB_LUT4 i13971_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n29714));   // verilog/coms.v(148[4] 304[11])
    defparam i13971_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48816_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65501));   // verilog/coms.v(158[12:15])
    defparam i48816_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1524 (.I0(n58882), .I1(\data_in_frame[14] [0]), 
            .I2(n25335), .I3(\data_in_frame[16]_c [1]), .O(n14_adj_5605));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1525 (.I0(\data_out_frame[15] [7]), .I1(n53666), 
            .I2(GND_net), .I3(GND_net), .O(n58585));
    defparam i1_2_lut_adj_1525.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5592));
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1527 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n58216));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i48809_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65500));   // verilog/coms.v(158[12:15])
    defparam i48809_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49292_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65499));   // verilog/coms.v(158[12:15])
    defparam i49292_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1528 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58449));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1528.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1529 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n43_adj_5494));
    defparam i1_2_lut_3_lut_adj_1529.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1530 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58650));
    defparam i1_2_lut_adj_1530.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_out_frame[9] [4]), .I1(n1312), 
            .I2(GND_net), .I3(GND_net), .O(n26085));
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1532 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n58197));   // verilog/coms.v(74[16:62])
    defparam i2_3_lut_adj_1532.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1533 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n58242));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1533.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1534 (.I0(\data_out_frame[7] [4]), .I1(n58276), 
            .I2(n58242), .I3(\data_out_frame[5] [1]), .O(n25639));   // verilog/coms.v(76[16:34])
    defparam i3_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1535 (.I0(\data_out_frame[10] [0]), .I1(n25639), 
            .I2(GND_net), .I3(GND_net), .O(n26088));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1535.LUT_INIT = 16'h6666;
    SB_LUT4 i13972_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n29715));   // verilog/coms.v(148[4] 304[11])
    defparam i13972_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58629));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1537 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(GND_net), .I3(GND_net), .O(n25259));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1538 (.I0(n58197), .I1(n26085), .I2(n58650), 
            .I3(n58742), .O(n15_adj_5606));   // verilog/coms.v(74[16:62])
    defparam i6_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1539 (.I0(n15_adj_5606), .I1(n58629), .I2(n14_adj_5607), 
            .I3(\data_out_frame[7] [6]), .O(n58254));   // verilog/coms.v(74[16:62])
    defparam i8_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [5]), 
            .I2(n58828), .I3(GND_net), .O(n22_adj_5608));
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1541 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n3579), .I3(n161), .O(n62));
    defparam i3_4_lut_adj_1541.LUT_INIT = 16'h2000;
    SB_LUT4 i13_4_lut_adj_1542 (.I0(n58585), .I1(\data_out_frame[8][6] ), 
            .I2(n58321), .I3(n1699), .O(n34_adj_5609));
    defparam i13_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i48804_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65495));   // verilog/coms.v(158[12:15])
    defparam i48804_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_4_lut_adj_1543 (.I0(\data_out_frame[14] [3]), .I1(n25269), 
            .I2(n25830), .I3(\data_out_frame[15] [4]), .O(n23_adj_5610));
    defparam i2_2_lut_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i48830_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65491));   // verilog/coms.v(158[12:15])
    defparam i48830_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13973_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n29716));   // verilog/coms.v(148[4] 304[11])
    defparam i13973_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i17_4_lut_adj_1544 (.I0(n23_adj_5610), .I1(n34_adj_5609), .I2(n54182), 
            .I3(n58925), .O(n38_adj_5611));
    defparam i17_4_lut_adj_1544.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1545 (.I0(n58491), .I1(n58562), .I2(n58258), 
            .I3(\data_out_frame[14] [1]), .O(n36));
    defparam i15_4_lut_adj_1545.LUT_INIT = 16'h9669;
    SB_LUT4 i19180_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n29717));   // verilog/coms.v(148[4] 304[11])
    defparam i19180_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut_adj_1546 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[14] [6]), .I3(n22_adj_5608), .O(n37));
    defparam i16_4_lut_adj_1546.LUT_INIT = 16'h6996;
    SB_LUT4 i48581_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65489));   // verilog/coms.v(158[12:15])
    defparam i48581_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14_4_lut_adj_1547 (.I0(\data_out_frame[15] [5]), .I1(n58617), 
            .I2(n58857), .I3(n58511), .O(n35_adj_5612));
    defparam i14_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35_adj_5612), .I1(n37), .I2(n36), .I3(n38_adj_5611), 
            .O(n53999));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1548 (.I0(n58216), .I1(\data_out_frame[12] [4]), 
            .I2(n58835), .I3(n58635), .O(n12_adj_5613));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1549 (.I0(\data_out_frame[4] [0]), .I1(n12_adj_5613), 
            .I2(n25992), .I3(\data_out_frame[14] [5]), .O(n60872));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i51358_4_lut (.I0(n58527), .I1(n54146), .I2(n60872), .I3(n40_adj_5587), 
            .O(n68374));
    defparam i51358_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i48766_2_lut (.I0(\data_out_frame[0][4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65443));
    defparam i48766_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1550 (.I0(n43_adj_5494), .I1(n68374), .I2(\data_out_frame[16] [4]), 
            .I3(n53999), .O(n10_adj_5614));
    defparam i4_4_lut_adj_1550.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1551 (.I0(\data_out_frame[18] [7]), .I1(n10_adj_5614), 
            .I2(\data_out_frame[19] [1]), .I3(GND_net), .O(n58151));
    defparam i5_3_lut_adj_1551.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25845));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1553 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58166));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1553.LUT_INIT = 16'h6666;
    SB_LUT4 i48701_2_lut (.I0(\data_out_frame[3][4] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65444));
    defparam i48701_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1554 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n58638));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1554.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1555 (.I0(\data_out_frame[5] [7]), .I1(n58638), 
            .I2(n58216), .I3(n58166), .O(n1513));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n58949));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(GND_net), .I3(GND_net), .O(n25814));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1558 (.I0(n25377), .I1(n58548), .I2(Kp_23__N_878), 
            .I3(n58363), .O(Kp_23__N_993));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1559 (.I0(n25377), .I1(n58548), .I2(n25370), 
            .I3(\data_in_frame[6] [7]), .O(n58620));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_5481));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n4_adj_5480));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1560 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n58617));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1560.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1561 (.I0(\data_out_frame[10] [0]), .I1(n25639), 
            .I2(\data_out_frame[14] [2]), .I3(\data_out_frame[12] [1]), 
            .O(n14_adj_5607));   // verilog/coms.v(74[16:62])
    defparam i5_3_lut_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25301));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 i48799_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65487));   // verilog/coms.v(158[12:15])
    defparam i48799_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13975_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n29718));   // verilog/coms.v(148[4] 304[11])
    defparam i13975_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48796_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65482));   // verilog/coms.v(158[12:15])
    defparam i48796_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1563 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n25656));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5478));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48951_2_lut (.I0(\data_out_frame[3][3] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65442));
    defparam i48951_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48794_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65481));   // verilog/coms.v(158[12:15])
    defparam i48794_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(n54253), .I1(n58608), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5615));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i48793_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65480));   // verilog/coms.v(158[12:15])
    defparam i48793_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1565 (.I0(\data_out_frame[21] [3]), .I1(n25845), 
            .I2(n58151), .I3(n6_adj_5615), .O(n54278));
    defparam i4_4_lut_adj_1565.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1566 (.I0(n58440), .I1(\data_out_frame[21] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5616));
    defparam i1_2_lut_adj_1566.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1567 (.I0(n58611), .I1(n26330), .I2(n26431), 
            .I3(n6_adj_5616), .O(n60532));
    defparam i4_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i48828_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65479));   // verilog/coms.v(158[12:15])
    defparam i48828_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1568 (.I0(n60532), .I1(n54278), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n53179));
    defparam i2_3_lut_adj_1568.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_3_lut_adj_1569 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26180));
    defparam i2_2_lut_3_lut_adj_1569.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_208_i3_4_lut (.I0(n5_adj_5603), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n58605), .I3(n58778), .O(n3_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i48666_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65476));   // verilog/coms.v(158[12:15])
    defparam i48666_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_776_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48820_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65465));   // verilog/coms.v(158[12:15])
    defparam i48820_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48765_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65451));   // verilog/coms.v(158[12:15])
    defparam i48765_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48633_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65428));   // verilog/coms.v(158[12:15])
    defparam i48633_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_776_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[19] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1570 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[10] [4]), 
            .I2(n10_adj_5604), .I3(n58231), .O(n53121));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_3_lut_adj_1571 (.I0(rx_data[1]), .I1(\data_in_frame[16]_c [1]), 
            .I2(n27994), .I3(GND_net), .O(n57608));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1571.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1572 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_5531));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_adj_1572.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_3_lut_adj_1573 (.I0(n10_adj_5531), .I1(n27913), .I2(n161), 
            .I3(GND_net), .O(n38022));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1573.LUT_INIT = 16'hefef;
    SB_LUT4 select_776_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i39_3_lut (.I0(n27994), .I1(rx_data[0]), .I2(\data_in_frame[16]_c [0]), 
            .I3(GND_net), .O(n31));   // verilog/coms.v(94[13:20])
    defparam i39_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13976_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n29719));   // verilog/coms.v(148[4] 304[11])
    defparam i13976_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13977_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n29720));   // verilog/coms.v(148[4] 304[11])
    defparam i13977_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [2]), 
            .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'ha088;
    SB_LUT4 select_776_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13978_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n29721));   // verilog/coms.v(148[4] 304[11])
    defparam i13978_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48736_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65401));   // verilog/coms.v(158[12:15])
    defparam i48736_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_776_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13979_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n29722));   // verilog/coms.v(148[4] 304[11])
    defparam i13979_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1575 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[6] [2]), .O(n58579));
    defparam i1_2_lut_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5566));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13980_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n29723));   // verilog/coms.v(148[4] 304[11])
    defparam i13980_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [2]), 
            .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'ha088;
    SB_LUT4 i5_3_lut_4_lut_adj_1577 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(n10_adj_5598), .I3(n25996), .O(n58683));
    defparam i5_3_lut_4_lut_adj_1577.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48735_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65400));   // verilog/coms.v(158[12:15])
    defparam i48735_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [7]), 
            .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'ha088;
    SB_LUT4 select_776_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_306_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5617));   // verilog/coms.v(157[7:23])
    defparam equal_306_i7_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i48734_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65399));   // verilog/coms.v(158[12:15])
    defparam i48734_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [4]), 
            .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'ha088;
    SB_LUT4 select_776_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48720_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65398));   // verilog/coms.v(158[12:15])
    defparam i48720_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48718_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65395));   // verilog/coms.v(158[12:15])
    defparam i48718_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1580 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [2]), 
            .I2(\encoder0_position_scaled[18] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1580.LUT_INIT = 16'ha088;
    SB_LUT4 i48715_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65394));   // verilog/coms.v(158[12:15])
    defparam i48715_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48709_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65393));   // verilog/coms.v(158[12:15])
    defparam i48709_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13981_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n29724));   // verilog/coms.v(148[4] 304[11])
    defparam i13981_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[17] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48706_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65387));   // verilog/coms.v(158[12:15])
    defparam i48706_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_776_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[16] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48702_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65386));   // verilog/coms.v(158[12:15])
    defparam i48702_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13982_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n29725));   // verilog/coms.v(148[4] 304[11])
    defparam i13982_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13983_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n29726));   // verilog/coms.v(148[4] 304[11])
    defparam i13983_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[12] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13984_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n29727));   // verilog/coms.v(148[4] 304[11])
    defparam i13984_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48678_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65382));   // verilog/coms.v(158[12:15])
    defparam i48678_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13985_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n29728));   // verilog/coms.v(148[4] 304[11])
    defparam i13985_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19754_3_lut (.I0(current_limit_c[15]), .I1(\current[15] ), 
            .I2(n30), .I3(GND_net), .O(n296));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i19754_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i13986_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n29729));   // verilog/coms.v(148[4] 304[11])
    defparam i13986_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13987_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n29730));   // verilog/coms.v(148[4] 304[11])
    defparam i13987_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13988_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n29731));   // verilog/coms.v(148[4] 304[11])
    defparam i13988_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48670_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65379));   // verilog/coms.v(158[12:15])
    defparam i48670_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_776_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13989_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n29732));   // verilog/coms.v(148[4] 304[11])
    defparam i13989_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13990_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n29733));   // verilog/coms.v(148[4] 304[11])
    defparam i13990_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48658_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65374));   // verilog/coms.v(158[12:15])
    defparam i48658_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48655_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65373));   // verilog/coms.v(158[12:15])
    defparam i48655_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48803_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65372));   // verilog/coms.v(158[12:15])
    defparam i48803_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14036_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n29779));   // verilog/coms.v(148[4] 304[11])
    defparam i14036_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12171_1_lut (.I0(n3579), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n27913));   // verilog/coms.v(148[4] 304[11])
    defparam i12171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i4_3_lut (.I0(\data_out_frame[4] [3]), 
            .I1(\data_out_frame[5] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n4_adj_5457));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_776_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19105_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n29780));   // verilog/coms.v(148[4] 304[11])
    defparam i19105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i19127_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n29781));   // verilog/coms.v(148[4] 304[11])
    defparam i19127_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14039_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n29782));   // verilog/coms.v(148[4] 304[11])
    defparam i14039_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14040_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n29783));   // verilog/coms.v(148[4] 304[11])
    defparam i14040_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14041_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n29784));   // verilog/coms.v(148[4] 304[11])
    defparam i14041_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5345_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n2092), 
            .I2(n60003), .I3(n4452), .O(n20750));   // verilog/coms.v(148[4] 304[11])
    defparam i5345_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i19179_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n29785));   // verilog/coms.v(148[4] 304[11])
    defparam i19179_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n20750), .I1(n2092), .I2(n22366), .I3(n62488), 
            .O(n27160));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'hbbba;
    SB_LUT4 i464_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2201));   // verilog/coms.v(148[4] 304[11])
    defparam i464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19028_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n29786));   // verilog/coms.v(148[4] 304[11])
    defparam i19028_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18979_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5]_c [7]), 
            .I3(\Ki[7] ), .O(n29787));   // verilog/coms.v(148[4] 304[11])
    defparam i18979_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14045_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5][6] ), 
            .I3(\Ki[6] ), .O(n29788));   // verilog/coms.v(148[4] 304[11])
    defparam i14045_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i45468_4_lut (.I0(n2092), .I1(n2095), .I2(n3303), .I3(n2098), 
            .O(n62469));   // verilog/coms.v(139[4] 141[7])
    defparam i45468_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1582 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n2095), 
            .I2(n62469), .I3(n60217), .O(n57202));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'hb3a0;
    SB_LUT4 select_776_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5338_4_lut (.I0(n2096), .I1(\FRAME_MATCHER.state[3] ), .I2(n2098), 
            .I3(n25082), .O(n20741));   // verilog/coms.v(148[4] 304[11])
    defparam i5338_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i453_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2190));   // verilog/coms.v(148[4] 304[11])
    defparam i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i452_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2189));   // verilog/coms.v(148[4] 304[11])
    defparam i452_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19029_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5]_c [5]), 
            .I3(\Ki[5] ), .O(n29789));   // verilog/coms.v(148[4] 304[11])
    defparam i19029_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23336_4_lut (.I0(n5_adj_5586), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [2]), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i23336_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i14047_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n29790));   // verilog/coms.v(148[4] 304[11])
    defparam i14047_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 equal_308_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5602));   // verilog/coms.v(157[7:23])
    defparam equal_308_i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(\FRAME_MATCHER.i [4]), .I1(n25154), .I2(GND_net), 
            .I3(GND_net), .O(n25001));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'heeee;
    SB_LUT4 i23339_4_lut (.I0(n8_adj_5584), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25001), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i23339_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i14048_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5][3] ), 
            .I3(\Ki[3] ), .O(n29791));   // verilog/coms.v(148[4] 304[11])
    defparam i14048_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48801_2_lut (.I0(\data_out_frame[9] [0]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65490));
    defparam i48801_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i9_3_lut (.I0(\data_out_frame[10] [0]), 
            .I1(\data_out_frame[11] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n9_adj_5565));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1584 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n22366));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1584.LUT_INIT = 16'h4444;
    SB_LUT4 i14049_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5][2] ), 
            .I3(\Ki[2] ), .O(n29792));   // verilog/coms.v(148[4] 304[11])
    defparam i14049_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_2_lut (.I0(n25082), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n26612));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1585 (.I0(n4452), .I1(n26612), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n22366), .O(n60942));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1585.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(n25090), .I1(n2098), .I2(n2096), .I3(n60942), 
            .O(n26617));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'hbaaa;
    SB_LUT4 i14050_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n29793));   // verilog/coms.v(148[4] 304[11])
    defparam i14050_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_2_lut_adj_1587 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5619));
    defparam i2_2_lut_adj_1587.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1588 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5620));
    defparam i6_4_lut_adj_1588.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1589 (.I0(\data_in[3] [6]), .I1(n14_adj_5620), 
            .I2(n10_adj_5619), .I3(\data_in[2] [1]), .O(n25127));
    defparam i7_4_lut_adj_1589.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1590 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n25127), .I3(\data_in[0] [1]), .O(n20_adj_5621));
    defparam i8_4_lut_adj_1590.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1591 (.I0(n25029), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_5622));
    defparam i7_4_lut_adj_1591.LUT_INIT = 16'hfeff;
    SB_LUT4 i14051_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [7]), 
            .I3(\Kp[15] ), .O(n29794));   // verilog/coms.v(148[4] 304[11])
    defparam i14051_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i45644_4_lut (.I0(\data_in[1] [3]), .I1(\data_in[0] [5]), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n62651));
    defparam i45644_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_1592 (.I0(n62651), .I1(n19_adj_5622), .I2(n20_adj_5621), 
            .I3(GND_net), .O(n2092));
    defparam i11_3_lut_adj_1592.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1593 (.I0(\data_in[2] [4]), .I1(n25127), .I2(\data_in[1] [5]), 
            .I3(n25157), .O(n18));
    defparam i7_4_lut_adj_1593.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1594 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n25096), .O(n20_adj_5623));
    defparam i9_4_lut_adj_1594.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_1595 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5624));
    defparam i4_2_lut_adj_1595.LUT_INIT = 16'heeee;
    SB_LUT4 i14052_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [6]), 
            .I3(\Kp[14] ), .O(n29795));   // verilog/coms.v(148[4] 304[11])
    defparam i14052_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1596 (.I0(n58495), .I1(n58771), .I2(n53999), 
            .I3(GND_net), .O(n58527));
    defparam i1_2_lut_3_lut_adj_1596.LUT_INIT = 16'h6969;
    SB_LUT4 i14053_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2][5] ), 
            .I3(\Kp[13] ), .O(n29796));   // verilog/coms.v(148[4] 304[11])
    defparam i14053_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19450_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [4]), 
            .I3(\Kp[12] ), .O(n29797));   // verilog/coms.v(148[4] 304[11])
    defparam i19450_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14055_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2][3] ), 
            .I3(\Kp[11] ), .O(n29798));   // verilog/coms.v(148[4] 304[11])
    defparam i14055_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut_adj_1597 (.I0(n15_adj_5624), .I1(n20_adj_5623), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n2095));
    defparam i10_4_lut_adj_1597.LUT_INIT = 16'hfeff;
    SB_LUT4 i4_4_lut_adj_1598 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5625));
    defparam i4_4_lut_adj_1598.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1599 (.I0(\data_in[3] [4]), .I1(n10_adj_5625), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n25157));
    defparam i5_3_lut_adj_1599.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1600 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5626));
    defparam i6_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1601 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [7]), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1601.LUT_INIT = 16'ha088;
    SB_LUT4 i7_4_lut_adj_1602 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_5627));
    defparam i7_4_lut_adj_1602.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1603 (.I0(n17_adj_5627), .I1(\data_in[1] [6]), 
            .I2(n16_adj_5626), .I3(\data_in[3] [7]), .O(n25096));
    defparam i9_4_lut_adj_1603.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_adj_1604 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5628));
    defparam i5_3_lut_adj_1604.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1605 (.I0(\data_in[0] [6]), .I1(n25157), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5629));
    defparam i6_4_lut_adj_1605.LUT_INIT = 16'hfeff;
    SB_LUT4 select_776_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14056_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [2]), 
            .I3(\Kp[10] ), .O(n29799));   // verilog/coms.v(148[4] 304[11])
    defparam i14056_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8_4_lut_adj_1606 (.I0(n15_adj_5629), .I1(\data_in[3] [0]), 
            .I2(n14_adj_5628), .I3(\data_in[2] [2]), .O(n25029));
    defparam i8_4_lut_adj_1606.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1607 (.I0(n25029), .I1(\data_in[0] [7]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [6]), .O(n16_adj_5630));
    defparam i6_4_lut_adj_1607.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1608 (.I0(n25096), .I1(\data_in[2] [1]), .I2(\data_in[3] [3]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5631));
    defparam i7_4_lut_adj_1608.LUT_INIT = 16'hbfff;
    SB_LUT4 select_776_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i9_4_lut_adj_1609 (.I0(n17_adj_5631), .I1(\data_in[2] [3]), 
            .I2(n16_adj_5630), .I3(\data_in[3] [5]), .O(n2098));
    defparam i9_4_lut_adj_1609.LUT_INIT = 16'hfbff;
    SB_LUT4 i370_2_lut (.I0(n2095), .I1(n2092), .I2(GND_net), .I3(GND_net), 
            .O(n2096));   // verilog/coms.v(142[4] 144[7])
    defparam i370_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1610 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(GND_net), .I3(GND_net), .O(n32799));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1610.LUT_INIT = 16'heeee;
    SB_LUT4 i23171_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), .I2(GND_net), 
            .I3(GND_net), .O(n38817));
    defparam i23171_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1611 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5632));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1611.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(byte_transmit_counter[4]), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_5633));
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'ha8a0;
    SB_LUT4 select_776_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23687_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5633), .I3(n4_adj_5632), .O(n39337));
    defparam i23687_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 select_776_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_adj_1613 (.I0(n39337), .I1(n60080), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(n38817), .O(n6_adj_5634));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1613.LUT_INIT = 16'hccec;
    SB_LUT4 i3_4_lut_adj_1614 (.I0(n32799), .I1(n6_adj_5634), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n69037));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1614.LUT_INIT = 16'hefee;
    SB_LUT4 select_776_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1615 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n58511), .I3(GND_net), .O(n54237));
    defparam i1_2_lut_3_lut_adj_1615.LUT_INIT = 16'h9696;
    SB_LUT4 i48865_2_lut (.I0(\data_out_frame[9] [2]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65441));
    defparam i48865_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21546_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n9_adj_5452));   // verilog/coms.v(105[12:33])
    defparam i21546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i12_3_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\data_out_frame[15] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n12_adj_5451));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i11_3_lut (.I0(\data_out_frame[12] [2]), 
            .I1(\data_out_frame[13] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n11_adj_5450));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49348_2_lut (.I0(\data_out_frame[9] [1]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65440));
    defparam i49348_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i9_3_lut (.I0(\data_out_frame[10] [1]), 
            .I1(\data_out_frame[11] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n9));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14057_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n29800));   // verilog/coms.v(148[4] 304[11])
    defparam i14057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i20082_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n29801));   // verilog/coms.v(148[4] 304[11])
    defparam i20082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1616 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3][3] ), .O(n25923));
    defparam i1_2_lut_3_lut_4_lut_adj_1616.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [4]), 
            .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'ha088;
    SB_LUT4 i18987_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3]_c [7]), 
            .I3(\Kp[7] ), .O(n29802));   // verilog/coms.v(148[4] 304[11])
    defparam i18987_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1618 (.I0(\data_out_frame[16] [6]), .I1(n58151), 
            .I2(n58495), .I3(n58771), .O(n58611));
    defparam i2_3_lut_4_lut_adj_1618.LUT_INIT = 16'h9669;
    SB_LUT4 select_776_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14060_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3] [6]), 
            .I3(\Kp[6] ), .O(n29803));   // verilog/coms.v(148[4] 304[11])
    defparam i14060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5293));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1619 (.I0(n54293), .I1(n53721), .I2(n54324), 
            .I3(\data_out_frame[21] [5]), .O(n58778));
    defparam i1_2_lut_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i12_3_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\data_out_frame[15] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n12_adj_5442));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_776_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5292));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1620 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n26199));
    defparam i1_2_lut_3_lut_adj_1620.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i11_3_lut (.I0(\data_out_frame[12] [1]), 
            .I1(\data_out_frame[13] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n11_adj_5441));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_776_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1621 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [1]), 
            .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5291));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1621.LUT_INIT = 16'ha088;
    SB_LUT4 i11858_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27598));   // verilog/coms.v(109[34:55])
    defparam i11858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45878_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62894));
    defparam i45878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45879_4_lut (.I0(n62894), .I1(n27598), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n62895));
    defparam i45879_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45877_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62893));
    defparam i45877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_776_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1622 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[20] [3]), 
            .I2(n60594), .I3(n25947), .O(n58689));
    defparam i2_3_lut_4_lut_adj_1622.LUT_INIT = 16'h9669;
    SB_LUT4 select_776_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5290));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [2]), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'ha088;
    SB_LUT4 i14061_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3]_c [5]), 
            .I3(\Kp[5] ), .O(n29804));   // verilog/coms.v(148[4] 304[11])
    defparam i14061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1624 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [1]), 
            .I2(\encoder0_position_scaled[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5429));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1624.LUT_INIT = 16'ha088;
    SB_LUT4 i14062_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][4] ), 
            .I3(\Kp[4] ), .O(n29805));   // verilog/coms.v(148[4] 304[11])
    defparam i14062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5425));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14063_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][3] ), 
            .I3(\Kp[3] ), .O(n29806));   // verilog/coms.v(148[4] 304[11])
    defparam i14063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_3_lut_4_lut_adj_1625 (.I0(\data_out_frame[15] [6]), .I1(n53285), 
            .I2(n10_adj_5581), .I3(n53666), .O(n60075));
    defparam i5_3_lut_4_lut_adj_1625.LUT_INIT = 16'h6996;
    SB_LUT4 i14064_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][2] ), 
            .I3(\Kp[2] ), .O(n29807));   // verilog/coms.v(148[4] 304[11])
    defparam i14064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[23] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5423));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14065_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n29808));   // verilog/coms.v(148[4] 304[11])
    defparam i14065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14066_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n29809));   // verilog/coms.v(148[4] 304[11])
    defparam i14066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51921 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n69002));
    defparam byte_transmit_counter_0__bdd_4_lut_51921.LUT_INIT = 16'he4aa;
    SB_LUT4 n69002_bdd_4_lut (.I0(n69002), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n69005));
    defparam n69002_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1626 (.I0(\data_out_frame[11] [5]), .I1(n58475), 
            .I2(n58561), .I3(\data_out_frame[13] [6]), .O(n58641));
    defparam i1_2_lut_4_lut_adj_1626.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1627 (.I0(n53279), .I1(n21), .I2(n19), 
            .I3(n20), .O(n58377));
    defparam i1_2_lut_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5289));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1628 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(n53285), .I3(n25269), .O(n54224));
    defparam i2_3_lut_4_lut_adj_1628.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_776_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1629 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5288));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1629.LUT_INIT = 16'ha088;
    SB_LUT4 i14067_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n29810));   // verilog/coms.v(148[4] 304[11])
    defparam i14067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14068_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n29811));   // verilog/coms.v(148[4] 304[11])
    defparam i14068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_adj_1630 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n58121), .O(n58146));
    defparam i1_2_lut_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n67569), .I2(n65591), .I3(byte_transmit_counter[4]), .O(n68996));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1631 (.I0(\data_in_frame[16]_c [0]), .I1(n14_adj_5605), 
            .I2(n10_adj_5638), .I3(\data_in_frame[13] [6]), .O(n23480));   // verilog/coms.v(88[17:63])
    defparam i7_4_lut_adj_1631.LUT_INIT = 16'h6996;
    SB_LUT4 n68996_bdd_4_lut (.I0(n68996), .I1(n68711), .I2(n68843), .I3(byte_transmit_counter[4]), 
            .O(tx_data[4]));
    defparam n68996_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14069_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n29812));   // verilog/coms.v(148[4] 304[11])
    defparam i14069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14070_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n29813));   // verilog/coms.v(148[4] 304[11])
    defparam i14070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14071_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n29814));   // verilog/coms.v(148[4] 304[11])
    defparam i14071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14072_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n29815));   // verilog/coms.v(148[4] 304[11])
    defparam i14072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14073_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n29816));   // verilog/coms.v(148[4] 304[11])
    defparam i14073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14074_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n29817));   // verilog/coms.v(148[4] 304[11])
    defparam i14074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14075_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n29818));   // verilog/coms.v(148[4] 304[11])
    defparam i14075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5543));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51782 (.I0(byte_transmit_counter[1]), 
            .I1(n62917), .I2(n62918), .I3(byte_transmit_counter[2]), .O(n68708));
    defparam byte_transmit_counter_1__bdd_4_lut_51782.LUT_INIT = 16'he4aa;
    SB_LUT4 i14076_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n29819));   // verilog/coms.v(148[4] 304[11])
    defparam i14076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14077_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n29820));   // verilog/coms.v(148[4] 304[11])
    defparam i14077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5287));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1632 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_5639));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1632.LUT_INIT = 16'h7bde;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51911 (.I0(byte_transmit_counter[3]), 
            .I1(n67535), .I2(n65559), .I3(byte_transmit_counter[4]), .O(n68984));
    defparam byte_transmit_counter_3__bdd_4_lut_51911.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut_adj_1633 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_5640));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1633.LUT_INIT = 16'h7bde;
    SB_LUT4 i14078_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n29821));   // verilog/coms.v(148[4] 304[11])
    defparam i14078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14079_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n29822));   // verilog/coms.v(148[4] 304[11])
    defparam i14079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14080_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n29823));   // verilog/coms.v(148[4] 304[11])
    defparam i14080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_4_lut_adj_1634 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n2092), .I3(n2095), .O(n25090));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1634.LUT_INIT = 16'h4000;
    SB_LUT4 i2_3_lut_4_lut_adj_1635 (.I0(n2092), .I1(n4452), .I2(n2095), 
            .I3(n2098), .O(n60003));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1635.LUT_INIT = 16'h2000;
    SB_LUT4 i14081_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n29824));   // verilog/coms.v(148[4] 304[11])
    defparam i14081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14082_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n29825));   // verilog/coms.v(148[4] 304[11])
    defparam i14082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_4_lut_4_lut (.I0(n2092), .I1(n4452), .I2(n62488), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n60217));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 n68984_bdd_4_lut (.I0(n68984), .I1(n68681), .I2(n7_adj_5641), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n68984_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1636 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n58288), .I3(\data_out_frame[20] [5]), .O(n2217));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1636.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1637 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [1]), .I3(\data_out_frame[20] [2]), 
            .O(n58288));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1637.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5314));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_776_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14083_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n29826));   // verilog/coms.v(148[4] 304[11])
    defparam i14083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_776_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5286));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1638 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[17] [6]), .I3(GND_net), .O(n58733));
    defparam i1_2_lut_3_lut_adj_1638.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1639 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[12] [4]), .I3(\data_out_frame[12] [6]), 
            .O(n6_adj_5556));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1640 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[18] [3]), .I3(GND_net), .O(n58848));
    defparam i1_2_lut_3_lut_adj_1640.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1641 (.I0(\data_in_frame[2]_c [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n26225));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1642 (.I0(n58207), .I1(\data_out_frame[16] [6]), 
            .I2(n58151), .I3(n54253), .O(n54243));
    defparam i1_2_lut_4_lut_adj_1642.LUT_INIT = 16'h9669;
    SB_LUT4 n68708_bdd_4_lut (.I0(n68708), .I1(n62867), .I2(n62866), .I3(byte_transmit_counter[2]), 
            .O(n68711));
    defparam n68708_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14084_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n29827));   // verilog/coms.v(148[4] 304[11])
    defparam i14084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1643 (.I0(\data_out_frame[21] [6]), .I1(\data_out_frame[21] [7]), 
            .I2(n26288), .I3(GND_net), .O(n58819));
    defparam i1_2_lut_3_lut_adj_1643.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1644 (.I0(reset), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [0]), .O(n58108));
    defparam i1_2_lut_4_lut_adj_1644.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1645 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[22] [6]), .I3(GND_net), .O(n58903));
    defparam i1_2_lut_3_lut_adj_1645.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1646 (.I0(n58794), .I1(n58906), .I2(\data_out_frame[20] [6]), 
            .I3(\data_out_frame[20] [7]), .O(n58940));
    defparam i2_3_lut_4_lut_adj_1646.LUT_INIT = 16'h6996;
    SB_LUT4 i12226_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5617), 
            .I2(n58133), .I3(reset), .O(n27968));   // verilog/coms.v(157[7:23])
    defparam i12226_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i5_3_lut_4_lut_adj_1647 (.I0(n53247), .I1(n10_adj_5542), .I2(n25814), 
            .I3(n58511), .O(n53191));
    defparam i5_3_lut_4_lut_adj_1647.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1648 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5617), 
            .I2(n58121), .I3(n10_adj_5642), .O(n58143));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1648.LUT_INIT = 16'hfffd;
    SB_LUT4 i14085_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n29828));   // verilog/coms.v(148[4] 304[11])
    defparam i14085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14086_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n29829));   // verilog/coms.v(148[4] 304[11])
    defparam i14086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14087_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n29830));   // verilog/coms.v(148[4] 304[11])
    defparam i14087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14088_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n29831));   // verilog/coms.v(148[4] 304[11])
    defparam i14088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14089_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n29832));   // verilog/coms.v(148[4] 304[11])
    defparam i14089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1649 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8][3] ), .I3(n25301), .O(n58919));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1649.LUT_INIT = 16'h6996;
    SB_LUT4 select_776_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1650 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n58258));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1650.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1651 (.I0(\data_in_frame[6] [7]), .I1(n25370), 
            .I2(n58701), .I3(\data_in_frame[4] [5]), .O(n25859));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1651.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1652 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [6]), .I3(n25666), .O(n26330));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1652.LUT_INIT = 16'h6996;
    SB_LUT4 i14091_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n29834));   // verilog/coms.v(148[4] 304[11])
    defparam i14091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1653 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n58632));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1653.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [3]), 
            .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5285));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'ha088;
    SB_LUT4 select_776_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_4_lut_adj_1655 (.I0(n53191), .I1(\data_out_frame[23] [3]), 
            .I2(n25947), .I3(n53925), .O(n6_adj_5518));
    defparam i2_2_lut_4_lut_adj_1655.LUT_INIT = 16'h9669;
    SB_LUT4 select_776_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5309));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51901 (.I0(byte_transmit_counter[3]), 
            .I1(n67533), .I2(n65546), .I3(byte_transmit_counter[4]), .O(n68978));
    defparam byte_transmit_counter_3__bdd_4_lut_51901.LUT_INIT = 16'he4aa;
    SB_LUT4 i14092_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n29835));   // verilog/coms.v(148[4] 304[11])
    defparam i14092_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1656 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n25656), .I3(n58276), .O(n1312));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1656.LUT_INIT = 16'h6996;
    SB_LUT4 n68978_bdd_4_lut (.I0(n68978), .I1(n68669), .I2(n7_adj_5643), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n68978_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51692 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n68696));
    defparam byte_transmit_counter_0__bdd_4_lut_51692.LUT_INIT = 16'he4aa;
    SB_LUT4 i14093_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n29836));   // verilog/coms.v(148[4] 304[11])
    defparam i14093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1657 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[8][5] ), .I3(GND_net), .O(n58343));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1657.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1658 (.I0(\data_out_frame[11] [5]), .I1(n58475), 
            .I2(n58707), .I3(n58370), .O(n53666));
    defparam i2_3_lut_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1659 (.I0(\data_out_frame[11] [5]), .I1(n58475), 
            .I2(n58561), .I3(GND_net), .O(n58562));
    defparam i1_2_lut_3_lut_adj_1659.LUT_INIT = 16'h9696;
    SB_LUT4 i14094_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n29837));   // verilog/coms.v(148[4] 304[11])
    defparam i14094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1660 (.I0(n58197), .I1(n58626), .I2(n25763), 
            .I3(\data_out_frame[4] [7]), .O(n24827));   // verilog/coms.v(74[16:62])
    defparam i2_3_lut_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 i14095_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n29838));   // verilog/coms.v(148[4] 304[11])
    defparam i14095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13_2_lut_3_lut (.I0(n58197), .I1(n58626), .I2(\data_out_frame[5] [0]), 
            .I3(GND_net), .O(n25456));   // verilog/coms.v(74[16:62])
    defparam i13_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14096_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n29839));   // verilog/coms.v(148[4] 304[11])
    defparam i14096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i42094_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5617), 
            .I2(n58133), .I3(reset), .O(n7));   // verilog/coms.v(157[7:23])
    defparam i42094_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14097_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n29840));   // verilog/coms.v(148[4] 304[11])
    defparam i14097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n68696_bdd_4_lut (.I0(n68696), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n68699));
    defparam n68696_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14098_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n29841));   // verilog/coms.v(148[4] 304[11])
    defparam i14098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1661 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5617), 
            .I2(n58121), .I3(n10_adj_5642), .O(n58142));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1662 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(n25456), .I3(GND_net), .O(n25763));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1662.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1663 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[8][7] ), .I3(n58189), .O(n58704));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1663.LUT_INIT = 16'h6996;
    SB_LUT4 i14099_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n29842));   // verilog/coms.v(148[4] 304[11])
    defparam i14099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_2_lut_3_lut (.I0(n25269), .I1(n25830), .I2(n53283), .I3(GND_net), 
            .O(n16_adj_5573));   // verilog/coms.v(77[16:43])
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1664 (.I0(n25269), .I1(n25830), .I2(\data_out_frame[15] [4]), 
            .I3(GND_net), .O(n58502));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1664.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1665 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(n58468), .I3(\data_in_frame[13] [7]), .O(n10_adj_5638));
    defparam i2_2_lut_3_lut_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(\data_in_frame[18] [7]), 
            .I3(rx_data[7]), .O(n57448));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i13812_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n29555));
    defparam i13812_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13809_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n29552));
    defparam i13809_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1666 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_5644));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1666.LUT_INIT = 16'h7bde;
    SB_LUT4 i51345_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(\data_in_frame[18] [4]), 
            .I3(rx_data[4]), .O(n57436));
    defparam i51345_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i13803_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n29546));
    defparam i13803_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i51344_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(\data_in_frame[18] [2]), 
            .I3(rx_data[2]), .O(n57430));
    defparam i51344_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i11_4_lut_4_lut (.I0(reset), .I1(n27918), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n57450));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13794_3_lut_4_lut (.I0(reset), .I1(n27918), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n29537));
    defparam i13794_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14100_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n29843));   // verilog/coms.v(148[4] 304[11])
    defparam i14100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51896 (.I0(byte_transmit_counter[3]), 
            .I1(n67527), .I2(n65478), .I3(byte_transmit_counter[4]), .O(n68972));
    defparam byte_transmit_counter_3__bdd_4_lut_51896.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51662 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n68690));
    defparam byte_transmit_counter_0__bdd_4_lut_51662.LUT_INIT = 16'he4aa;
    SB_LUT4 i14101_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n29844));   // verilog/coms.v(148[4] 304[11])
    defparam i14101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14102_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n29845));   // verilog/coms.v(148[4] 304[11])
    defparam i14102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n68972_bdd_4_lut (.I0(n68972), .I1(n62994), .I2(n7_adj_5645), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n68972_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1667 (.I0(\data_out_frame[16] [4]), .I1(n53247), 
            .I2(n58736), .I3(\data_out_frame[18] [5]), .O(n25645));
    defparam i2_3_lut_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 i14103_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n29846));   // verilog/coms.v(148[4] 304[11])
    defparam i14103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1668 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5646));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5544), .I3(\FRAME_MATCHER.i_31__N_2512 ), .O(n26494));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'haaa8;
    SB_LUT4 i14104_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n29847));   // verilog/coms.v(148[4] 304[11])
    defparam i14104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1670 (.I0(n59852), .I1(n58794), .I2(n58906), 
            .I3(n25800), .O(n6_adj_5504));
    defparam i1_2_lut_4_lut_adj_1670.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1671 (.I0(n26225), .I1(n58359), .I2(\data_in_frame[7] [1]), 
            .I3(GND_net), .O(n58701));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1671.LUT_INIT = 16'h9696;
    SB_LUT4 i13844_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29587));
    defparam i13844_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1672 (.I0(n9_adj_5646), .I1(n11_adj_5644), .I2(n10_adj_5640), 
            .I3(n12_adj_5639), .O(n60269));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i13841_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29584));
    defparam i13841_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n68690_bdd_4_lut (.I0(n68690), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n68693));
    defparam n68690_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14105_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n29848));   // verilog/coms.v(148[4] 304[11])
    defparam i14105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_4_lut_4_lut_adj_1673 (.I0(n27916), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n57482));
    defparam i11_4_lut_4_lut_adj_1673.LUT_INIT = 16'hfe10;
    SB_LUT4 i13834_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29577));
    defparam i13834_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13827_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29570));
    defparam i13827_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13824_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29567));
    defparam i13824_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13821_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29564));
    defparam i13821_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14106_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16][7] ), 
            .I3(deadband[7]), .O(n29849));   // verilog/coms.v(148[4] 304[11])
    defparam i14106_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14107_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n29850));   // verilog/coms.v(148[4] 304[11])
    defparam i14107_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13818_3_lut_4_lut (.I0(n27916), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29561));
    defparam i13818_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14108_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16][5] ), 
            .I3(deadband[5]), .O(n29851));   // verilog/coms.v(148[4] 304[11])
    defparam i14108_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14109_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16][4] ), 
            .I3(deadband[4]), .O(n29852));   // verilog/coms.v(148[4] 304[11])
    defparam i14109_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1674 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_748), 
            .I2(n58337), .I3(\data_in_frame[2] [1]), .O(n23_adj_5647));
    defparam i6_4_lut_adj_1674.LUT_INIT = 16'h1248;
    SB_LUT4 i1_2_lut_3_lut_adj_1675 (.I0(Kp_23__N_974), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n25335));
    defparam i1_2_lut_3_lut_adj_1675.LUT_INIT = 16'h9696;
    SB_LUT4 i14110_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n29853));   // verilog/coms.v(148[4] 304[11])
    defparam i14110_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_3_lut (.I0(n25377), .I1(n25936), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n26_adj_5648));
    defparam i9_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i14111_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n29854));   // verilog/coms.v(148[4] 304[11])
    defparam i14111_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12_4_lut_adj_1676 (.I0(n23_adj_5647), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[2]_c [7]), .I3(n58179), .O(n29_c));
    defparam i12_4_lut_adj_1676.LUT_INIT = 16'h8008;
    SB_LUT4 i19906_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(deadband[1]), 
            .I3(\data_in_frame[16]_c [1]), .O(n29855));   // verilog/coms.v(148[4] 304[11])
    defparam i19906_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_adj_1677 (.I0(n25259), .I1(n58443), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n54146));
    defparam i1_2_lut_3_lut_adj_1677.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1678 (.I0(n25259), .I1(n58443), .I2(\data_out_frame[16] [3]), 
            .I3(\data_out_frame[14] [3]), .O(n58736));
    defparam i2_3_lut_4_lut_adj_1678.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1679 (.I0(Kp_23__N_878), .I1(\data_in_frame[6] [5]), 
            .I2(Kp_23__N_875), .I3(\data_in_frame[6] [4]), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1679.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1680 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5602), 
            .I2(n53), .I3(\FRAME_MATCHER.i [5]), .O(n27997));   // verilog/coms.v(157[7:23])
    defparam i2_3_lut_4_lut_adj_1680.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1681 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5602), 
            .I2(n58121), .I3(n10_adj_5642), .O(n58141));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1681.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_3_lut_4_lut (.I0(n25830), .I1(n58185), .I2(n58733), .I3(n2217), 
            .O(n20_adj_5575));   // verilog/coms.v(77[16:43])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13256_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][0] ), 
            .I3(\Kp[0] ), .O(n28999));   // verilog/coms.v(148[4] 304[11])
    defparam i13256_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13269_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[5][0] ), 
            .I3(\Ki[0] ), .O(n29012));   // verilog/coms.v(148[4] 304[11])
    defparam i13269_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1682 (.I0(n26330), .I1(n58623), .I2(\data_out_frame[19] [4]), 
            .I3(n53988), .O(n54293));
    defparam i2_3_lut_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1683 (.I0(n26330), .I1(n58623), .I2(\data_out_frame[19] [3]), 
            .I3(n58608), .O(n54324));
    defparam i2_3_lut_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 i13529_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n29272));
    defparam i13529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13532_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n29275));
    defparam i13532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13535_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n29278));
    defparam i13535_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13538_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n29281));
    defparam i13538_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13541_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n29284));
    defparam i13541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1684 (.I0(n26031), .I1(\data_in_frame[11] [6]), 
            .I2(n25549), .I3(GND_net), .O(n58468));
    defparam i1_2_lut_3_lut_adj_1684.LUT_INIT = 16'h9696;
    SB_LUT4 i13544_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n29287));
    defparam i13544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13276_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n29019));   // verilog/coms.v(148[4] 304[11])
    defparam i13276_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13547_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n29290));
    defparam i13547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13550_3_lut_4_lut (.I0(n39291), .I1(n58146), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29293));
    defparam i13550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13901_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29644));
    defparam i13901_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1685 (.I0(Kp_23__N_1748), .I1(n30_c), .I2(n32809), 
            .I3(GND_net), .O(n5_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1685.LUT_INIT = 16'hf8f8;
    SB_LUT4 mux_1045_i7_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[19] [6]), .O(n4793[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i14178_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29921));
    defparam i14178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14181_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29924));
    defparam i14181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1045_i8_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3]_c [7]), 
            .I3(\data_in_frame[19] [7]), .O(n4793[7]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i14184_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29927));
    defparam i14184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14187_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29930));
    defparam i14187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14190_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29933));
    defparam i14190_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14193_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29936));
    defparam i14193_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14196_3_lut_4_lut (.I0(n8_adj_5584), .I1(n58146), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29939));
    defparam i14196_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13484_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n29227));
    defparam i13484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13481_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n29224));
    defparam i13481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13488_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n29231));
    defparam i13488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13478_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n29221));
    defparam i13478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1045_i9_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[18] [0]), .O(n4793[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51672 (.I0(byte_transmit_counter[1]), 
            .I1(n62812), .I2(n62813), .I3(byte_transmit_counter[2]), .O(n68678));
    defparam byte_transmit_counter_1__bdd_4_lut_51672.LUT_INIT = 16'he4aa;
    SB_LUT4 i13517_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n29260));
    defparam i13517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1686 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(n58173), .I3(n58620), .O(n8_adj_5489));
    defparam i1_2_lut_4_lut_adj_1686.LUT_INIT = 16'h6996;
    SB_LUT4 i13520_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n29263));
    defparam i13520_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13523_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n29266));
    defparam i13523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i12_3_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\data_out_frame[15] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n12_adj_5541));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19803_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[18] [1]), .O(n4793[9]));   // verilog/coms.v(148[4] 304[11])
    defparam i19803_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i11_3_lut (.I0(\data_out_frame[12] [0]), 
            .I1(\data_out_frame[13] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n11_adj_5540));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1687 (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(n10_adj_5501), .I3(\data_in_frame[11] [2]), .O(n58297));
    defparam i1_2_lut_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1688 (.I0(n58173), .I1(n58620), .I2(n26031), 
            .I3(GND_net), .O(n26297));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1688.LUT_INIT = 16'h9696;
    SB_LUT4 i13526_3_lut_4_lut (.I0(n8_adj_5519), .I1(n58146), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n29269));
    defparam i13526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n68678_bdd_4_lut (.I0(n68678), .I1(n62858), .I2(n62857), .I3(byte_transmit_counter[2]), 
            .O(n68681));
    defparam n68678_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19444_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [2]), 
            .I3(\data_in_frame[18] [2]), .O(n4793[10]));   // verilog/coms.v(148[4] 304[11])
    defparam i19444_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1045_i12_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2][3] ), 
            .I3(\data_in_frame[18] [3]), .O(n4793[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_adj_1689 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[17] [5]), 
            .I2(n58185), .I3(GND_net), .O(n58647));
    defparam i1_2_lut_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1690 (.I0(\data_in_frame[5]_c [5]), .I1(n58534), 
            .I2(n25479), .I3(\data_in_frame[7] [6]), .O(n25569));
    defparam i2_3_lut_4_lut_adj_1690.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1691 (.I0(\data_in_frame[1] [5]), .I1(n58219), 
            .I2(\data_in_frame[6] [0]), .I3(\data_in_frame[3] [6]), .O(n26388));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_4_lut_adj_1691.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1692 (.I0(n25944), .I1(\data_in_frame[16] [6]), 
            .I2(n53130), .I3(GND_net), .O(n54274));
    defparam i1_2_lut_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1693 (.I0(\data_in_frame[18] [7]), .I1(n60010), 
            .I2(\data_in_frame[19] [1]), .I3(GND_net), .O(n54156));
    defparam i1_2_lut_3_lut_adj_1693.LUT_INIT = 16'h6969;
    SB_LUT4 i13655_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n29398));   // verilog/coms.v(148[4] 304[11])
    defparam i13655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1694 (.I0(\data_in_frame[14] [7]), .I1(n25437), 
            .I2(\data_in_frame[15] [0]), .I3(\data_in_frame[12] [6]), .O(n6_adj_5470));
    defparam i1_2_lut_4_lut_adj_1694.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1695 (.I0(\data_in_frame[16][7] ), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[9] [7]), .I3(n58551), .O(n58291));
    defparam i1_2_lut_4_lut_adj_1695.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1696 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[9] [7]), 
            .I2(n58551), .I3(GND_net), .O(n58400));
    defparam i1_2_lut_3_lut_adj_1696.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1697 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n26424));
    defparam i1_2_lut_3_lut_adj_1697.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1698 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(n60272), .I3(n60594), .O(n23344));
    defparam i2_3_lut_4_lut_adj_1698.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1699 (.I0(n53703), .I1(\data_in_frame[12] [4]), 
            .I2(n25604), .I3(\data_in_frame[12] [5]), .O(n54180));
    defparam i2_3_lut_4_lut_adj_1699.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1700 (.I0(\data_in_frame[8] [6]), .I1(n25549), 
            .I2(n25569), .I3(\data_in_frame[8] [7]), .O(n58864));   // verilog/coms.v(74[16:27])
    defparam i1_3_lut_4_lut_adj_1700.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1701 (.I0(n25830), .I1(n58185), .I2(\data_out_frame[17] [5]), 
            .I3(\data_out_frame[15] [4]), .O(n26288));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1701.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1045_i2_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3] [1]), 
            .I3(\data_in_frame[19] [1]), .O(n4793[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i2_3_lut_4_lut_adj_1702 (.I0(\data_in_frame[1] [5]), .I1(n58182), 
            .I2(\data_in_frame[8] [2]), .I3(\data_in_frame[8] [1]), .O(n58695));
    defparam i2_3_lut_4_lut_adj_1702.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1703 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_748), 
            .I2(\data_in_frame[1] [1]), .I3(n58300), .O(n22_adj_5649));
    defparam i5_4_lut_adj_1703.LUT_INIT = 16'h2184;
    SB_LUT4 i1_2_lut_3_lut_adj_1704 (.I0(\data_in_frame[14] [2]), .I1(n24758), 
            .I2(n25757), .I3(GND_net), .O(n58349));
    defparam i1_2_lut_3_lut_adj_1704.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1705 (.I0(LED_c), .I1(n32797), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5537));
    defparam i1_2_lut_adj_1705.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1706 (.I0(n53703), .I1(\data_in_frame[14] [4]), 
            .I2(n53398), .I3(n58825), .O(n25944));
    defparam i1_2_lut_4_lut_adj_1706.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1045_i3_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][2] ), 
            .I3(\data_in_frame[19] [2]), .O(n4793[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i17066_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n32809));   // verilog/coms.v(118[11:12])
    defparam i17066_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i2_3_lut_4_lut_adj_1707 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(n58677), .I3(n23480), .O(n53772));
    defparam i2_3_lut_4_lut_adj_1707.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1045_i4_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][3] ), 
            .I3(\data_in_frame[19] [3]), .O(n4793[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51647 (.I0(byte_transmit_counter[1]), 
            .I1(n62836), .I2(n62837), .I3(byte_transmit_counter[2]), .O(n68672));
    defparam byte_transmit_counter_1__bdd_4_lut_51647.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1708 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[19] [0]), 
            .I2(\data_in_frame[20]_c [7]), .I3(GND_net), .O(n6_adj_5434));
    defparam i1_2_lut_3_lut_adj_1708.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5305));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1709 (.I0(\data_in_frame[16][4] ), .I1(n58349), 
            .I2(n58854), .I3(\data_in_frame[16] [3]), .O(n58383));
    defparam i2_3_lut_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1710 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[14] [2]), 
            .I2(n24758), .I3(GND_net), .O(n6_adj_5433));
    defparam i1_2_lut_3_lut_adj_1710.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5304));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1711 (.I0(\data_in_frame[11] [5]), .I1(Kp_23__N_993), 
            .I2(n53463), .I3(GND_net), .O(n58810));
    defparam i1_2_lut_3_lut_adj_1711.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1045_i5_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][4] ), 
            .I3(\data_in_frame[19] [4]), .O(n4793[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i5_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_776_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5303));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_776_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5302));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1712 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n58346));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1712.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1713 (.I0(n26055), .I1(n25604), .I2(\data_in_frame[12] [5]), 
            .I3(GND_net), .O(n25596));
    defparam i1_2_lut_3_lut_adj_1713.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1045_i1_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3][0] ), 
            .I3(\data_in_frame[19] [0]), .O(n4793[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i19238_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[3]_c [5]), 
            .I3(\data_in_frame[19] [5]), .O(n4793[5]));   // verilog/coms.v(148[4] 304[11])
    defparam i19238_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_adj_1714 (.I0(n25859), .I1(n53463), .I2(\data_in_frame[9] [4]), 
            .I3(\data_in_frame[11] [5]), .O(n58588));
    defparam i1_2_lut_4_lut_adj_1714.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [6]), 
            .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'ha088;
    SB_LUT4 i15_4_lut_adj_1716 (.I0(n29_c), .I1(n25908), .I2(n26_adj_5648), 
            .I3(n26225), .O(n32));
    defparam i15_4_lut_adj_1716.LUT_INIT = 16'h0020;
    SB_LUT4 i19907_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[17]_c [7]), .O(n4793[23]));   // verilog/coms.v(148[4] 304[11])
    defparam i19907_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_1626_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5538));   // verilog/coms.v(148[4] 304[11])
    defparam select_1626_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1045_i23_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[17] [6]), .O(n4793[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1045_i22_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[17] [5]), .O(n4793[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1045_i21_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[17] [4]), .O(n4793[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_3_lut_4_lut_adj_1717 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(n58194), .I3(Kp_23__N_1080), .O(n53187));
    defparam i1_3_lut_4_lut_adj_1717.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1045_i20_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[17] [3]), .O(n4793[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 n68672_bdd_4_lut (.I0(n68672), .I1(n62852), .I2(n62851), .I3(byte_transmit_counter[2]), 
            .O(n68675));
    defparam n68672_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1045_i19_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [2]), 
            .I3(\data_in_frame[17] [2]), .O(n4793[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i19_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1045_i18_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[17] [1]), .O(n4793[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i18_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1045_i17_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[1] [0]), 
            .I3(\data_in_frame[17][0] ), .O(n4793[16]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i17_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i19383_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [7]), 
            .I3(\data_in_frame[18] [7]), .O(n4793[15]));   // verilog/coms.v(148[4] 304[11])
    defparam i19383_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_adj_1718 (.I0(n58724), .I1(n25511), .I2(n25859), 
            .I3(n25426), .O(n62150));
    defparam i1_2_lut_4_lut_adj_1718.LUT_INIT = 16'h6996;
    SB_LUT4 i19384_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [6]), 
            .I3(\data_in_frame[18] [6]), .O(n4793[14]));   // verilog/coms.v(148[4] 304[11])
    defparam i19384_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1045_i14_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2][5] ), 
            .I3(\data_in_frame[18] [5]), .O(n4793[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1045_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_adj_1719 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[21] [0]), .I3(GND_net), .O(n58906));
    defparam i1_2_lut_3_lut_adj_1719.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1720 (.I0(n59916), .I1(n54284), .I2(n54184), 
            .I3(\data_in_frame[17] [5]), .O(Kp_23__N_1551));
    defparam i1_2_lut_4_lut_adj_1720.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1721 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[18] [5]), .I3(n58440), .O(n53119));
    defparam i2_3_lut_4_lut_adj_1721.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1722 (.I0(\data_out_frame[18] [4]), .I1(n59852), 
            .I2(\data_out_frame[16] [1]), .I3(n58478), .O(n53169));
    defparam i2_3_lut_4_lut_adj_1722.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1723 (.I0(\data_out_frame[18] [4]), .I1(n59852), 
            .I2(\data_out_frame[22] [5]), .I3(GND_net), .O(n6_adj_5545));
    defparam i1_2_lut_3_lut_adj_1723.LUT_INIT = 16'h6969;
    SB_LUT4 i19445_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n30_c), .I2(\data_in_frame[2]_c [4]), 
            .I3(\data_in_frame[18] [4]), .O(n4793[12]));   // verilog/coms.v(148[4] 304[11])
    defparam i19445_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i11871_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3579), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n27612));   // verilog/coms.v(158[12:15])
    defparam i11871_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 select_778_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5546));
    defparam select_778_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1724 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n58092));
    defparam i1_2_lut_3_lut_adj_1724.LUT_INIT = 16'hfefe;
    SB_LUT4 select_778_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5418));
    defparam select_778_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i5_3_lut_4_lut_adj_1725 (.I0(\data_out_frame[13] [7]), .I1(n58585), 
            .I2(n54243), .I3(n60509), .O(n14_adj_5508));
    defparam i5_3_lut_4_lut_adj_1725.LUT_INIT = 16'h9669;
    SB_LUT4 select_778_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5416));
    defparam select_778_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_3_lut_4_lut_adj_1726 (.I0(\data_in_frame[15] [1]), .I1(n53096), 
            .I2(\data_in_frame[13] [7]), .I3(\data_in_frame[13] [6]), .O(n58816));
    defparam i1_3_lut_4_lut_adj_1726.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1727 (.I0(n54307), .I1(\data_out_frame[20] [4]), 
            .I2(n10_adj_5493), .I3(n58903), .O(n54235));
    defparam i5_3_lut_4_lut_adj_1727.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1728 (.I0(n53247), .I1(n58804), .I2(n10_adj_5568), 
            .I3(n58602), .O(n58412));
    defparam i5_3_lut_4_lut_adj_1728.LUT_INIT = 16'h6996;
    SB_LUT4 select_778_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5415));
    defparam select_778_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1729 (.I0(n53247), .I1(n58804), .I2(n54237), 
            .I3(GND_net), .O(n58961));
    defparam i1_2_lut_3_lut_adj_1729.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1730 (.I0(n53247), .I1(n58804), .I2(n25673), 
            .I3(n58478), .O(n53055));
    defparam i2_3_lut_4_lut_adj_1730.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut (.I0(n25426), .I1(Kp_23__N_974), .I2(\data_in_frame[8] [6]), 
            .I3(\data_in_frame[11] [0]), .O(n60197));   // verilog/coms.v(74[16:27])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 equal_313_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5578));   // verilog/coms.v(157[7:23])
    defparam equal_313_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_312_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5569));   // verilog/coms.v(157[7:23])
    defparam equal_312_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1731 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n53187), .I3(n25525), .O(n54148));
    defparam i1_3_lut_4_lut_adj_1731.LUT_INIT = 16'h9669;
    SB_LUT4 select_778_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n1_adj_5414));
    defparam select_778_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51642 (.I0(byte_transmit_counter[1]), 
            .I1(n62863), .I2(n62864), .I3(byte_transmit_counter[2]), .O(n68666));
    defparam byte_transmit_counter_1__bdd_4_lut_51642.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1732 (.I0(\data_in_frame[17] [1]), .I1(n58394), 
            .I2(\data_in_frame[19] [3]), .I3(n58520), .O(n23529));
    defparam i1_2_lut_4_lut_adj_1732.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1733 (.I0(\data_in_frame[17] [1]), .I1(n58394), 
            .I2(\data_in_frame[19] [3]), .I3(GND_net), .O(n58452));
    defparam i1_2_lut_3_lut_adj_1733.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_215_i3_3_lut_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(n23344), .I2(n58418), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5397));
    defparam select_776_Select_215_i3_3_lut_4_lut.LUT_INIT = 16'h6900;
    SB_LUT4 n68666_bdd_4_lut (.I0(n68666), .I1(n62846), .I2(n62845), .I3(byte_transmit_counter[2]), 
            .O(n68669));
    defparam n68666_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_776_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(n23344), .I2(n58306), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5394));
    defparam select_776_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h9600;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51637 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[25] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(\byte_transmit_counter[0] ), .O(n68660));
    defparam byte_transmit_counter_1__bdd_4_lut_51637.LUT_INIT = 16'he4aa;
    SB_LUT4 select_778_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n1_adj_5413));
    defparam select_778_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1734 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[23] [3]), .I3(n53191), .O(n6_adj_5458));
    defparam i2_2_lut_3_lut_4_lut_adj_1734.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_4_lut_adj_1735 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(n58605), .I3(\data_out_frame[25] [3]), .O(n8_adj_5552));
    defparam i3_3_lut_4_lut_adj_1735.LUT_INIT = 16'h6996;
    SB_LUT4 n68660_bdd_4_lut (.I0(n68660), .I1(\data_out_frame[26] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(\byte_transmit_counter[0] ), 
            .O(n68663));
    defparam n68660_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1736 (.I0(\data_in_frame[0] [5]), .I1(n58282), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[5][2] ), .O(n58270));
    defparam i2_3_lut_4_lut_adj_1736.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1737 (.I0(n10_adj_5642), .I1(n58121), .I2(n8_adj_5584), 
            .I3(GND_net), .O(n58140));
    defparam i1_2_lut_3_lut_adj_1737.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1738 (.I0(\data_in_frame[20][6] ), .I1(\data_in_frame[18] [3]), 
            .I2(n24742), .I3(GND_net), .O(n58727));
    defparam i1_2_lut_3_lut_adj_1738.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1739 (.I0(n10_adj_5642), .I1(n58121), .I2(n8_adj_5578), 
            .I3(GND_net), .O(n58144));
    defparam i1_2_lut_3_lut_adj_1739.LUT_INIT = 16'hfefe;
    SB_LUT4 select_778_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5412));
    defparam select_778_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1740 (.I0(n10_adj_5642), .I1(n58121), .I2(n8_adj_5519), 
            .I3(GND_net), .O(n58145));
    defparam i1_2_lut_3_lut_adj_1740.LUT_INIT = 16'hfefe;
    SB_LUT4 select_778_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_c));
    defparam select_778_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_4_lut_adj_1741 (.I0(Kp_23__N_1551), .I1(n53903), .I2(n25343), 
            .I3(\data_in_frame[17] [6]), .O(n6_adj_5393));
    defparam i1_2_lut_4_lut_adj_1741.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1742 (.I0(n10_adj_5642), .I1(n58121), .I2(n39291), 
            .I3(GND_net), .O(n58139));
    defparam i1_2_lut_3_lut_adj_1742.LUT_INIT = 16'hefef;
    SB_LUT4 equal_311_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5519));
    defparam equal_311_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i23643_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n39291));
    defparam i23643_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_4_lut_adj_1743 (.I0(n3579), .I1(n161), .I2(n10_adj_5642), 
            .I3(n58108), .O(n60939));
    defparam i2_3_lut_4_lut_adj_1743.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_adj_1744 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3579));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1744.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51632 (.I0(byte_transmit_counter[1]), 
            .I1(n63001), .I2(n63002), .I3(byte_transmit_counter[2]), .O(n68636));
    defparam byte_transmit_counter_1__bdd_4_lut_51632.LUT_INIT = 16'he4aa;
    SB_LUT4 n68636_bdd_4_lut (.I0(n68636), .I1(n63005), .I2(n63004), .I3(byte_transmit_counter[2]), 
            .O(n68639));
    defparam n68636_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1745 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n58092), .I3(LED_c), .O(n26862));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1745.LUT_INIT = 16'hfe00;
    SB_LUT4 equal_310_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_5642));   // verilog/coms.v(158[12:15])
    defparam equal_310_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_318_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_5530));   // verilog/coms.v(158[12:15])
    defparam equal_318_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n62901), .I3(n62899), .O(n7_adj_5645));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n62904), .I3(n62902), .O(n7_adj_5643));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n62889), .I3(n62887), .O(n7_adj_5641));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51619 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n68630));
    defparam byte_transmit_counter_0__bdd_4_lut_51619.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n62895), .I3(n62893), .O(n7_adj_8));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n62874), .I3(n62872), .O(n7_adj_9));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n62877), .I3(n62875), .O(n7_adj_10));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13895_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29638));
    defparam i13895_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13890_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29633));
    defparam i13890_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_776_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13887_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29630));
    defparam i13887_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_3_lut_4_lut_adj_1746 (.I0(n38022), .I1(n58108), .I2(\data_in_frame[21] [4]), 
            .I3(rx_data[4]), .O(n57414));
    defparam i11_3_lut_4_lut_adj_1746.LUT_INIT = 16'hf1e0;
    SB_LUT4 i41_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(\data_in_frame[21]_c [3]), 
            .I3(rx_data[3]), .O(n33_adj_5570));
    defparam i41_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i18134_3_lut (.I0(\current[0] ), .I1(n1828), .I2(n209), .I3(GND_net), 
            .O(n270));
    defparam i18134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n68630_bdd_4_lut (.I0(n68630), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n68633));
    defparam n68630_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13877_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29620));
    defparam i13877_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13874_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29617));
    defparam i13874_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13871_3_lut_4_lut (.I0(n38022), .I1(n58108), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29614));
    defparam i13871_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1747 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n58363));
    defparam i1_2_lut_3_lut_adj_1747.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1748 (.I0(\data_in_frame[5]_c [7]), .I1(\data_in_frame[5][6] ), 
            .I2(n25479), .I3(\data_in_frame[1] [4]), .O(n58219));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_4_lut_adj_1748.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1749 (.I0(\data_in_frame[9] [2]), .I1(n25871), 
            .I2(n26031), .I3(n58759), .O(n58571));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1749.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51610 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n68612));
    defparam byte_transmit_counter_0__bdd_4_lut_51610.LUT_INIT = 16'he4aa;
    SB_LUT4 n68612_bdd_4_lut (.I0(n68612), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n68615));
    defparam n68612_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1750 (.I0(n25908), .I1(n25377), .I2(\data_in_frame[6] [4]), 
            .I3(GND_net), .O(n58698));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1750.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1751 (.I0(\data_in_frame[2][3] ), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n25908));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1751.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1752 (.I0(n25908), .I1(n25377), .I2(\data_in_frame[5][0] ), 
            .I3(\data_in_frame[4] [7]), .O(n58359));   // verilog/coms.v(78[16:43])
    defparam i1_3_lut_4_lut_adj_1752.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1753 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(n58864), .I3(GND_net), .O(n6_adj_5447));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1753.LUT_INIT = 16'h9696;
    SB_LUT4 i13934_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29677));
    defparam i13934_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1754 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n25405));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1754.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1755 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(n58614), .I3(\data_in_frame[1] [0]), .O(n25448));   // verilog/coms.v(88[17:63])
    defparam i1_3_lut_4_lut_adj_1755.LUT_INIT = 16'h6996;
    SB_LUT4 i13931_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29674));
    defparam i13931_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1756 (.I0(n25405), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n58614));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1756.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1757 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2]_c [4]), .I3(GND_net), .O(n25377));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1757.LUT_INIT = 16'h9696;
    SB_LUT4 select_776_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1758 (.I0(\data_in_frame[9] [2]), .I1(n25871), 
            .I2(n26031), .I3(n58200), .O(n25544));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1758.LUT_INIT = 16'h6996;
    SB_LUT4 i13928_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29671));
    defparam i13928_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1759 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(n25936), .I3(GND_net), .O(n6_c));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1759.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1760 (.I0(n60269), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[1] [2]), .O(n27_adj_5653));
    defparam i10_4_lut_adj_1760.LUT_INIT = 16'h4000;
    SB_LUT4 i16_4_lut_adj_1761 (.I0(n27_adj_5653), .I1(n32), .I2(n62621), 
            .I3(n22_adj_5649), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1761.LUT_INIT = 16'h0800;
    SB_LUT4 select_776_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1762 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(n58674), .I3(\data_in_frame[4] [4]), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut_adj_1762.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_4_lut_adj_1763 (.I0(n27926), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n57420));
    defparam i11_4_lut_4_lut_adj_1763.LUT_INIT = 16'hfe10;
    SB_LUT4 i13915_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29658));
    defparam i13915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13912_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n29655));
    defparam i13912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13905_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29648));
    defparam i13905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1764 (.I0(n25405), .I1(n58285), .I2(Kp_23__N_875), 
            .I3(GND_net), .O(n6_adj_5299));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1764.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1765 (.I0(\data_in_frame[3][3] ), .I1(n10_c), 
            .I2(n25405), .I3(n58162), .O(n53770));
    defparam i5_3_lut_4_lut_adj_1765.LUT_INIT = 16'h6996;
    SB_LUT4 i13898_3_lut_4_lut (.I0(n27926), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n29641));
    defparam i13898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_776_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_776_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1766 (.I0(\data_in_frame[2][5] ), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n25370));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1766.LUT_INIT = 16'h9696;
    uart_tx tx (.GND_net(GND_net), .r_Clock_Count({r_Clock_Count}), .VCC_net(VCC_net), 
            .n1(n1), .tx_o(tx_o), .clk16MHz(clk16MHz), .tx_data({tx_data[7], 
            \tx_data[6] , tx_data[5:4], \tx_data[3] , \tx_data[2] , 
            \tx_data[1] , tx_data[0]}), .r_SM_Main({r_SM_Main}), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .n57758(n57758), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n61290(n61290), .n27(n27), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
            .n58968(n58968), .n29040(n29040), .tx_active(tx_active), .n69042(n69042), 
            .n29653(n29653), .n27295(n27295), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .n4894(n4894), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n29(n29), .n23(n23), .n59805(n59805), .n61278(n61278), 
            .n6(n6), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.baudrate({baudrate}), .GND_net(GND_net), .VCC_net(VCC_net), 
            .r_Clock_Count({r_Clock_Count_adj_22}), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n25117(n25117), .n29(n29), .n23(n23), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .clk16MHz(clk16MHz), 
            .\r_SM_Main[2] (\r_SM_Main[2]_adj_19 ), .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), 
            .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n4894(n4894), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
            .n57758(n57758), .n61290(n61290), .n4891(n4891), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_20 ), 
            .\r_SM_Main[1] (\r_SM_Main[1]_adj_21 ), .n58022(n58022), .n27288(n27288), 
            .n58970(n58970), .n61676(n61676), .n61604(n61604), .n61658(n61658), 
            .n61640(n61640), .n61586(n61586), .n61622(n61622), .n61550(n61550), 
            .n29912(n29912), .rx_data({rx_data}), .n29911(n29911), .n29910(n29910), 
            .n29909(n29909), .n29908(n29908), .n29907(n29907), .n29906(n29906), 
            .n29663(n29663), .n54370(n54370), .rx_data_ready(rx_data_ready), 
            .n29667(n29667), .n27292(n27292), .n61568(n61568), .\r_SM_Main[0] (r_SM_Main[0]), 
            .n59805(n59805), .n61280(n61280)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (GND_net, r_Clock_Count, VCC_net, n1, tx_o, clk16MHz, 
            tx_data, r_SM_Main, \r_Bit_Index[0] , n57758, \r_SM_Main_2__N_3545[0] , 
            n61290, n27, \r_SM_Main_2__N_3536[1] , n58968, n29040, 
            tx_active, n69042, n29653, n27295, \o_Rx_DV_N_3488[12] , 
            n4894, \o_Rx_DV_N_3488[24] , n29, n23, n59805, n61278, 
            n6, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [8:0]r_Clock_Count;
    input VCC_net;
    output n1;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    output \r_Bit_Index[0] ;
    output n57758;
    input \r_SM_Main_2__N_3545[0] ;
    input n61290;
    input n27;
    input \r_SM_Main_2__N_3536[1] ;
    output n58968;
    input n29040;
    output tx_active;
    input n69042;
    input n29653;
    output n27295;
    input \o_Rx_DV_N_3488[12] ;
    input n4894;
    input \o_Rx_DV_N_3488[24] ;
    input n29;
    input n23;
    input n59805;
    output n61278;
    output n6;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    
    wire n52182, n52181, n52180, n52179, n52178, n52177, n52176, 
        n52175, n3, n22384;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n21376;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n21375, n3_adj_5282, n59102, o_Tx_Serial_N_3598, n28715, 
        n62764, n62765, n62783, n62782;
    wire [2:0]n460;
    
    wire n28643, n61258, n61264, n65529, n65526, n68648;
    
    SB_LUT4 r_Clock_Count_1946_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n52182), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1946_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n52181), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_9 (.CI(n52181), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n52182));
    SB_LUT4 r_Clock_Count_1946_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n52180), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_8 (.CI(n52180), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n52181));
    SB_LUT4 r_Clock_Count_1946_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n52179), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_7 (.CI(n52179), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n52180));
    SB_LUT4 r_Clock_Count_1946_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n52178), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_6 (.CI(n52178), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n52179));
    SB_LUT4 r_Clock_Count_1946_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n52177), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_5 (.CI(n52177), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n52178));
    SB_LUT4 r_Clock_Count_1946_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n52176), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_4 (.CI(n52176), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n52177));
    SB_LUT4 r_Clock_Count_1946_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n52175), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_3 (.CI(n52175), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n52176));
    SB_LUT4 r_Clock_Count_1946_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1946_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1946_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n52175));
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n21376), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n57758));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i5952_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n61290), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n21375));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i5952_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i5953_3_lut (.I0(n21375), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21376));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i5953_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5282), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n22384), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i42134_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n59102));
    defparam i42134_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3598), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_1946__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_LUT4 i42008_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n58968));
    defparam i42008_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR r_Clock_Count_1946__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1946__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n28715));   // verilog/uart_tx.v(119[34:51])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29040));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i45748_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n62764));
    defparam i45748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45749_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n62765));
    defparam i45749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45767_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n62783));
    defparam i45767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45766_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n62782));
    defparam i45766_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n69042));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29653));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27295), 
            .D(n460[1]), .R(n28643));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27295), 
            .D(n460[2]), .R(n28643));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2176_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(99[36:51])
    defparam i2176_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_3_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4894), .I2(n57758), 
            .I3(GND_net), .O(n61258));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), .I3(n61258), 
            .O(n61264));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1108 (.I0(n61264), .I1(n59102), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n28643));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_4_lut_adj_1108.LUT_INIT = 16'h0323;
    SB_LUT4 i2169_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(99[36:51])
    defparam i2169_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51526_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3536[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n28715));
    defparam i51526_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i49259_3_lut (.I0(n4894), .I1(\o_Rx_DV_N_3488[12] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n65529));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i49259_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i49255_4_lut (.I0(n65529), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65526));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i49255_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n65526), .I1(n59805), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5282));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_3_lut_4_lut (.I0(n57758), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n61278));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i51586_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n27295));
    defparam i51586_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n59805), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n22384));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n62782), 
            .I2(n62783), .I3(r_Bit_Index[2]), .O(n68648));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n68648_bdd_4_lut (.I0(n68648), .I1(n62765), .I2(n62764), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3598));
    defparam n68648_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (baudrate, GND_net, VCC_net, r_Clock_Count, \o_Rx_DV_N_3488[24] , 
            n27, n25117, n29, n23, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[8] , 
            clk16MHz, \r_SM_Main[2] , \o_Rx_DV_N_3488[7] , r_Rx_Data, 
            RX_N_2, \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , 
            \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , 
            \o_Rx_DV_N_3488[0] , n4894, \r_SM_Main_2__N_3536[1] , n57758, 
            n61290, n4891, \r_Bit_Index[0] , \r_SM_Main[1] , n58022, 
            n27288, n58970, n61676, n61604, n61658, n61640, n61586, 
            n61622, n61550, n29912, rx_data, n29911, n29910, n29909, 
            n29908, n29907, n29906, n29663, n54370, rx_data_ready, 
            n29667, n27292, n61568, \r_SM_Main[0] , n59805, n61280) /* synthesis syn_module_defined=1 */ ;
    input [31:0]baudrate;
    input GND_net;
    input VCC_net;
    output [7:0]r_Clock_Count;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    output n25117;
    output n29;
    output n23;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[8] ;
    input clk16MHz;
    output \r_SM_Main[2] ;
    output \o_Rx_DV_N_3488[7] ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    input n4894;
    output \r_SM_Main_2__N_3536[1] ;
    input n57758;
    output n61290;
    input n4891;
    output \r_Bit_Index[0] ;
    output \r_SM_Main[1] ;
    input n58022;
    output n27288;
    output n58970;
    output n61676;
    output n61604;
    output n61658;
    output n61640;
    output n61586;
    output n61622;
    output n61550;
    input n29912;
    output [7:0]rx_data;
    input n29911;
    input n29910;
    input n29909;
    input n29908;
    input n29907;
    input n29906;
    input n29663;
    input n54370;
    output rx_data_ready;
    input n29667;
    output n27292;
    output n61568;
    input \r_SM_Main[0] ;
    output n59805;
    output n61280;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n67986, n67356, n45, n66623, n67358, n2715, n43, n2720, 
        n33, n2719, n35, n2723, n27_c, n1557;
    wire [23:0]n7651;
    wire [23:0]n294;
    
    wire n1698;
    wire [23:0]n7677;
    
    wire n1836;
    wire [23:0]n7885;
    
    wire n2713, n2977, n51750, n2722, n29_c, n2714, n2867, n51749, 
        n2721, n31, n2728, n17, n2727, n19, n2754, n51748, n2716, 
        n2638, n51747, n2717, n2519, n51746, n2718, n2397, n51745, 
        n2272, n51744, n2144, n51743, n2013, n51742, n1879, n51741, 
        n2726, n21, n1742, n51740, n2724, n1602, n51739, n2725, 
        n23_c, n1459, n51738, n1460, n51737, n1011, n51736, n856, 
        n51735, n25, n2729, n698, n51734, n2730, n858, n51733, 
        n61172, n538, n59295, n37;
    wire [23:0]n7859;
    
    wire n2596, n51717, n2597, n51716, n2598, n51715, n2599, n51714, 
        n2600, n51713, n2601, n51712, n2602, n51711, n2603, n51710, 
        n2604, n51709, n2605, n51708, n2606, n51707, n2607, n51706, 
        n2608, n51705, n2609, n51704, n2610, n51703, n2611, n51702, 
        n2612, n51701, n65669, n61170, n59299, n66579, n67314, 
        n67312, n37_adj_5006, n1554, n1695, n1833, n65672, n61166, 
        n48, n2491;
    wire [23:0]n7833;
    
    wire n14, n67803, n39, n67804, n22, n45_adj_5007, n40, n41, 
        n65665, n20, n65659, n67361, n67716, n62002, n61148, n61146, 
        n61992, n25206, n18, n26, n16, n65690, n68191;
    wire [7:0]n1;
    
    wire n52174, n52173, n52172, n52171, n52170, n52169, n43_adj_5012, 
        n52168, n68192, n68013, n2476, n51666, n67631, n2477, 
        n51665, n2478, n51664, n2479, n51663, n2480, n51662, n67991, 
        n2481, n51661, n2482, n51660, n67990, n1559, n1700, n2483, 
        n51659, n2484, n51658, n2485, n51657, n2486, n51656, n2487, 
        n51655, n17_adj_5014, n2488, n51654, n2489, n51653, n2490, 
        n51652, n23_adj_5015, n21_adj_5016, n19_adj_5017, n65741, 
        n51651, n61168, n59303, n67993, n51278, n1558, n1699, 
        n51277, n61066, n62747, n51276, n61210, n51275;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n51274, n61208;
    wire [23:0]n7807;
    
    wire n2353, n51632, n2354, n51631, n51273, n61206, n1837, 
        n2355, n51630, n51272, n2356, n51629, n29_adj_5021, n27_adj_5022, 
        n25_adj_5023, n65732, n51271, n61204, n35_adj_5024, n33_adj_5025, 
        n31_adj_5026, n67646, n2357, n51628, n1560, n1701, n51270, 
        n61202, n1839, n2358, n51627, n51269, n61064, n1838, n16_adj_5027, 
        n2359, n51626, n2360, n51625, n2361, n51624, n2362, n51623, 
        n2363, n51622, n31_adj_5028, n39_adj_5029, n67809, n51268, 
        n61200, n2364, n51621, n2365, n51620, n2366, n51619, n51267, 
        n41_adj_5030, n67810, n51266, n2367, n51618, n59307, n51265, 
        n51264, n51263, n51262, n65737, n66585, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n51261, r_Rx_Data_R, n22_adj_5031, n67359, n51260, n43_adj_5032, 
        n67709, n33_adj_5033, n1265, n38_adj_5034, n1266, n66017, 
        n51259, n51258;
    wire [23:0]n7781;
    
    wire n2227, n51601, n51257, n2228, n51600, n20_adj_5035, n28, 
        n2229, n51599, n2230, n51598, n51256, n2231, n51597, n18_adj_5036, 
        n65729, n68189, n51255, n2232, n51596, n2233, n51595, 
        n60086, n68190, n35_adj_5037, n2234, n51594, n68015, n37_adj_5038, 
        n66589, n67807, n67988, n2235, n51593, n68201, n2236, 
        n51592, n1555, n1696, n68202, n2237, n51591, n2238, n51590, 
        n1834, n41_adj_5039, n2239, n51589, n1414;
    wire [23:0]n7625;
    
    wire n1408, n1552, n1410, n43_adj_5040, n61126, n1409, n1553, 
        n1413, n37_adj_5041, n2240, n51588, n61164, n59311, n1411, 
        n41_adj_5042, n61284;
    wire [23:0]n7755;
    
    wire n2098, n51577, n1412, n1556, n39_adj_5043, n2099, n51576, 
        n2100, n51575, n61160, n48_adj_5044, n1261;
    wire [23:0]n7599;
    
    wire n1111;
    wire [23:0]n7573;
    
    wire n1264, n41_adj_5045, n1267, n36, n61884, n40_adj_5046, 
        n3_adj_5047, n68181, n61888, n5, n61892, n1263, n68182, 
        n8, n57790, n61104, n1262, n68039;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n48_adj_5048, n1112;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n57762, n45_adj_5049, n39001, n61296, n61302, n62625, n62723, 
        n2, n9679, n961, n962, n21487, n2101, n51574, n2102, 
        n51573, n2103, n51572, n804, n42_adj_5050, n960, n62673, 
        n2104, n51571, n3_adj_5051, n2105, n51570, n2106, n51569, 
        n2107, n51568, n42_adj_5052, n1113, n27409, n28713, n2108, 
        n51567, n2109, n51566, n2110, n65437, n65434;
    wire [23:0]n7729;
    
    wire n1966, n51556, n1967, n51555, n1968, n51554, n1969, n51553, 
        n1970, n51552, n43_adj_5053, n1971, n51551, n61964, n1972, 
        n51550, n20_adj_5054, n65789, n2843, n14_adj_5055, n2838, 
        n2842, n65643, n16_adj_5056, n2840, n18_adj_5057, n22_adj_5058, 
        n2830, n2839, n65625, n20_adj_5059, n68260, n25194, n1973, 
        n51549, n24, n1115, n18_adj_5060, n39_adj_5061, n1974, n51548, 
        n24_adj_5062, n1975, n51547, n65882, n26_adj_5063, n65893, 
        n65795, n28_adj_5064, n62711, n48_adj_5065, n2955, n12, 
        n2950, n2954, n65594, n14_adj_5066, n1976, n51546, n2952, 
        n16_adj_5067, n1977, n51545, n2942, n2951, n66456, n18_adj_5068;
    wire [23:0]n7703;
    
    wire n1831, n51544, n22_adj_5069, n14_adj_5070, n1832, n51543, 
        n15, n69043, n65847, n51542, n24_adj_5071, n48_adj_5072, 
        n20_adj_5073, n65854, n4, n6, n61664, n61670, n26_adj_5074, 
        n3064, n10, n61592, n61598, n51541, n1835, n51540, n3061, 
        n14_adj_5075, n25163, n65779, n48_adj_5076, n3051, n3060, 
        n66346, n51539, n16_adj_5077, n3059, n12_adj_5078, n3063, 
        n66402, n51538, n51537, n51536, n1840, n51535, n1841, 
        n51534, n61162, n59320, n805, n42_adj_5079, n1693, n51533, 
        n61646, n61652, n1694, n51532, n51531, n67785, n51530, 
        n803, n67786, n58994, n61988, n68155, n3151, n25221, n1697, 
        n51529, n61628, n61634, n61942, n51528, n61994, n51527, 
        n61872, n61946, n25212, n39003, n28_adj_5080, n65904, n30, 
        n3170, n8_adj_5081, n65498, n68388, n46, n3167, n12_adj_5082, 
        n61574, n61580, n58992, n48_adj_5083, n3157, n3166, n66243, 
        n61844, n61908, n61910, n61906, n61856, n14_adj_5084, n3165, 
        n10_adj_5085, n61848, n62004, n25166, n3169, n66298, n40_adj_5086, 
        n62106, n1114, n41_adj_5087, n21489, n9470, n44_adj_5088, 
        n959, n62498, n61710, n61712, n62500, n61714, n61092, 
        n62683, n62593, n60160, n61442, n61460, n62597, n62739, 
        n62719, n59034, n59802, n61990, n61610, n61616, n21473, 
        n21475, n68262, n62659, n61926, n43_adj_5089, n62655, n61936, 
        n61948, n61538, n61544, n62689, n61730, n61750, n25209, 
        n48_adj_5090, n26_adj_5091, n61706, n61702, n61704, n61724, 
        n51526, n61708, n61726, n51525, n1702, n51524, n51523, 
        n51522, n51521, n28_adj_5092, n51520, n51519, n51518, n51517, 
        n51516, n65931, n30_adj_5093, n51507, n51506, n51505, n51504, 
        n51503, n30_adj_5094, n51502, n65952, n51501, n1415, n51500, 
        n32, n59329, n51499, n61916, n61996, n61790;
    wire [2:0]n479;
    
    wire n28645, n67768, n25185, n32_adj_5095, n51498, n51497, n51496, 
        n51495, n51494, n65420, n59291, n51493, n61158, n59333, 
        n51492, n51491, n51490, n51489, n61918, n65421, n62516, 
        n51488, n1116, n51487, n61156, n59337, n62713, n59287;
    wire [23:0]n7989;
    
    wire n3186, n51892, n3152, n3082, n51891, n3153, n3188, n51890, 
        n3154, n3084, n51889, n25218, n59283, n3155, n51888, n3156, 
        n51887, n51886, n3158, n51885, n3159, n51884, n3160, n51883, 
        n3161, n51882, n3162, n51881, n3163, n51880, n3164, n51879, 
        n51878, n51877, n61904, n51876, n3168, n51875, n51874, 
        n51873, n3171, n51872, n3172, n51871, n61180, n51870, 
        n59279;
    wire [23:0]n7963;
    
    wire n3046, n51851, n3047, n51850, n3048, n51849, n3049, n51848, 
        n3050, n51847, n51846, n3052, n51845, n3053, n51844, n3054, 
        n51843, n3055, n51842, n3056, n51841, n3057, n51840, n3058, 
        n51839, n51838, n51837, n51836, n3062, n51835, n51834, 
        n51833, n3065, n51832, n3066, n51831, n61178;
    wire [23:0]n7937;
    
    wire n2938, n51830, n2939, n51829, n2940, n51828, n2941, n51827, 
        n51826, n2943, n51825, n2944, n51824, n2945, n51823, n2946, 
        n51822, n2947, n51821, n2948, n51820, n2949, n51819, n51818, 
        n51817, n51816, n2953, n51815, n51814, n51813, n2956, 
        n51812, n2957, n51811, n61176, n62609;
    wire [23:0]n7911;
    
    wire n2827, n51785, n2828, n51784, n2829, n51783, n51782, 
        n2831, n51781, n2832, n51780, n2833, n51779, n2834, n51778, 
        n2835, n51777, n2836, n51776, n2837, n51775, n51774, n51773, 
        n51772, n2841, n51771, n51770, n51769, n2844, n51768, 
        n2845, n51767, n61174, n61270, n61276, n61498, n62667, 
        n62100, n61526, n61556, n61562, n62737, n34, n65777, n44_adj_5096, 
        n9463, n9299, n44_adj_5097, n48_adj_5098, n25172, n46_adj_5099, 
        n58996, n46_adj_5100, n61976, n62102, n65409, n59340, n65406, 
        n42_adj_5101, n65403, n67781, n61234, n67782, n61240, n38_adj_5102, 
        n40_adj_5103, n42_adj_5104, n66027, n68024, n68025, n67775, 
        n67776, n65514, n65520, n65511, n66007, n66908, n65517, 
        n36_adj_5105, n38_adj_5106, n66709, n61682, n67686, n65985, 
        n34_adj_5108, n68327, n62104, n61944, n67773, n62657, n62743, 
        n67774, n65999, n66902, n34_adj_5109, n67688, n66711, n67771, 
        n67772, n48_adj_5110, n68353, n67796, n29_adj_5111, n65970, 
        n41_adj_5112, n39_adj_5113, n40_adj_5114, n28_adj_5115, n33_adj_5116, 
        n35_adj_5117, n37_adj_5118, n29_adj_5119, n31_adj_5120, n67765, 
        n23_adj_5121, n67766, n25_adj_5122, n7, n45_adj_5123, n43_adj_5124, 
        n39_adj_5125, n65957, n11, n68022, n13, n15_adj_5126, n66717, 
        n68322, n68323, n27_adj_5127, n9, n48_adj_5128, n19_adj_5129, 
        n21_adj_5130, n17_adj_5131, n66175, n66191, n16_adj_5132, 
        n27_adj_5133, n33_adj_5134, n31_adj_5135, n29_adj_5136, n65937, 
        n66117, n8_adj_5137, n24_adj_5138, n3274, n66209, n67072, 
        n67064, n68078, n67499, n68209, n41_adj_5139, n38_adj_5140, 
        n12_adj_5141, n48_adj_5142, n4_adj_5143, n67674, n67675, n67763, 
        n66154, n35_adj_5144, n67764, n39_adj_5145, n37_adj_5146, 
        n65933, n10_adj_5147, n30_adj_5148, n68183, n66160, n68058, 
        n66779, n68282, n68283, n6_adj_5149, n67676, n67677, n66719, 
        n68314, n66125, n67729, n66777, n68236, n66127, n68161, 
        n66785, n68315, n61572, n61114, n3253, n68163, n61122, 
        n48_adj_5150, n61608, n33_adj_5151, n31_adj_5152, n37_adj_5153, 
        n35_adj_5154, n25_adj_5155, n27_adj_5156, n21_adj_5157, n23_adj_5158, 
        n9_adj_5159, n29_adj_5160, n11_adj_5161, n31_adj_5162, n19_adj_5163, 
        n13_adj_5164, n15_adj_5165, n17_adj_5166, n33_adj_5167, n29_adj_5168, 
        n66251, n27_adj_5169, n67144, n67553, n65920, n67549, n66267, 
        n6_adj_5170, n67682, n32_adj_5171, n67683, n66245, n68026, 
        n66765, n67731, n67732, n67126, n67727, n66763, n67901, 
        n41_adj_5172, n38_adj_5173, n68246, n67969, n68350, n59314, 
        n68351, n26_adj_5174, n68239, n67759, n68154, n35_adj_5175, 
        n67760, n39_adj_5176, n37_adj_5177, n65910, n39_adj_5178, 
        n68030, n35_adj_5179, n33_adj_5180, n37_adj_5181, n27_adj_5182, 
        n29_adj_5183, n23_adj_5184, n25_adj_5185, n11_adj_5186, n66727, 
        n68316, n13_adj_5187, n21_adj_5188, n68317, n15_adj_5189, 
        n48_adj_5190, n17_adj_5191, n19_adj_5192, n31_adj_5193, n66367, 
        n61998, n67224, n67591, n67587, n66369, n62006, n8_adj_5194, 
        n67739, n67740, n21_adj_5195, n34_adj_5196, n27_adj_5197, 
        n25_adj_5198, n23_adj_5199, n65857, n33_adj_5200, n31_adj_5201, 
        n29_adj_5202, n65852, n66351, n68004, n66755, n67741, n67742, 
        n67200, n20_adj_5203, n66753, n67913, n68320, n67723, n68348, 
        n68349, n67795, n28_adj_5204, n37_adj_5205, n41_adj_5206, 
        n35_adj_5207, n35_adj_5208, n32_adj_5209, n68244, n39_adj_5210, 
        n37_adj_5211, n68245, n29_adj_5212, n39_adj_5213, n68243, 
        n67733, n31_adj_5214, n68185, n41_adj_5215, n40_adj_5216, 
        n68257, n68258, n68198, n23_adj_5217, n25_adj_5218, n27_adj_5219, 
        n13_adj_5220, n15_adj_5221, n17_adj_5222, n19_adj_5223, n21_adj_5224, 
        n33_adj_5225, n66466, n66515, n67282, n67276, n66468, n10_adj_5226, 
        n25_adj_5227, n67747, n67748, n27_adj_5228, n36_adj_5229, 
        n66458, n39_adj_5230, n68002, n66743, n43_adj_5231, n41_adj_5232, 
        n22_adj_5233, n68195, n68196, n33_adj_5234, n68009, n67927, 
        n35_adj_5235, n37_adj_5236, n68318, n66741, n29_adj_5237, 
        n31_adj_5238, n21_adj_5239, n23_adj_5240, n68354, n68355, 
        n39_adj_5241, n43_adj_5242, n37_adj_5243, n41_adj_5244, n43_adj_5245, 
        n39_adj_5246, n41_adj_5247, n31_adj_5248, n33_adj_5249, n37_adj_5250, 
        n25_adj_5251, n27_adj_5252, n29_adj_5253, n31_adj_5254, n25_adj_5255, 
        n33_adj_5256, n35_adj_5257, n23_adj_5258, n65896, n27_adj_5259, 
        n29_adj_5260, n65887, n19_adj_5261, n22_adj_5262, n30_adj_5263, 
        n34_adj_5264, n67783, n65797, n65791, n67672, n67815, n67784, 
        n67754, n67749, n15_adj_5265, n67816, n67825, n66737, n68020, 
        n68021, n17_adj_5266, n19_adj_5267, n66621, n21_adj_5268, 
        n23_adj_5269, n35_adj_5270, n65633, n66549, n26_adj_5271, 
        n67298, n67296, n65635, n12_adj_5272, n67799, n42_adj_5273, 
        n38_adj_5274, n67800, n65627, n67797, n67720, n24_adj_5275, 
        n68193, n68194, n68011, n30_adj_5276, n67627, n68165, n67995, 
        n68326, n68187, n43_adj_5277, n37_adj_5278, n39_adj_5279, 
        n41_adj_5280, n68188, n61974, n59323, n32_adj_5281, n68017, 
        n67769, n67770, n66890, n67690, n66714, n67767;
    
    SB_LUT4 i50342_4_lut (.I0(n67986), .I1(n67356), .I2(n45), .I3(n66623), 
            .O(n67358));   // verilog/uart_rx.v(119[33:55])
    defparam i50342_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7651[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n7677[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2650_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n51750), 
            .O(n7885[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2650_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n51749), 
            .O(n7885[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2650_19 (.CI(n51749), .I0(n2714), .I1(n2867), .CO(n51750));
    SB_LUT4 add_2650_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n51748), 
            .O(n7885[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_18 (.CI(n51748), .I0(n2715), .I1(n2754), .CO(n51749));
    SB_LUT4 add_2650_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n51747), 
            .O(n7885[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_17 (.CI(n51747), .I0(n2716), .I1(n2638), .CO(n51748));
    SB_LUT4 add_2650_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n51746), 
            .O(n7885[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_16 (.CI(n51746), .I0(n2717), .I1(n2519), .CO(n51747));
    SB_LUT4 add_2650_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n51745), 
            .O(n7885[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_15 (.CI(n51745), .I0(n2718), .I1(n2397), .CO(n51746));
    SB_LUT4 add_2650_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n51744), 
            .O(n7885[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_14 (.CI(n51744), .I0(n2719), .I1(n2272), .CO(n51745));
    SB_LUT4 add_2650_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n51743), 
            .O(n7885[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_13 (.CI(n51743), .I0(n2720), .I1(n2144), .CO(n51744));
    SB_LUT4 add_2650_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n51742), 
            .O(n7885[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_12 (.CI(n51742), .I0(n2721), .I1(n2013), .CO(n51743));
    SB_LUT4 add_2650_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n51741), 
            .O(n7885[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2650_11 (.CI(n51741), .I0(n2722), .I1(n1879), .CO(n51742));
    SB_LUT4 add_2650_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n51740), 
            .O(n7885[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_10 (.CI(n51740), .I0(n2723), .I1(n1742), .CO(n51741));
    SB_LUT4 add_2650_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n51739), 
            .O(n7885[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2650_9 (.CI(n51739), .I0(n2724), .I1(n1602), .CO(n51740));
    SB_LUT4 add_2650_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n51738), 
            .O(n7885[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_8 (.CI(n51738), .I0(n2725), .I1(n1459), .CO(n51739));
    SB_LUT4 add_2650_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n51737), 
            .O(n7885[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_7 (.CI(n51737), .I0(n2726), .I1(n1460), .CO(n51738));
    SB_LUT4 add_2650_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n51736), 
            .O(n7885[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_6 (.CI(n51736), .I0(n2727), .I1(n1011), .CO(n51737));
    SB_LUT4 add_2650_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n51735), 
            .O(n7885[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2650_5 (.CI(n51735), .I0(n2728), .I1(n856), .CO(n51736));
    SB_LUT4 add_2650_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n51734), 
            .O(n7885[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_4 (.CI(n51734), .I0(n2729), .I1(n698), .CO(n51735));
    SB_LUT4 add_2650_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n51733), 
            .O(n7885[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2650_3 (.CI(n51733), .I0(n2730), .I1(n858), .CO(n51734));
    SB_LUT4 add_2650_2_lut (.I0(n59295), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2650_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2650_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51733));
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2649_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n51717), 
            .O(n7859[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2649_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n51716), 
            .O(n7859[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_18 (.CI(n51716), .I0(n2597), .I1(n2754), .CO(n51717));
    SB_LUT4 add_2649_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n51715), 
            .O(n7859[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_17 (.CI(n51715), .I0(n2598), .I1(n2638), .CO(n51716));
    SB_LUT4 add_2649_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n51714), 
            .O(n7859[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_16 (.CI(n51714), .I0(n2599), .I1(n2519), .CO(n51715));
    SB_LUT4 add_2649_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n51713), 
            .O(n7859[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_15 (.CI(n51713), .I0(n2600), .I1(n2397), .CO(n51714));
    SB_LUT4 add_2649_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n51712), 
            .O(n7859[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_14 (.CI(n51712), .I0(n2601), .I1(n2272), .CO(n51713));
    SB_LUT4 add_2649_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n51711), 
            .O(n7859[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_13 (.CI(n51711), .I0(n2602), .I1(n2144), .CO(n51712));
    SB_LUT4 add_2649_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n51710), 
            .O(n7859[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_12 (.CI(n51710), .I0(n2603), .I1(n2013), .CO(n51711));
    SB_LUT4 add_2649_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n51709), 
            .O(n7859[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_11 (.CI(n51709), .I0(n2604), .I1(n1879), .CO(n51710));
    SB_LUT4 add_2649_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n51708), 
            .O(n7859[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_10 (.CI(n51708), .I0(n2605), .I1(n1742), .CO(n51709));
    SB_LUT4 add_2649_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n51707), 
            .O(n7859[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_9 (.CI(n51707), .I0(n2606), .I1(n1602), .CO(n51708));
    SB_LUT4 add_2649_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n51706), 
            .O(n7859[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_8 (.CI(n51706), .I0(n2607), .I1(n1459), .CO(n51707));
    SB_LUT4 add_2649_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n51705), 
            .O(n7859[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_7 (.CI(n51705), .I0(n2608), .I1(n1460), .CO(n51706));
    SB_LUT4 add_2649_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n51704), 
            .O(n7859[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_6 (.CI(n51704), .I0(n2609), .I1(n1011), .CO(n51705));
    SB_LUT4 add_2649_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n51703), 
            .O(n7859[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_5 (.CI(n51703), .I0(n2610), .I1(n856), .CO(n51704));
    SB_LUT4 add_2649_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n51702), 
            .O(n7859[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2649_4 (.CI(n51702), .I0(n2611), .I1(n698), .CO(n51703));
    SB_LUT4 add_2649_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n51701), 
            .O(n7859[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48653_4_lut (.I0(n37), .I1(n25), .I2(n23_c), .I3(n21), 
            .O(n65669));
    defparam i48653_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2649_3 (.CI(n51701), .I0(n2612), .I1(n858), .CO(n51702));
    SB_LUT4 add_2649_2_lut (.I0(n59299), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2649_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2649_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51701));
    SB_LUT4 i49563_4_lut (.I0(n19), .I1(n17), .I2(n2729), .I3(baudrate[2]), 
            .O(n66579));
    defparam i49563_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50298_4_lut (.I0(n25), .I1(n23_c), .I2(n21), .I3(n66579), 
            .O(n67314));
    defparam i50298_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50296_4_lut (.I0(n31), .I1(n29_c), .I2(n27_c), .I3(n67314), 
            .O(n67312));
    defparam i50296_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5006));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7651[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n7677[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48656_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67312), 
            .O(n65672));
    defparam i48656_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut (.I0(n61166), .I1(n48), .I2(GND_net), .I3(GND_net), 
            .O(n2491));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n7833[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50787_3_lut (.I0(n14), .I1(baudrate[13]), .I2(n37), .I3(GND_net), 
            .O(n67803));   // verilog/uart_rx.v(119[33:55])
    defparam i50787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50788_3_lut (.I0(n67803), .I1(baudrate[14]), .I2(n39), .I3(GND_net), 
            .O(n67804));   // verilog/uart_rx.v(119[33:55])
    defparam i50788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22), .I1(baudrate[17]), 
            .I2(n45_adj_5007), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48649_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n65669), 
            .O(n65665));
    defparam i48649_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50345_4_lut (.I0(n40), .I1(n20), .I2(n45_adj_5007), .I3(n65659), 
            .O(n67361));   // verilog/uart_rx.v(119[33:55])
    defparam i50345_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50700_3_lut (.I0(n67804), .I1(baudrate[15]), .I2(n41), .I3(GND_net), 
            .O(n67716));   // verilog/uart_rx.v(119[33:55])
    defparam i50700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n62002), .I1(n61148), .I2(n61146), .I3(n61992), 
            .O(n25206));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18), .I1(baudrate[9]), 
            .I2(n29_c), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51175_4_lut (.I0(n26), .I1(n16), .I2(n29_c), .I3(n65690), 
            .O(n68191));   // verilog/uart_rx.v(119[33:55])
    defparam i51175_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 r_Clock_Count_1944_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n52174), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1944_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n52173), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_8 (.CI(n52173), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n52174));
    SB_LUT4 r_Clock_Count_1944_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n52172), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_7 (.CI(n52172), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n52173));
    SB_LUT4 r_Clock_Count_1944_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n52171), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_6 (.CI(n52171), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n52172));
    SB_LUT4 r_Clock_Count_1944_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n52170), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_5 (.CI(n52170), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n52171));
    SB_LUT4 r_Clock_Count_1944_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n52169), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_4 (.CI(n52169), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n52170));
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5012));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Clock_Count_1944_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n52168), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_3 (.CI(n52168), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n52169));
    SB_LUT4 r_Clock_Count_1944_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1944_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1944_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n52168));
    SB_LUT4 i51176_3_lut (.I0(n68191), .I1(baudrate[10]), .I2(n31), .I3(GND_net), 
            .O(n68192));   // verilog/uart_rx.v(119[33:55])
    defparam i51176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50997_3_lut (.I0(n68192), .I1(baudrate[11]), .I2(n33), .I3(GND_net), 
            .O(n68013));   // verilog/uart_rx.v(119[33:55])
    defparam i50997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2648_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n51666), 
            .O(n7833[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50615_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n65672), 
            .O(n67631));
    defparam i50615_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2648_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n51665), 
            .O(n7833[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_17 (.CI(n51665), .I0(n2477), .I1(n2638), .CO(n51666));
    SB_LUT4 add_2648_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n51664), 
            .O(n7833[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_16 (.CI(n51664), .I0(n2478), .I1(n2519), .CO(n51665));
    SB_LUT4 add_2648_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n51663), 
            .O(n7833[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_15 (.CI(n51663), .I0(n2479), .I1(n2397), .CO(n51664));
    SB_LUT4 add_2648_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n51662), 
            .O(n7833[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_14 (.CI(n51662), .I0(n2480), .I1(n2272), .CO(n51663));
    SB_LUT4 i50975_4_lut (.I0(n67716), .I1(n67361), .I2(n45_adj_5007), 
            .I3(n65665), .O(n67991));   // verilog/uart_rx.v(119[33:55])
    defparam i50975_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2648_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n51661), 
            .O(n7833[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_13 (.CI(n51661), .I0(n2481), .I1(n2144), .CO(n51662));
    SB_LUT4 add_2648_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n51660), 
            .O(n7833[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_12 (.CI(n51660), .I0(n2482), .I1(n2013), .CO(n51661));
    SB_LUT4 i50974_3_lut (.I0(n68013), .I1(baudrate[12]), .I2(n35), .I3(GND_net), 
            .O(n67990));   // verilog/uart_rx.v(119[33:55])
    defparam i50974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7651[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2648_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n51659), 
            .O(n7833[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_11 (.CI(n51659), .I0(n2483), .I1(n1879), .CO(n51660));
    SB_LUT4 add_2648_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n51658), 
            .O(n7833[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_10 (.CI(n51658), .I0(n2484), .I1(n1742), .CO(n51659));
    SB_LUT4 add_2648_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n51657), 
            .O(n7833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_9 (.CI(n51657), .I0(n2485), .I1(n1602), .CO(n51658));
    SB_LUT4 add_2648_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n51656), 
            .O(n7833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_8 (.CI(n51656), .I0(n2486), .I1(n1459), .CO(n51657));
    SB_LUT4 add_2648_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n51655), 
            .O(n7833[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_7 (.CI(n51655), .I0(n2487), .I1(n1460), .CO(n51656));
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5014));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2648_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n51654), 
            .O(n7833[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_6 (.CI(n51654), .I0(n2488), .I1(n1011), .CO(n51655));
    SB_LUT4 add_2648_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n51653), 
            .O(n7833[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_5 (.CI(n51653), .I0(n2489), .I1(n856), .CO(n51654));
    SB_LUT4 add_2648_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n51652), 
            .O(n7833[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_4 (.CI(n51652), .I0(n2490), .I1(n698), .CO(n51653));
    SB_LUT4 i48725_4_lut (.I0(n23_adj_5015), .I1(n21_adj_5016), .I2(n19_adj_5017), 
            .I3(n17_adj_5014), .O(n65741));
    defparam i48725_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2648_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n51651), 
            .O(n7833[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2648_3 (.CI(n51651), .I0(n2491), .I1(n858), .CO(n51652));
    SB_LUT4 add_2648_2_lut (.I0(n59303), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2648_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2648_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51651));
    SB_LUT4 i50977_4_lut (.I0(n67990), .I1(n67991), .I2(n45_adj_5007), 
            .I3(n67631), .O(n67993));   // verilog/uart_rx.v(119[33:55])
    defparam i50977_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n51278), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7651[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n61066), .I1(n25117), .I2(VCC_net), 
            .I3(n51277), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_25 (.CI(n51277), .I0(n25117), .I1(VCC_net), 
            .CO(n51278));
    SB_LUT4 sub_38_add_2_24_lut (.I0(n61210), .I1(n62747), .I2(VCC_net), 
            .I3(n51276), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_24 (.CI(n51276), .I0(n62747), .I1(VCC_net), 
            .CO(n51277));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n51275), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_23 (.CI(n51275), .I0(n294[21]), .I1(VCC_net), 
            .CO(n51276));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n61208), .I1(n294[20]), .I2(VCC_net), 
            .I3(n51274), .O(n61210)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2647_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n51632), 
            .O(n7807[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2647_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n51631), 
            .O(n7807[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_22 (.CI(n51274), .I0(n294[20]), .I1(VCC_net), 
            .CO(n51275));
    SB_LUT4 sub_38_add_2_21_lut (.I0(n61206), .I1(n294[19]), .I2(VCC_net), 
            .I3(n51273), .O(n61208)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n7677[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2647_16 (.CI(n51631), .I0(n2354), .I1(n2519), .CO(n51632));
    SB_LUT4 add_2647_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n51630), 
            .O(n7807[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_21 (.CI(n51273), .I0(n294[19]), .I1(VCC_net), 
            .CO(n51274));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n51272), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_15 (.CI(n51630), .I0(n2355), .I1(n2397), .CO(n51631));
    SB_LUT4 add_2647_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n51629), 
            .O(n7807[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n51272), .I0(n294[18]), .I1(VCC_net), 
            .CO(n51273));
    SB_LUT4 i48716_4_lut (.I0(n29_adj_5021), .I1(n27_adj_5022), .I2(n25_adj_5023), 
            .I3(n65741), .O(n65732));
    defparam i48716_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 sub_38_add_2_19_lut (.I0(n61204), .I1(n294[17]), .I2(VCC_net), 
            .I3(n51271), .O(n61206)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i50630_4_lut (.I0(n35_adj_5024), .I1(n33_adj_5025), .I2(n31_adj_5026), 
            .I3(n65732), .O(n67646));
    defparam i50630_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2647_14 (.CI(n51629), .I0(n2356), .I1(n2272), .CO(n51630));
    SB_CARRY sub_38_add_2_19 (.CI(n51271), .I0(n294[17]), .I1(VCC_net), 
            .CO(n51272));
    SB_LUT4 add_2647_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n51628), 
            .O(n7807[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7651[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_18_lut (.I0(n61202), .I1(n294[16]), .I2(VCC_net), 
            .I3(n51270), .O(n61204)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n7677[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_18 (.CI(n51270), .I0(n294[16]), .I1(VCC_net), 
            .CO(n51271));
    SB_CARRY add_2647_13 (.CI(n51628), .I0(n2357), .I1(n2144), .CO(n51629));
    SB_LUT4 add_2647_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n51627), 
            .O(n7807[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n61064), .I1(n294[15]), .I2(VCC_net), 
            .I3(n51269), .O(n61066)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_17 (.CI(n51269), .I0(n294[15]), .I1(VCC_net), 
            .CO(n51270));
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n7677[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2647_12 (.CI(n51627), .I0(n2358), .I1(n2013), .CO(n51628));
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2647_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n51626), 
            .O(n7807[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_11 (.CI(n51626), .I0(n2359), .I1(n1879), .CO(n51627));
    SB_LUT4 add_2647_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n51625), 
            .O(n7807[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_10 (.CI(n51625), .I0(n2360), .I1(n1742), .CO(n51626));
    SB_LUT4 add_2647_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n51624), 
            .O(n7807[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_9 (.CI(n51624), .I0(n2361), .I1(n1602), .CO(n51625));
    SB_LUT4 add_2647_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n51623), 
            .O(n7807[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_8 (.CI(n51623), .I0(n2362), .I1(n1459), .CO(n51624));
    SB_LUT4 add_2647_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n51622), 
            .O(n7807[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_7 (.CI(n51622), .I0(n2363), .I1(n1460), .CO(n51623));
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50793_3_lut (.I0(n16_adj_5027), .I1(baudrate[13]), .I2(n39_adj_5029), 
            .I3(GND_net), .O(n67809));   // verilog/uart_rx.v(119[33:55])
    defparam i50793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n61200), .I1(n294[14]), .I2(VCC_net), 
            .I3(n51268), .O(n61202)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2647_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n51621), 
            .O(n7807[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_6 (.CI(n51621), .I0(n2364), .I1(n1011), .CO(n51622));
    SB_LUT4 add_2647_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n51620), 
            .O(n7807[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_16 (.CI(n51268), .I0(n294[14]), .I1(VCC_net), 
            .CO(n51269));
    SB_CARRY add_2647_5 (.CI(n51620), .I0(n2365), .I1(n856), .CO(n51621));
    SB_LUT4 add_2647_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n51619), 
            .O(n7807[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n51267), .O(n61200)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i50794_3_lut (.I0(n67809), .I1(baudrate[14]), .I2(n41_adj_5030), 
            .I3(GND_net), .O(n67810));   // verilog/uart_rx.v(119[33:55])
    defparam i50794_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_15 (.CI(n51267), .I0(n294[13]), .I1(VCC_net), 
            .CO(n51268));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n51266), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_4 (.CI(n51619), .I0(n2366), .I1(n698), .CO(n51620));
    SB_LUT4 add_2647_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n51618), 
            .O(n7807[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2647_3 (.CI(n51618), .I0(n2367), .I1(n858), .CO(n51619));
    SB_LUT4 add_2647_2_lut (.I0(n59307), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2647_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_38_add_2_14 (.CI(n51266), .I0(n294[12]), .I1(VCC_net), 
            .CO(n51267));
    SB_CARRY add_2647_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51618));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n51265), .O(n61064)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n51265), .I0(n294[11]), .I1(VCC_net), 
            .CO(n51266));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n51264), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n51264), .I0(n294[10]), .I1(VCC_net), 
            .CO(n51265));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n51263), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n51263), .I0(n294[9]), .I1(VCC_net), 
            .CO(n51264));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n51262), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_10 (.CI(n51262), .I0(n294[8]), .I1(VCC_net), 
            .CO(n51263));
    SB_LUT4 i49569_4_lut (.I0(n41_adj_5030), .I1(n39_adj_5029), .I2(n27_adj_5022), 
            .I3(n65737), .O(n66585));
    defparam i49569_4_lut.LUT_INIT = 16'heeef;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n51261), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY sub_38_add_2_9 (.CI(n51261), .I0(n294[7]), .I1(VCC_net), 
            .CO(n51262));
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 i50343_3_lut (.I0(n22_adj_5031), .I1(baudrate[7]), .I2(n27_adj_5022), 
            .I3(GND_net), .O(n67359));   // verilog/uart_rx.v(119[33:55])
    defparam i50343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n51260), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50693_3_lut (.I0(n67810), .I1(baudrate[15]), .I2(n43_adj_5032), 
            .I3(GND_net), .O(n67709));   // verilog/uart_rx.v(119[33:55])
    defparam i50693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49001_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n66017));   // verilog/uart_rx.v(119[33:55])
    defparam i49001_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY sub_38_add_2_8 (.CI(n51260), .I0(n294[6]), .I1(VCC_net), 
            .CO(n51261));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n51259), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n51259), .I0(n294[5]), .I1(VCC_net), 
            .CO(n51260));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n51258), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n51258), .I0(n294[4]), .I1(VCC_net), 
            .CO(n51259));
    SB_LUT4 add_2646_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n51601), 
            .O(n7781[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n51257), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2646_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n51600), 
            .O(n7781[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_15 (.CI(n51600), .I0(n2228), .I1(n2397), .CO(n51601));
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5035), .I1(baudrate[9]), 
            .I2(n31_adj_5026), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2646_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n51599), 
            .O(n7781[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_14 (.CI(n51599), .I0(n2229), .I1(n2272), .CO(n51600));
    SB_LUT4 add_2646_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n51598), 
            .O(n7781[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n51257), .I0(n294[3]), .I1(VCC_net), 
            .CO(n51258));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n51256), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_13 (.CI(n51598), .I0(n2230), .I1(n2144), .CO(n51599));
    SB_LUT4 add_2646_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n51597), 
            .O(n7781[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51173_4_lut (.I0(n28), .I1(n18_adj_5036), .I2(n31_adj_5026), 
            .I3(n65729), .O(n68189));   // verilog/uart_rx.v(119[33:55])
    defparam i51173_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2646_12 (.CI(n51597), .I0(n2231), .I1(n2013), .CO(n51598));
    SB_CARRY sub_38_add_2_4 (.CI(n51256), .I0(n294[2]), .I1(VCC_net), 
            .CO(n51257));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n51255), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2646_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n51596), 
            .O(n7781[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_11 (.CI(n51596), .I0(n2232), .I1(n1879), .CO(n51597));
    SB_CARRY sub_38_add_2_3 (.CI(n51255), .I0(n294[1]), .I1(VCC_net), 
            .CO(n51256));
    SB_LUT4 add_2646_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n51595), 
            .O(n7781[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_10 (.CI(n51595), .I0(n2233), .I1(n1742), .CO(n51596));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n60086), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51174_3_lut (.I0(n68189), .I1(baudrate[10]), .I2(n33_adj_5025), 
            .I3(GND_net), .O(n68190));   // verilog/uart_rx.v(119[33:55])
    defparam i51174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2646_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n51594), 
            .O(n7781[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50999_3_lut (.I0(n68190), .I1(baudrate[11]), .I2(n35_adj_5024), 
            .I3(GND_net), .O(n68015));   // verilog/uart_rx.v(119[33:55])
    defparam i50999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49573_4_lut (.I0(n41_adj_5030), .I1(n39_adj_5029), .I2(n37_adj_5038), 
            .I3(n67646), .O(n66589));
    defparam i49573_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2646_9 (.CI(n51594), .I0(n2234), .I1(n1602), .CO(n51595));
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n60086), .I1(GND_net), 
            .CO(n51255));
    SB_LUT4 i50791_4_lut (.I0(n67709), .I1(n67359), .I2(n43_adj_5032), 
            .I3(n66585), .O(n67807));   // verilog/uart_rx.v(119[33:55])
    defparam i50791_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50972_3_lut (.I0(n68015), .I1(baudrate[12]), .I2(n37_adj_5038), 
            .I3(GND_net), .O(n67988));   // verilog/uart_rx.v(119[33:55])
    defparam i50972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2646_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n51593), 
            .O(n7781[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_8 (.CI(n51593), .I0(n2235), .I1(n1459), .CO(n51594));
    SB_LUT4 i51185_4_lut (.I0(n67988), .I1(n67807), .I2(n43_adj_5032), 
            .I3(n66589), .O(n68201));   // verilog/uart_rx.v(119[33:55])
    defparam i51185_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2646_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n51592), 
            .O(n7781[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7651[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51186_3_lut (.I0(n68201), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n68202));   // verilog/uart_rx.v(119[33:55])
    defparam i51186_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2646_7 (.CI(n51592), .I0(n2236), .I1(n1460), .CO(n51593));
    SB_LUT4 add_2646_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n51591), 
            .O(n7781[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_6 (.CI(n51591), .I0(n2237), .I1(n1011), .CO(n51592));
    SB_LUT4 add_2646_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n51590), 
            .O(n7781[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n7677[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2646_5 (.CI(n51590), .I0(n2238), .I1(n856), .CO(n51591));
    SB_LUT4 add_2646_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n51589), 
            .O(n7781[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7625[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7625[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n7833[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7625[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n7859[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2646_4 (.CI(n51589), .I0(n2239), .I1(n698), .CO(n51590));
    SB_LUT4 i1_3_lut (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4894), 
            .I3(GND_net), .O(n61126));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_983 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n61126), .O(\r_SM_Main_2__N_3536[1] ));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_983.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7625[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7625[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2646_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n51588), 
            .O(n7781[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2646_3 (.CI(n51588), .I0(n2240), .I1(n858), .CO(n51589));
    SB_LUT4 i1_2_lut_4_lut (.I0(n68202), .I1(baudrate[17]), .I2(n2596), 
            .I3(n61170), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 add_2646_2_lut (.I0(n59311), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2646_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2646_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51588));
    SB_LUT4 i51446_2_lut_4_lut (.I0(n68202), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25206), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i51446_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7625[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_984 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4894), .I2(n57758), 
            .I3(GND_net), .O(n61284));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_adj_984.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_985 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61284), .O(n61290));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_985.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2645_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n51577), 
            .O(n7755[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7625[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2645_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n51576), 
            .O(n7755[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_13 (.CI(n51576), .I0(n2099), .I1(n2272), .CO(n51577));
    SB_LUT4 add_2645_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n51575), 
            .O(n7755[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_986 (.I0(n61160), .I1(n48_adj_5044), .I2(GND_net), 
            .I3(GND_net), .O(n1560));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7599[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7573[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_987 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n61884));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_987.LUT_INIT = 16'h7bde;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5034), .I1(baudrate[4]), 
            .I2(n41_adj_5045), .I3(GND_net), .O(n40_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_275_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5047));   // verilog/uart_rx.v(69[17:62])
    defparam equal_275_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51165_4_lut (.I0(n40_adj_5046), .I1(n36), .I2(n41_adj_5045), 
            .I3(n66017), .O(n68181));   // verilog/uart_rx.v(119[33:55])
    defparam i51165_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_988 (.I0(r_Clock_Count[3]), .I1(n3_adj_5047), .I2(\o_Rx_DV_N_3488[4] ), 
            .I3(n61884), .O(n61888));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_988.LUT_INIT = 16'hffde;
    SB_LUT4 equal_275_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_275_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_989 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n61888), .O(n61892));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_989.LUT_INIT = 16'hffde;
    SB_LUT4 i51166_3_lut (.I0(n68181), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n68182));   // verilog/uart_rx.v(119[33:55])
    defparam i51166_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 equal_275_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(69[17:62])
    defparam equal_275_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_990 (.I0(r_Clock_Count[6]), .I1(n8), .I2(n61892), 
            .I3(\o_Rx_DV_N_3488[7] ), .O(n57790));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_4_lut_adj_991 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4891), 
            .I3(\o_Rx_DV_N_3488[8] ), .O(n61104));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_991.LUT_INIT = 16'hfffe;
    SB_LUT4 i51023_3_lut (.I0(n68182), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n68039));   // verilog/uart_rx.v(119[33:55])
    defparam i51023_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_992 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n61104), .O(r_SM_Main_2__N_3446[1]));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i49691_3_lut (.I0(n68039), .I1(baudrate[7]), .I2(n1261), .I3(GND_net), 
            .O(n48_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam i49691_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7573[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n57762));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7599[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i23355_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n39001));
    defparam i23355_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_993 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n57762), .O(n61296));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_993.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_994 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61296), .O(n61302));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_994.LUT_INIT = 16'hfffe;
    SB_LUT4 i45618_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n57790), .I2(GND_net), 
            .I3(GND_net), .O(n62625));
    defparam i45618_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45716_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n62625), .O(n62723));
    defparam i45716_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n61302), .I1(r_SM_Main_2__N_3446[1]), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n62723), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n9679));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i6058_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21487));   // verilog/uart_rx.v(119[33:55])
    defparam i6058_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n9679), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY add_2645_12 (.CI(n51575), .I0(n2100), .I1(n2144), .CO(n51576));
    SB_LUT4 add_2645_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n51574), 
            .O(n7755[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_11 (.CI(n51574), .I0(n2101), .I1(n2013), .CO(n51575));
    SB_LUT4 add_2645_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n51573), 
            .O(n7755[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_10 (.CI(n51573), .I0(n2102), .I1(n1879), .CO(n51574));
    SB_LUT4 add_2645_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n51572), 
            .O(n7755[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_9 (.CI(n51572), .I0(n2103), .I1(n1742), .CO(n51573));
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5050), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i45666_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n62673));
    defparam i45666_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2645_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n51571), 
            .O(n7755[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_5051), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2645_8 (.CI(n51571), .I0(n2104), .I1(n1602), .CO(n51572));
    SB_LUT4 add_2645_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n51570), 
            .O(n7755[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_7 (.CI(n51570), .I0(n2105), .I1(n1459), .CO(n51571));
    SB_LUT4 add_2645_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n51569), 
            .O(n7755[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_6 (.CI(n51569), .I0(n2106), .I1(n1460), .CO(n51570));
    SB_LUT4 add_2645_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n51568), 
            .O(n7755[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5052), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_CARRY add_2645_5 (.CI(n51568), .I0(n2107), .I1(n1011), .CO(n51569));
    SB_DFFESR r_Clock_Count_1944__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27409), .D(n1[0]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 add_2645_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n51567), 
            .O(n7755[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_4 (.CI(n51567), .I0(n2108), .I1(n856), .CO(n51568));
    SB_LUT4 add_2645_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n51566), 
            .O(n7755[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_3 (.CI(n51566), .I0(n2109), .I1(n698), .CO(n51567));
    SB_LUT4 add_2645_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n7755[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2645_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2645_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n51566));
    SB_LUT4 i49341_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4891), .I3(n58022), .O(n65437));
    defparam i49341_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i49332_4_lut (.I0(n65437), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65434));
    defparam i49332_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n65434), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27288));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 add_2644_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n51556), 
            .O(n7729[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2644_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n51555), 
            .O(n7729[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_13 (.CI(n51555), .I0(n1967), .I1(n2144), .CO(n51556));
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7573[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2644_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n51554), 
            .O(n7729[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42010_2_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n58970));
    defparam i42010_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_2644_12 (.CI(n51554), .I0(n1968), .I1(n2013), .CO(n51555));
    SB_LUT4 add_2644_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n51553), 
            .O(n7729[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_11 (.CI(n51553), .I0(n1969), .I1(n1879), .CO(n51554));
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7599[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2644_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n51552), 
            .O(n7729[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_10 (.CI(n51552), .I0(n1970), .I1(n1742), .CO(n51553));
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2644_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n51551), 
            .O(n7729[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_995 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n61964));
    defparam i1_2_lut_4_lut_adj_995.LUT_INIT = 16'hfffe;
    SB_CARRY add_2644_9 (.CI(n51551), .I0(n1971), .I1(n1602), .CO(n51552));
    SB_LUT4 add_2644_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n51550), 
            .O(n7729[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2644_8 (.CI(n51550), .I0(n1972), .I1(n1459), .CO(n51551));
    SB_LUT4 i48773_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n65789));
    defparam i48773_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48627_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n65643));
    defparam i48627_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48609_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n65625));
    defparam i48609_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51538_2_lut_4_lut (.I0(n68260), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25194), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i51538_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2644_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n51549), 
            .O(n7729[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7573[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7599[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61166), .I3(n48), .O(n18_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_CARRY add_2644_7 (.CI(n51549), .I0(n1973), .I1(n1460), .CO(n51550));
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2644_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n51548), 
            .O(n7729[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2644_6 (.CI(n51548), .I0(n1974), .I1(n1011), .CO(n51549));
    SB_LUT4 add_2644_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n51547), 
            .O(n7729[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_5 (.CI(n51547), .I0(n1975), .I1(n856), .CO(n51548));
    SB_LUT4 i48866_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n65882));
    defparam i48866_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48877_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n65893));
    defparam i48877_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48779_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n65795));
    defparam i48779_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51389_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n62711), .I3(n48_adj_5065), .O(n294[19]));
    defparam i51389_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48578_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n65594));
    defparam i48578_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2644_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n51546), 
            .O(n7729[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFESR r_Clock_Count_1944__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27409), .D(n1[7]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1944__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27409), .D(n1[6]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1944__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27409), .D(n1[5]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1944__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27409), .D(n1[4]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1944__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27409), .D(n1[3]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1944__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27409), .D(n1[2]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1944__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27409), .D(n1[1]), .R(n28713));   // verilog/uart_rx.v(121[34:51])
    SB_CARRY add_2644_4 (.CI(n51546), .I0(n1976), .I1(n698), .CO(n51547));
    SB_LUT4 add_2644_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n51545), 
            .O(n7729[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49440_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n66456));
    defparam i49440_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2644_3 (.CI(n51545), .I0(n1977), .I1(n858), .CO(n51546));
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2644_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7729[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2644_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2644_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51545));
    SB_LUT4 add_2643_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n51544), 
            .O(n7703[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5070));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 add_2643_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n51543), 
            .O(n7703[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4891), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5070), 
            .I3(n58022), .O(n69043));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i48831_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n65847));
    defparam i48831_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2643_12 (.CI(n51543), .I0(n1832), .I1(n2013), .CO(n51544));
    SB_LUT4 add_2643_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n51542), 
            .O(n7703[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61164), .I3(n48_adj_5072), .O(n20_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i48838_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n65854));
    defparam i48838_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 equal_353_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(98[17:39])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_996 (.I0(\r_SM_Main[1] ), .I1(n6), .I2(\r_Bit_Index[0] ), 
            .I3(n4), .O(n61664));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_996.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut_adj_997 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61664), .O(n61670));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_998 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61670), .O(n61676));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_998.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_999 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61592), .O(n61598));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1000 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61598), .O(n61604));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_CARRY add_2643_11 (.CI(n51542), .I0(n1833), .I1(n1879), .CO(n51543));
    SB_LUT4 add_2643_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n51541), 
            .O(n7703[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_10 (.CI(n51541), .I0(n1834), .I1(n1742), .CO(n51542));
    SB_LUT4 add_2643_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n51540), 
            .O(n7703[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_9 (.CI(n51540), .I0(n1835), .I1(n1602), .CO(n51541));
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49415_4_lut (.I0(n25163), .I1(n65779), .I2(n48_adj_5076), 
            .I3(baudrate[0]), .O(n804));
    defparam i49415_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i49330_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n66346));
    defparam i49330_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_2643_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n51539), 
            .O(n7703[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49386_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n66402));
    defparam i49386_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2643_8 (.CI(n51539), .I0(n1836), .I1(n1459), .CO(n51540));
    SB_LUT4 add_2643_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n51538), 
            .O(n7703[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_7 (.CI(n51538), .I0(n1837), .I1(n1460), .CO(n51539));
    SB_LUT4 add_2643_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n51537), 
            .O(n7703[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_6 (.CI(n51537), .I0(n1838), .I1(n1011), .CO(n51538));
    SB_LUT4 add_2643_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n51536), 
            .O(n7703[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_5 (.CI(n51536), .I0(n1839), .I1(n856), .CO(n51537));
    SB_LUT4 add_2643_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n51535), 
            .O(n7703[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_4 (.CI(n51535), .I0(n1840), .I1(n698), .CO(n51536));
    SB_LUT4 add_2643_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n51534), 
            .O(n7703[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2643_3 (.CI(n51534), .I0(n1841), .I1(n858), .CO(n51535));
    SB_LUT4 add_2643_2_lut (.I0(n59320), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2643_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2643_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51534));
    SB_LUT4 add_2642_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n51533), 
            .O(n7677[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61646), .O(n61652));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2642_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n51532), 
            .O(n7677[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_10 (.CI(n51532), .I0(n1694), .I1(n1879), .CO(n51533));
    SB_LUT4 add_2642_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n51531), 
            .O(n7677[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_9 (.CI(n51531), .I0(n1695), .I1(n1742), .CO(n51532));
    SB_LUT4 i1_4_lut_adj_1002 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61652), .O(n61658));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 i50769_3_lut (.I0(n42_adj_5079), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n67785));   // verilog/uart_rx.v(119[33:55])
    defparam i50769_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2642_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n51530), 
            .O(n7677[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_8 (.CI(n51530), .I0(n1696), .I1(n1602), .CO(n51531));
    SB_LUT4 i50770_3_lut (.I0(n67785), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n67786));   // verilog/uart_rx.v(119[33:55])
    defparam i50770_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n67786), .I1(baudrate[4]), 
            .I2(n58994), .I3(GND_net), .O(n48_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[27]), 
            .I3(baudrate[24]), .O(n61146));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n61988));
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'heeee;
    SB_LUT4 i51535_2_lut_4_lut (.I0(n68155), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25221), .O(n294[1]));
    defparam i51535_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2642_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n51529), 
            .O(n7677[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_7 (.CI(n51529), .I0(n1697), .I1(n1459), .CO(n51530));
    SB_LUT4 i1_4_lut_adj_1004 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61628), .O(n61634));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n61942));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61634), .O(n61640));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2642_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n51528), 
            .O(n7677[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n61992));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n61994));
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'heeee;
    SB_CARRY add_2642_6 (.CI(n51528), .I0(n1698), .I1(n1460), .CO(n51529));
    SB_LUT4 add_2642_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n51527), 
            .O(n7677[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n61872));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'hfffe;
    SB_CARRY add_2642_5 (.CI(n51527), .I0(n1699), .I1(n1011), .CO(n51528));
    SB_LUT4 i1_4_lut_adj_1010 (.I0(n61872), .I1(n62002), .I2(n61946), 
            .I3(n61942), .O(n25212));
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 i23357_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n39003));
    defparam i23357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48888_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n65904));
    defparam i48888_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n65498), .I1(baudrate[2]), 
            .I2(n68388), .I3(n48_adj_5076), .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61574), .O(n61580));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46), .I1(baudrate[3]), .I2(n58992), 
            .I3(GND_net), .O(n48_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i49227_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n66243));
    defparam i49227_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(n61844), .I1(n61908), .I2(n61910), 
            .I3(n61906), .O(n61856));
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(n61856), .I1(n25212), .I2(n61848), 
            .I3(n62004), .O(n25166));
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1014 (.I0(n25166), .I1(n48_adj_5083), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1014.LUT_INIT = 16'hefef;
    SB_LUT4 i49282_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n66298));
    defparam i49282_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61580), .O(n61586));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'hfffe;
    SB_LUT4 i4094_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam i4094_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n62106));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5086), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7573[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7599[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4109_2_lut (.I0(n21489), .I1(n9470), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam i4109_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5088), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i45494_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62498));
    defparam i45494_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n61710));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n61712));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n62500));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1019 (.I0(baudrate[17]), .I1(n61714), .I2(baudrate[2]), 
            .I3(n39001), .O(n61092));
    defparam i1_4_lut_adj_1019.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1020 (.I0(n62683), .I1(n61092), .I2(n25206), 
            .I3(n62593), .O(n60160));
    defparam i1_4_lut_adj_1020.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n39003), .O(n61442));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1022 (.I0(n61442), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n61460));
    defparam i1_4_lut_adj_1022.LUT_INIT = 16'h0002;
    SB_LUT4 i45732_4_lut (.I0(n62673), .I1(n62593), .I2(n62597), .I3(n62500), 
            .O(n62739));
    defparam i45732_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1023 (.I0(n62719), .I1(n62739), .I2(n59034), 
            .I3(n61460), .O(n59802));
    defparam i1_4_lut_adj_1023.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n61946));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n61990));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61610), .O(n61616));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n61714));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'heeee;
    SB_LUT4 i6048_4_lut (.I0(n804), .I1(n39001), .I2(n21473), .I3(baudrate[2]), 
            .O(n21475));   // verilog/uart_rx.v(119[33:55])
    defparam i6048_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i51417_2_lut_4_lut (.I0(n68262), .I1(baudrate[12]), .I2(n1966), 
            .I3(n62659), .O(n294[11]));
    defparam i51417_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_1028 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61616), .O(n61622));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n61926));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42132_2_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i42132_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45648_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n62655));
    defparam i45648_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n61936));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n61948));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61538), .O(n61544));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i45682_2_lut_3_lut_4_lut (.I0(baudrate[12]), .I1(n62659), .I2(baudrate[10]), 
            .I3(baudrate[11]), .O(n62689));
    defparam i45682_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(n61988), .I1(n61926), .I2(n61730), 
            .I3(baudrate[19]), .O(n61750));
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1033 (.I0(n61750), .I1(n61948), .I2(n61990), 
            .I3(n61946), .O(n25209));
    defparam i1_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61162), .I3(n48_adj_5090), .O(n26_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61544), .O(n61550));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n61706), .I1(n61702), .I2(n61704), 
            .I3(n62500), .O(n61724));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2642_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n51526), 
            .O(n7677[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_4 (.CI(n51526), .I0(n1700), .I1(n856), .CO(n51527));
    SB_LUT4 i1_4_lut_adj_1036 (.I0(n61714), .I1(n61710), .I2(n61712), 
            .I3(n61708), .O(n61726));
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1037 (.I0(n61726), .I1(n25209), .I2(n61724), 
            .I3(GND_net), .O(n25163));
    defparam i1_3_lut_adj_1037.LUT_INIT = 16'hfefe;
    SB_LUT4 add_2642_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n51525), 
            .O(n7677[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_3 (.CI(n51525), .I0(n1701), .I1(n698), .CO(n51526));
    SB_LUT4 add_2642_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n7677[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2642_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2642_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n51525));
    SB_LUT4 add_2641_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n51524), 
            .O(n7651[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2641_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n51523), 
            .O(n7651[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_10 (.CI(n51523), .I0(n1553), .I1(n1742), .CO(n51524));
    SB_LUT4 add_2641_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n51522), 
            .O(n7651[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_9 (.CI(n51522), .I0(n1554), .I1(n1602), .CO(n51523));
    SB_LUT4 add_2641_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n51521), 
            .O(n7651[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2641_8 (.CI(n51521), .I0(n1555), .I1(n1459), .CO(n51522));
    SB_LUT4 add_2641_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n51520), 
            .O(n7651[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_7 (.CI(n51520), .I0(n1556), .I1(n1460), .CO(n51521));
    SB_LUT4 add_2641_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n51519), 
            .O(n7651[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_6 (.CI(n51519), .I0(n1557), .I1(n1011), .CO(n51520));
    SB_LUT4 add_2641_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n51518), 
            .O(n7651[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_5 (.CI(n51518), .I0(n1558), .I1(n856), .CO(n51519));
    SB_LUT4 add_2641_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n51517), 
            .O(n7651[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_4 (.CI(n51517), .I0(n1559), .I1(n698), .CO(n51518));
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n59802), .I1(baudrate[2]), 
            .I2(n60160), .I3(GND_net), .O(n48_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 add_2641_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n51516), 
            .O(n7651[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_3 (.CI(n51516), .I0(n1560), .I1(n858), .CO(n51517));
    SB_LUT4 add_2641_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7651[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2641_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2641_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51516));
    SB_LUT4 i48915_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n65931));
    defparam i48915_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51578_2_lut (.I0(n48_adj_5076), .I1(n25163), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i51578_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45517_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25206), .I3(baudrate[15]), .O(n59311));
    defparam i45517_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i45513_1_lut_2_lut (.I0(baudrate[17]), .I1(n25206), .I2(GND_net), 
            .I3(GND_net), .O(n59303));
    defparam i45513_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n61844));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'heeee;
    SB_LUT4 i42066_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n59034));
    defparam i42066_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51429_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25206), .I3(n48), .O(n294[8]));
    defparam i51429_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i45515_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25206), .I3(GND_net), .O(n59307));
    defparam i45515_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 add_2640_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n51507), 
            .O(n7625[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29912));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29911));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29910));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29909));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29908));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29907));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29906));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n69043));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29663));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .D(n54370));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2640_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n51506), 
            .O(n7625[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_9 (.CI(n51506), .I0(n1409), .I1(n1602), .CO(n51507));
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n29667));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2640_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n51505), 
            .O(n7625[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_8 (.CI(n51505), .I0(n1410), .I1(n1459), .CO(n51506));
    SB_LUT4 add_2640_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n51504), 
            .O(n7625[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_7 (.CI(n51504), .I0(n1411), .I1(n1460), .CO(n51505));
    SB_LUT4 add_2640_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n51503), 
            .O(n7625[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2640_6 (.CI(n51503), .I0(n1412), .I1(n1011), .CO(n51504));
    SB_LUT4 add_2640_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n51502), 
            .O(n7625[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48936_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n65952));
    defparam i48936_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2640_5 (.CI(n51502), .I0(n1413), .I1(n856), .CO(n51503));
    SB_LUT4 add_2640_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n51501), 
            .O(n7625[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_4 (.CI(n51501), .I0(n1414), .I1(n698), .CO(n51502));
    SB_LUT4 add_2640_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n51500), 
            .O(n7625[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2640_3 (.CI(n51500), .I0(n1415), .I1(n858), .CO(n51501));
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2640_2_lut (.I0(n59329), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61160)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2640_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2640_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51500));
    SB_LUT4 add_2639_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n51499), 
            .O(n7599[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(n61916), .I1(n61996), .I2(baudrate[16]), 
            .I3(n39001), .O(n61790));
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'h0100;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27292), 
            .D(n479[1]), .R(n28645));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27292), 
            .D(n479[2]), .R(n28645));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i51532_2_lut_4_lut (.I0(n67768), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25185), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i51532_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61160), .I3(n48_adj_5044), .O(n32_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 add_2639_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n51498), 
            .O(n7599[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_8 (.CI(n51498), .I0(n1262), .I1(n1459), .CO(n51499));
    SB_LUT4 add_2639_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n51497), 
            .O(n7599[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_7 (.CI(n51497), .I0(n1263), .I1(n1460), .CO(n51498));
    SB_LUT4 add_2639_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n51496), 
            .O(n7599[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_6 (.CI(n51496), .I0(n1264), .I1(n1011), .CO(n51497));
    SB_LUT4 add_2639_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n51495), 
            .O(n7599[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_5 (.CI(n51495), .I0(n1265), .I1(n856), .CO(n51496));
    SB_LUT4 add_2639_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n51494), 
            .O(n7599[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49477_3_lut (.I0(n59802), .I1(n60160), .I2(baudrate[2]), 
            .I3(GND_net), .O(n65420));   // verilog/uart_rx.v(119[33:55])
    defparam i49477_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i42322_1_lut (.I0(n25212), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59291));
    defparam i42322_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2639_4 (.CI(n51494), .I0(n1266), .I1(n698), .CO(n51495));
    SB_LUT4 add_2639_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n51493), 
            .O(n7599[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2639_3 (.CI(n51493), .I0(n1267), .I1(n858), .CO(n51494));
    SB_LUT4 add_2639_2_lut (.I0(n59333), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61158)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2639_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2639_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51493));
    SB_LUT4 add_2638_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n51492), 
            .O(n7573[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2638_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n51491), 
            .O(n7573[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_7 (.CI(n51491), .I0(n1112), .I1(n1460), .CO(n51492));
    SB_LUT4 add_2638_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n51490), 
            .O(n7573[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_6 (.CI(n51490), .I0(n1113), .I1(n1011), .CO(n51491));
    SB_LUT4 add_2638_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n51489), 
            .O(n7573[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_5 (.CI(n51489), .I0(n1114), .I1(n856), .CO(n51490));
    SB_LUT4 i49237_4_lut (.I0(n59034), .I1(n61790), .I2(n61918), .I3(n61844), 
            .O(n65421));   // verilog/uart_rx.v(119[33:55])
    defparam i49237_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n65421), .I1(n65420), .I2(n294[21]), 
            .I3(n62516), .O(n58992));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 add_2638_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n51488), 
            .O(n7573[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_4 (.CI(n51488), .I0(n1115), .I1(n698), .CO(n51489));
    SB_LUT4 add_2638_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n51487), 
            .O(n7573[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2638_3 (.CI(n51487), .I0(n1116), .I1(n858), .CO(n51488));
    SB_LUT4 add_2638_2_lut (.I0(n59337), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61156)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2638_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2638_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51487));
    SB_LUT4 i45707_1_lut (.I0(n62713), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59287));
    defparam i45707_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2654_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n51892), 
            .O(n7989[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2654_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n51891), 
            .O(n7989[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_24 (.CI(n51891), .I0(n3152), .I1(n3082), .CO(n51892));
    SB_LUT4 add_2654_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n51890), 
            .O(n7989[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_23 (.CI(n51890), .I0(n3153), .I1(n3188), .CO(n51891));
    SB_LUT4 add_2654_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n51889), 
            .O(n7989[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_22 (.CI(n51889), .I0(n3154), .I1(n3084), .CO(n51890));
    SB_LUT4 i42314_1_lut (.I0(n25218), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59283));
    defparam i42314_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2654_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n51888), 
            .O(n7989[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_21 (.CI(n51888), .I0(n3155), .I1(n2977), .CO(n51889));
    SB_LUT4 add_2654_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n51887), 
            .O(n7989[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_20 (.CI(n51887), .I0(n3156), .I1(n2867), .CO(n51888));
    SB_LUT4 add_2654_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n51886), 
            .O(n7989[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_19 (.CI(n51886), .I0(n3157), .I1(n2754), .CO(n51887));
    SB_LUT4 add_2654_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n51885), 
            .O(n7989[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_18 (.CI(n51885), .I0(n3158), .I1(n2638), .CO(n51886));
    SB_LUT4 add_2654_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n51884), 
            .O(n7989[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i534_3_lut (.I0(n58992), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n58994));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_CARRY add_2654_17 (.CI(n51884), .I0(n3159), .I1(n2519), .CO(n51885));
    SB_LUT4 add_2654_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n51883), 
            .O(n7989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_16 (.CI(n51883), .I0(n3160), .I1(n2397), .CO(n51884));
    SB_LUT4 add_2654_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n51882), 
            .O(n7989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_15 (.CI(n51882), .I0(n3161), .I1(n2272), .CO(n51883));
    SB_LUT4 add_2654_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n51881), 
            .O(n7989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_14 (.CI(n51881), .I0(n3162), .I1(n2144), .CO(n51882));
    SB_LUT4 add_2654_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n51880), 
            .O(n7989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_13 (.CI(n51880), .I0(n3163), .I1(n2013), .CO(n51881));
    SB_LUT4 add_2654_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n51879), 
            .O(n7989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_12 (.CI(n51879), .I0(n3164), .I1(n1879), .CO(n51880));
    SB_LUT4 add_2654_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n51878), 
            .O(n7989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_11 (.CI(n51878), .I0(n3165), .I1(n1742), .CO(n51879));
    SB_LUT4 add_2654_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n51877), 
            .O(n7989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_10 (.CI(n51877), .I0(n3166), .I1(n1602), .CO(n51878));
    SB_LUT4 i1_2_lut_adj_1040 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n61996));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n61904));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'heeee;
    SB_LUT4 add_2654_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n51876), 
            .O(n7989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_9 (.CI(n51876), .I0(n3167), .I1(n1459), .CO(n51877));
    SB_LUT4 add_2654_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n51875), 
            .O(n7989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_8 (.CI(n51875), .I0(n3168), .I1(n1460), .CO(n51876));
    SB_LUT4 add_2654_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n51874), 
            .O(n7989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_7 (.CI(n51874), .I0(n3169), .I1(n1011), .CO(n51875));
    SB_LUT4 add_2654_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n51873), 
            .O(n7989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_6 (.CI(n51873), .I0(n3170), .I1(n856), .CO(n51874));
    SB_LUT4 add_2654_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n51872), 
            .O(n7989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_5 (.CI(n51872), .I0(n3171), .I1(n698), .CO(n51873));
    SB_LUT4 add_2654_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n51871), 
            .O(n7989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_4 (.CI(n51871), .I0(n3172), .I1(n858), .CO(n51872));
    SB_LUT4 add_2654_3_lut (.I0(n59279), .I1(GND_net), .I2(n538), .I3(n51870), 
            .O(n61180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2654_3 (.CI(n51870), .I0(GND_net), .I1(n538), .CO(n51871));
    SB_CARRY add_2654_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n51870));
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n61906));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'heeee;
    SB_LUT4 add_2653_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n51851), 
            .O(n7963[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2653_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n51850), 
            .O(n7963[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_22 (.CI(n51850), .I0(n3047), .I1(n3188), .CO(n51851));
    SB_LUT4 add_2653_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n51849), 
            .O(n7963[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_21 (.CI(n51849), .I0(n3048), .I1(n3084), .CO(n51850));
    SB_LUT4 add_2653_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n51848), 
            .O(n7963[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_20 (.CI(n51848), .I0(n3049), .I1(n2977), .CO(n51849));
    SB_LUT4 add_2653_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n51847), 
            .O(n7963[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_19 (.CI(n51847), .I0(n3050), .I1(n2867), .CO(n51848));
    SB_LUT4 add_2653_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n51846), 
            .O(n7963[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_18 (.CI(n51846), .I0(n3051), .I1(n2754), .CO(n51847));
    SB_LUT4 add_2653_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n51845), 
            .O(n7963[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_17 (.CI(n51845), .I0(n3052), .I1(n2638), .CO(n51846));
    SB_LUT4 add_2653_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n51844), 
            .O(n7963[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_16 (.CI(n51844), .I0(n3053), .I1(n2519), .CO(n51845));
    SB_LUT4 add_2653_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n51843), 
            .O(n7963[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_15 (.CI(n51843), .I0(n3054), .I1(n2397), .CO(n51844));
    SB_LUT4 add_2653_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n51842), 
            .O(n7963[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_14 (.CI(n51842), .I0(n3055), .I1(n2272), .CO(n51843));
    SB_LUT4 add_2653_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n51841), 
            .O(n7963[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_13 (.CI(n51841), .I0(n3056), .I1(n2144), .CO(n51842));
    SB_LUT4 add_2653_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n51840), 
            .O(n7963[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_12 (.CI(n51840), .I0(n3057), .I1(n2013), .CO(n51841));
    SB_LUT4 add_2653_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n51839), 
            .O(n7963[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_11 (.CI(n51839), .I0(n3058), .I1(n1879), .CO(n51840));
    SB_LUT4 add_2653_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n51838), 
            .O(n7963[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_10 (.CI(n51838), .I0(n3059), .I1(n1742), .CO(n51839));
    SB_LUT4 add_2653_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n51837), 
            .O(n7963[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_9 (.CI(n51837), .I0(n3060), .I1(n1602), .CO(n51838));
    SB_LUT4 add_2653_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n51836), 
            .O(n7963[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_8 (.CI(n51836), .I0(n3061), .I1(n1459), .CO(n51837));
    SB_LUT4 add_2653_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n51835), 
            .O(n7963[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_7 (.CI(n51835), .I0(n3062), .I1(n1460), .CO(n51836));
    SB_LUT4 add_2653_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n51834), 
            .O(n7963[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_6 (.CI(n51834), .I0(n3063), .I1(n1011), .CO(n51835));
    SB_LUT4 add_2653_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n51833), 
            .O(n7963[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_5 (.CI(n51833), .I0(n3064), .I1(n856), .CO(n51834));
    SB_LUT4 add_2653_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n51832), 
            .O(n7963[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_4 (.CI(n51832), .I0(n3065), .I1(n698), .CO(n51833));
    SB_LUT4 add_2653_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n51831), 
            .O(n7963[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2653_3 (.CI(n51831), .I0(n3066), .I1(n858), .CO(n51832));
    SB_LUT4 add_2653_2_lut (.I0(n59283), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2653_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2653_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51831));
    SB_LUT4 add_2652_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n51830), 
            .O(n7937[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2652_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n51829), 
            .O(n7937[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_21 (.CI(n51829), .I0(n2939), .I1(n3084), .CO(n51830));
    SB_LUT4 add_2652_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n51828), 
            .O(n7937[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_20 (.CI(n51828), .I0(n2940), .I1(n2977), .CO(n51829));
    SB_LUT4 add_2652_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n51827), 
            .O(n7937[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_19 (.CI(n51827), .I0(n2941), .I1(n2867), .CO(n51828));
    SB_LUT4 add_2652_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n51826), 
            .O(n7937[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_18 (.CI(n51826), .I0(n2942), .I1(n2754), .CO(n51827));
    SB_LUT4 add_2652_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n51825), 
            .O(n7937[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_17 (.CI(n51825), .I0(n2943), .I1(n2638), .CO(n51826));
    SB_LUT4 add_2652_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n51824), 
            .O(n7937[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_16 (.CI(n51824), .I0(n2944), .I1(n2519), .CO(n51825));
    SB_LUT4 add_2652_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n51823), 
            .O(n7937[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_15 (.CI(n51823), .I0(n2945), .I1(n2397), .CO(n51824));
    SB_LUT4 add_2652_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n51822), 
            .O(n7937[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_14 (.CI(n51822), .I0(n2946), .I1(n2272), .CO(n51823));
    SB_LUT4 add_2652_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n51821), 
            .O(n7937[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_13 (.CI(n51821), .I0(n2947), .I1(n2144), .CO(n51822));
    SB_LUT4 add_2652_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n51820), 
            .O(n7937[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_12 (.CI(n51820), .I0(n2948), .I1(n2013), .CO(n51821));
    SB_LUT4 add_2652_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n51819), 
            .O(n7937[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_11 (.CI(n51819), .I0(n2949), .I1(n1879), .CO(n51820));
    SB_LUT4 add_2652_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n51818), 
            .O(n7937[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_10 (.CI(n51818), .I0(n2950), .I1(n1742), .CO(n51819));
    SB_LUT4 add_2652_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n51817), 
            .O(n7937[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_9 (.CI(n51817), .I0(n2951), .I1(n1602), .CO(n51818));
    SB_LUT4 add_2652_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n51816), 
            .O(n7937[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_8 (.CI(n51816), .I0(n2952), .I1(n1459), .CO(n51817));
    SB_LUT4 add_2652_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n51815), 
            .O(n7937[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_7 (.CI(n51815), .I0(n2953), .I1(n1460), .CO(n51816));
    SB_LUT4 add_2652_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n51814), 
            .O(n7937[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_6 (.CI(n51814), .I0(n2954), .I1(n1011), .CO(n51815));
    SB_LUT4 add_2652_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n51813), 
            .O(n7937[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_5 (.CI(n51813), .I0(n2955), .I1(n856), .CO(n51814));
    SB_LUT4 add_2652_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n51812), 
            .O(n7937[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_4 (.CI(n51812), .I0(n2956), .I1(n698), .CO(n51813));
    SB_LUT4 add_2652_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n51811), 
            .O(n7937[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2652_3 (.CI(n51811), .I0(n2957), .I1(n858), .CO(n51812));
    SB_LUT4 add_2652_2_lut (.I0(n59287), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2652_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i45602_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n62609));
    defparam i45602_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2652_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51811));
    SB_LUT4 i45712_4_lut (.I0(n62609), .I1(n61848), .I2(n61906), .I3(baudrate[9]), 
            .O(n62719));
    defparam i45712_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45705_1_lut (.I0(n62711), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59337));
    defparam i45705_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2651_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n51785), 
            .O(n7911[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2651_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n51784), 
            .O(n7911[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_20 (.CI(n51784), .I0(n2828), .I1(n2977), .CO(n51785));
    SB_LUT4 add_2651_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n51783), 
            .O(n7911[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_19 (.CI(n51783), .I0(n2829), .I1(n2867), .CO(n51784));
    SB_LUT4 add_2651_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n51782), 
            .O(n7911[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_18 (.CI(n51782), .I0(n2830), .I1(n2754), .CO(n51783));
    SB_LUT4 add_2651_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n51781), 
            .O(n7911[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_17 (.CI(n51781), .I0(n2831), .I1(n2638), .CO(n51782));
    SB_LUT4 add_2651_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n51780), 
            .O(n7911[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_16 (.CI(n51780), .I0(n2832), .I1(n2519), .CO(n51781));
    SB_LUT4 add_2651_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n51779), 
            .O(n7911[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_15 (.CI(n51779), .I0(n2833), .I1(n2397), .CO(n51780));
    SB_LUT4 add_2651_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n51778), 
            .O(n7911[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_14 (.CI(n51778), .I0(n2834), .I1(n2272), .CO(n51779));
    SB_LUT4 add_2651_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n51777), 
            .O(n7911[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_13 (.CI(n51777), .I0(n2835), .I1(n2144), .CO(n51778));
    SB_LUT4 add_2651_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n51776), 
            .O(n7911[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_12 (.CI(n51776), .I0(n2836), .I1(n2013), .CO(n51777));
    SB_LUT4 add_2651_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n51775), 
            .O(n7911[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_11 (.CI(n51775), .I0(n2837), .I1(n1879), .CO(n51776));
    SB_LUT4 add_2651_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n51774), 
            .O(n7911[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_10 (.CI(n51774), .I0(n2838), .I1(n1742), .CO(n51775));
    SB_LUT4 add_2651_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n51773), 
            .O(n7911[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_9 (.CI(n51773), .I0(n2839), .I1(n1602), .CO(n51774));
    SB_LUT4 add_2651_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n51772), 
            .O(n7911[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_8 (.CI(n51772), .I0(n2840), .I1(n1459), .CO(n51773));
    SB_LUT4 add_2651_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n51771), 
            .O(n7911[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_7 (.CI(n51771), .I0(n2841), .I1(n1460), .CO(n51772));
    SB_LUT4 add_2651_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n51770), 
            .O(n7911[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_6 (.CI(n51770), .I0(n2842), .I1(n1011), .CO(n51771));
    SB_LUT4 add_2651_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n51769), 
            .O(n7911[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_5 (.CI(n51769), .I0(n2843), .I1(n856), .CO(n51770));
    SB_LUT4 add_2651_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n51768), 
            .O(n7911[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_4 (.CI(n51768), .I0(n2844), .I1(n698), .CO(n51769));
    SB_LUT4 add_2651_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n51767), 
            .O(n7911[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2651_3 (.CI(n51767), .I0(n2845), .I1(n858), .CO(n51768));
    SB_LUT4 add_2651_2_lut (.I0(n59291), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n61174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2651_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2651_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n51767));
    SB_LUT4 i51523_2_lut (.I0(n48_adj_5083), .I1(n25166), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i51523_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2154_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2154_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n57762), .O(n61270));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61270), .O(n61276));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(n61276), .I1(n6), .I2(\r_SM_Main[1] ), 
            .I3(n27), .O(n28645));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'h0323;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n61498));
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'h0100;
    SB_LUT4 i2147_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2147_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45660_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n62667));
    defparam i45660_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1047 (.I0(n59034), .I1(n61498), .I2(n62100), 
            .I3(baudrate[16]), .O(n61526));
    defparam i1_4_lut_adj_1047.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1048 (.I0(n4), .I1(\r_SM_Main[1] ), .I2(n6), 
            .I3(\r_Bit_Index[0] ), .O(n61556));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1048.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4891), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61556), .O(n61562));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1050 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61562), .O(n61568));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'hfffe;
    SB_LUT4 i45730_4_lut (.I0(n62667), .I1(n62593), .I2(n62597), .I3(n62500), 
            .O(n62737));
    defparam i45730_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_965_i34_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61158), .I3(n48_adj_5048), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1051 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n61918));
    defparam i1_2_lut_4_lut_adj_1051.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1052 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n61916));
    defparam i1_2_lut_4_lut_adj_1052.LUT_INIT = 16'hfffe;
    SB_LUT4 i51372_4_lut (.I0(n62719), .I1(n65777), .I2(n62737), .I3(n61526), 
            .O(n68388));
    defparam i51372_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_i535_4_lut (.I0(n68388), .I1(n44_adj_5096), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 i6059_4_lut (.I0(n960), .I1(n9463), .I2(n21487), .I3(baudrate[3]), 
            .O(n21489));   // verilog/uart_rx.v(119[33:55])
    defparam i6059_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 i4107_2_lut (.I0(baudrate[3]), .I1(n42_adj_5052), .I2(GND_net), 
            .I3(GND_net), .O(n9470));   // verilog/uart_rx.v(119[33:55])
    defparam i4107_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3938_2_lut (.I0(n21475), .I1(n9299), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam i3938_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5097), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i51529_2_lut (.I0(n48_adj_5098), .I1(n25172), .I2(GND_net), 
            .I3(GND_net), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i51529_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i3945_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n9299), .I3(n21475), 
            .O(n46_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam i3945_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i639_4_lut (.I0(n58994), .I1(n294[19]), .I2(n46_adj_5099), 
            .I3(baudrate[4]), .O(n58996));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 i4116_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n9470), .I3(n21489), 
            .O(n46_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam i4116_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i742_4_lut (.I0(n58996), .I1(n294[18]), .I2(n46_adj_5100), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 i1_2_lut_4_lut_adj_1053 (.I0(n67358), .I1(baudrate[16]), .I2(n2476), 
            .I3(n61168), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1053.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n61908));
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n61910));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n61996), .I1(n61992), .I2(n61994), 
            .I3(n61990), .O(n61976));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i51443_2_lut_4_lut (.I0(n67358), .I1(baudrate[16]), .I2(n2476), 
            .I3(n62516), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i51443_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_1057 (.I0(n62102), .I1(n61936), .I2(n61988), 
            .I3(n61926), .O(n25218));
    defparam i1_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i49398_2_lut (.I0(n57790), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n65409));
    defparam i49398_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23365_rep_5_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59340));   // verilog/uart_rx.v(119[33:55])
    defparam i23365_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49390_4_lut (.I0(n65409), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n65406));
    defparam i49390_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n59340), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48739_4_lut (.I0(n65406), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n65403));
    defparam i48739_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i50765_3_lut (.I0(n42_adj_5101), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n67781));   // verilog/uart_rx.v(119[33:55])
    defparam i50765_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51515_4_lut (.I0(\r_SM_Main[2] ), .I1(n65403), .I2(r_SM_Main_2__N_3446[1]), 
            .I3(\r_SM_Main[1] ), .O(n28713));
    defparam i51515_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(n57790), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n61234));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'h1000;
    SB_LUT4 i50766_3_lut (.I0(n67781), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n67782));   // verilog/uart_rx.v(119[33:55])
    defparam i50766_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n67782), .I1(baudrate[5]), 
            .I2(n58996), .I3(GND_net), .O(n48_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_3_lut_4_lut_adj_1059 (.I0(n25163), .I1(n48_adj_5076), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5096));
    defparam i1_3_lut_4_lut_adj_1059.LUT_INIT = 16'hefff;
    SB_LUT4 i1_4_lut_adj_1060 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n61234), .O(n61240));
    defparam i1_4_lut_adj_1060.LUT_INIT = 16'h0100;
    SB_LUT4 i51399_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n61240), .O(n27409));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51399_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n61918), .I1(n25218), .I2(n61976), 
            .I3(n61916), .O(n25172));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'hfffe;
    SB_LUT4 i48761_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5076), .I2(n25163), 
            .I3(GND_net), .O(n65777));   // verilog/uart_rx.v(119[33:55])
    defparam i48761_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5103), .I1(baudrate[4]), 
            .I2(n43_adj_5089), .I3(GND_net), .O(n42_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51008_4_lut (.I0(n42_adj_5104), .I1(n38_adj_5102), .I2(n43_adj_5089), 
            .I3(n66027), .O(n68024));   // verilog/uart_rx.v(119[33:55])
    defparam i51008_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51009_3_lut (.I0(n68024), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n68025));   // verilog/uart_rx.v(119[33:55])
    defparam i51009_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1062 (.I0(n25172), .I1(n48_adj_5098), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1062.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7573[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7599[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7599[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1063 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n61848));
    defparam i1_2_lut_4_lut_adj_1063.LUT_INIT = 16'hfffe;
    SB_LUT4 i50759_3_lut (.I0(n34), .I1(baudrate[5]), .I2(n41_adj_5087), 
            .I3(GND_net), .O(n67775));   // verilog/uart_rx.v(119[33:55])
    defparam i50759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50760_3_lut (.I0(n67775), .I1(baudrate[6]), .I2(n43_adj_5053), 
            .I3(GND_net), .O(n67776));   // verilog/uart_rx.v(119[33:55])
    defparam i50760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49134_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4891), .I3(\o_Rx_DV_N_3488[8] ), .O(n65514));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49134_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i49245_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n57790), 
            .I3(r_SM_Main[0]), .O(n65520));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49245_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i49129_4_lut (.I0(n65514), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65511));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49129_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49892_4_lut (.I0(n43_adj_5053), .I1(n41_adj_5087), .I2(n39_adj_5061), 
            .I3(n66007), .O(n66908));
    defparam i49892_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49137_4_lut (.I0(n65520), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65517));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49137_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n65517), .I1(n65511), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_5051));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5105), .I1(baudrate[4]), 
            .I2(n39_adj_5061), .I3(GND_net), .O(n38_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49693_3_lut (.I0(n67776), .I1(baudrate[7]), .I2(n45_adj_5049), 
            .I3(GND_net), .O(n66709));   // verilog/uart_rx.v(119[33:55])
    defparam i49693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1064 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4894), 
            .I3(\r_SM_Main[0] ), .O(n61682));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1064.LUT_INIT = 16'hfeff;
    SB_LUT4 i50670_4_lut (.I0(n66709), .I1(n38_adj_5106), .I2(n45_adj_5049), 
            .I3(n66908), .O(n67686));   // verilog/uart_rx.v(119[33:55])
    defparam i50670_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1065 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n61682), .O(n59805));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 i48969_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n65985));   // verilog/uart_rx.v(119[33:55])
    defparam i48969_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1066 (.I0(n68327), .I1(baudrate[19]), .I2(n2827), 
            .I3(n61174), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1066.LUT_INIT = 16'h7100;
    SB_LUT4 i51504_2_lut_4_lut (.I0(n68327), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25212), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i51504_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50671_3_lut (.I0(n67686), .I1(baudrate[8]), .I2(n1408), .I3(GND_net), 
            .O(n48_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam i50671_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i42310_1_lut_4_lut (.I0(n62104), .I1(n62106), .I2(n61944), 
            .I3(n62102), .O(n59279));
    defparam i42310_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(n61158), .I1(n48_adj_5048), .I2(GND_net), 
            .I3(GND_net), .O(n1415));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7625[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n61702));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n61706));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n61708));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'heeee;
    SB_LUT4 i45676_4_lut (.I0(n61708), .I1(n61704), .I2(n61706), .I3(n61702), 
            .O(n62683));
    defparam i45676_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50757_3_lut (.I0(n32_adj_5095), .I1(baudrate[5]), .I2(n39_adj_5043), 
            .I3(GND_net), .O(n67773));   // verilog/uart_rx.v(119[33:55])
    defparam i50757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45650_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n62657));
    defparam i45650_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i45706_4_lut (.I0(n62657), .I1(n61988), .I2(n62655), .I3(n61942), 
            .O(n62713));
    defparam i45706_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45736_4_lut (.I0(n62713), .I1(n62593), .I2(n59034), .I3(baudrate[4]), 
            .O(n62743));
    defparam i45736_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51541_4_lut (.I0(n62683), .I1(n62500), .I2(n62743), .I3(n62498), 
            .O(n62747));
    defparam i51541_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i50758_3_lut (.I0(n67773), .I1(baudrate[6]), .I2(n41_adj_5042), 
            .I3(GND_net), .O(n67774));   // verilog/uart_rx.v(119[33:55])
    defparam i50758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49886_4_lut (.I0(n41_adj_5042), .I1(n39_adj_5043), .I2(n37_adj_5041), 
            .I3(n65999), .O(n66902));
    defparam i49886_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50672_3_lut (.I0(n34_adj_5109), .I1(baudrate[4]), .I2(n37_adj_5041), 
            .I3(GND_net), .O(n67688));   // verilog/uart_rx.v(119[33:55])
    defparam i50672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51520_3_lut (.I0(n25163), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25117));   // verilog/uart_rx.v(119[33:55])
    defparam i51520_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i49695_3_lut (.I0(n67774), .I1(baudrate[7]), .I2(n43_adj_5040), 
            .I3(GND_net), .O(n66711));   // verilog/uart_rx.v(119[33:55])
    defparam i49695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50755_4_lut (.I0(n66711), .I1(n67688), .I2(n43_adj_5040), 
            .I3(n66902), .O(n67771));   // verilog/uart_rx.v(119[33:55])
    defparam i50755_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50756_3_lut (.I0(n67771), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n67772));   // verilog/uart_rx.v(119[33:55])
    defparam i50756_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n67772), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1071 (.I0(n68353), .I1(baudrate[20]), .I2(n2938), 
            .I3(n61176), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1071.LUT_INIT = 16'h7100;
    SB_LUT4 i1_3_lut_adj_1072 (.I0(n62689), .I1(n48_adj_5110), .I2(n7651[14]), 
            .I3(GND_net), .O(n1702));
    defparam i1_3_lut_adj_1072.LUT_INIT = 16'h1010;
    SB_LUT4 i51507_2_lut_4_lut (.I0(n68353), .I1(baudrate[20]), .I2(n2938), 
            .I3(n62713), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i51507_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1073 (.I0(n67796), .I1(baudrate[21]), .I2(n3046), 
            .I3(n61178), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1073.LUT_INIT = 16'h7100;
    SB_LUT4 i51510_2_lut_4_lut (.I0(n67796), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25218), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i51510_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n7677[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48954_4_lut (.I0(n35_adj_5037), .I1(n33_adj_5033), .I2(n31_adj_5028), 
            .I3(n29_adj_5111), .O(n65970));
    defparam i48954_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n7989[20]), .I3(n294[1]), .O(n41_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n7989[19]), .I3(n294[1]), .O(n39_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32), .I1(baudrate[9]), 
            .I2(n43_adj_5012), .I3(GND_net), .O(n40_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n7989[16]), .I3(n294[1]), .O(n33_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n7989[17]), .I3(n294[1]), .O(n35_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n7989[18]), .I3(n294[1]), .O(n37_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i51420_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n62516), .I2(n48_adj_5072), 
            .I3(baudrate[15]), .O(n294[9]));
    defparam i51420_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n7989[14]), .I3(n294[1]), .O(n29_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n7989[15]), .I3(n294[1]), .O(n31_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i50749_3_lut (.I0(n28_adj_5115), .I1(baudrate[5]), .I2(n35_adj_5037), 
            .I3(GND_net), .O(n67765));   // verilog/uart_rx.v(119[33:55])
    defparam i50749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n7989[11]), .I3(n294[1]), .O(n23_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i50750_3_lut (.I0(n67765), .I1(baudrate[6]), .I2(n37_adj_5006), 
            .I3(GND_net), .O(n67766));   // verilog/uart_rx.v(119[33:55])
    defparam i50750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n7989[12]), .I3(n294[1]), .O(n25_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n7989[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n7989[22]), .I3(n294[1]), .O(n45_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n7989[21]), .I3(n294[1]), .O(n43_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i48941_4_lut (.I0(n41_adj_5039), .I1(n39_adj_5125), .I2(n37_adj_5006), 
            .I3(n65970), .O(n65957));
    defparam i48941_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n7989[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i45652_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n62516), .I2(n61704), 
            .I3(baudrate[15]), .O(n62659));
    defparam i45652_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51006_4_lut (.I0(n40_adj_5114), .I1(n30_adj_5094), .I2(n43_adj_5012), 
            .I3(n65952), .O(n68022));   // verilog/uart_rx.v(119[33:55])
    defparam i51006_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n7989[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n7989[7]), .I3(n294[1]), .O(n15_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i49701_3_lut (.I0(n67766), .I1(baudrate[7]), .I2(n39_adj_5125), 
            .I3(GND_net), .O(n66717));   // verilog/uart_rx.v(119[33:55])
    defparam i49701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51306_4_lut (.I0(n66717), .I1(n68022), .I2(n43_adj_5012), 
            .I3(n65957), .O(n68322));   // verilog/uart_rx.v(119[33:55])
    defparam i51306_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51307_3_lut (.I0(n68322), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n68323));   // verilog/uart_rx.v(119[33:55])
    defparam i51307_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n7989[13]), .I3(n294[1]), .O(n27_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i51236_3_lut (.I0(n68323), .I1(baudrate[11]), .I2(n1831), 
            .I3(GND_net), .O(n48_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam i51236_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n7989[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_3_lut_adj_1074 (.I0(n25185), .I1(n48_adj_5128), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1074.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n7989[9]), .I3(n294[1]), .O(n19_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n7989[10]), .I3(n294[1]), .O(n21_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n7703[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n7989[8]), .I3(n294[1]), .O(n17_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i49159_4_lut (.I0(n27_adj_5127), .I1(n15_adj_5126), .I2(n13), 
            .I3(n11), .O(n66175));
    defparam i49159_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n61704));
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'heeee;
    SB_LUT4 i49175_4_lut (.I0(n21_adj_5130), .I1(n19_adj_5129), .I2(n17_adj_5131), 
            .I3(n9), .O(n66191));
    defparam i49175_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5124), .I3(GND_net), .O(n16_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48921_4_lut (.I0(n33_adj_5134), .I1(n31_adj_5135), .I2(n29_adj_5136), 
            .I3(n27_adj_5133), .O(n65937));
    defparam i48921_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49101_2_lut (.I0(n43_adj_5124), .I1(n19_adj_5129), .I2(GND_net), 
            .I3(GND_net), .O(n66117));
    defparam i49101_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5131), .I3(GND_net), .O(n8_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5132), .I1(baudrate[22]), 
            .I2(n45_adj_5123), .I3(GND_net), .O(n24_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n7989[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49193_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n66209));
    defparam i49193_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i50056_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n66209), 
            .O(n67072));
    defparam i50056_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50048_4_lut (.I0(n19_adj_5129), .I1(n17_adj_5131), .I2(n15_adj_5126), 
            .I3(n67072), .O(n67064));
    defparam i50048_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51062_4_lut (.I0(n25_adj_5122), .I1(n23_adj_5121), .I2(n21_adj_5130), 
            .I3(n67064), .O(n68078));
    defparam i51062_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50483_4_lut (.I0(n31_adj_5120), .I1(n29_adj_5119), .I2(n27_adj_5127), 
            .I3(n68078), .O(n67499));
    defparam i50483_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51193_4_lut (.I0(n37_adj_5118), .I1(n35_adj_5117), .I2(n33_adj_5116), 
            .I3(n67499), .O(n68209));
    defparam i51193_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5093), .I1(baudrate[9]), 
            .I2(n41_adj_5139), .I3(GND_net), .O(n38_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5116), .I3(GND_net), .O(n12_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n61180), .I3(n48_adj_5142), .O(n4_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i50658_3_lut (.I0(n4_adj_5143), .I1(baudrate[13]), .I2(n27_adj_5127), 
            .I3(GND_net), .O(n67674));   // verilog/uart_rx.v(119[33:55])
    defparam i50658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50659_3_lut (.I0(n67674), .I1(baudrate[14]), .I2(n29_adj_5119), 
            .I3(GND_net), .O(n67675));   // verilog/uart_rx.v(119[33:55])
    defparam i50659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50747_3_lut (.I0(n26_adj_5091), .I1(baudrate[5]), .I2(n33_adj_5134), 
            .I3(GND_net), .O(n67763));   // verilog/uart_rx.v(119[33:55])
    defparam i50747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49138_2_lut (.I0(n33_adj_5116), .I1(n15_adj_5126), .I2(GND_net), 
            .I3(GND_net), .O(n66154));
    defparam i49138_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50748_3_lut (.I0(n67763), .I1(baudrate[6]), .I2(n35_adj_5144), 
            .I3(GND_net), .O(n67764));   // verilog/uart_rx.v(119[33:55])
    defparam i50748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48917_4_lut (.I0(n39_adj_5145), .I1(n37_adj_5146), .I2(n35_adj_5144), 
            .I3(n65937), .O(n65933));
    defparam i48917_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45679_1_lut_2_lut (.I0(baudrate[12]), .I1(n62659), .I2(GND_net), 
            .I3(GND_net), .O(n59320));
    defparam i45679_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i51414_2_lut_3_lut (.I0(baudrate[12]), .I1(n62659), .I2(n48_adj_5090), 
            .I3(GND_net), .O(n294[12]));
    defparam i51414_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_5141), .I1(baudrate[17]), 
            .I2(n35_adj_5117), .I3(GND_net), .O(n30_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51167_4_lut (.I0(n38_adj_5140), .I1(n28_adj_5092), .I2(n41_adj_5139), 
            .I3(n65931), .O(n68183));   // verilog/uart_rx.v(119[33:55])
    defparam i51167_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49144_4_lut (.I0(n33_adj_5116), .I1(n31_adj_5120), .I2(n29_adj_5119), 
            .I3(n66175), .O(n66160));
    defparam i49144_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51042_4_lut (.I0(n30_adj_5148), .I1(n10_adj_5147), .I2(n35_adj_5117), 
            .I3(n66154), .O(n68058));   // verilog/uart_rx.v(119[33:55])
    defparam i51042_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49763_3_lut (.I0(n67675), .I1(baudrate[15]), .I2(n31_adj_5120), 
            .I3(GND_net), .O(n66779));   // verilog/uart_rx.v(119[33:55])
    defparam i49763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51266_4_lut (.I0(n66779), .I1(n68058), .I2(n35_adj_5117), 
            .I3(n66160), .O(n68282));   // verilog/uart_rx.v(119[33:55])
    defparam i51266_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51267_3_lut (.I0(n68282), .I1(baudrate[18]), .I2(n37_adj_5118), 
            .I3(GND_net), .O(n68283));   // verilog/uart_rx.v(119[33:55])
    defparam i51267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50660_3_lut (.I0(n6_adj_5149), .I1(baudrate[10]), .I2(n21_adj_5130), 
            .I3(GND_net), .O(n67676));   // verilog/uart_rx.v(119[33:55])
    defparam i50660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50661_3_lut (.I0(n67676), .I1(baudrate[11]), .I2(n23_adj_5121), 
            .I3(GND_net), .O(n67677));   // verilog/uart_rx.v(119[33:55])
    defparam i50661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49703_3_lut (.I0(n67764), .I1(baudrate[7]), .I2(n37_adj_5146), 
            .I3(GND_net), .O(n66719));   // verilog/uart_rx.v(119[33:55])
    defparam i49703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51298_4_lut (.I0(n66719), .I1(n68183), .I2(n41_adj_5139), 
            .I3(n65933), .O(n68314));   // verilog/uart_rx.v(119[33:55])
    defparam i51298_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48983_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n65999));   // verilog/uart_rx.v(119[33:55])
    defparam i48983_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49109_4_lut (.I0(n43_adj_5124), .I1(n25_adj_5122), .I2(n23_adj_5121), 
            .I3(n66191), .O(n66125));
    defparam i49109_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50713_4_lut (.I0(n24_adj_5138), .I1(n8_adj_5137), .I2(n45_adj_5123), 
            .I3(n66117), .O(n67729));   // verilog/uart_rx.v(119[33:55])
    defparam i50713_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49761_3_lut (.I0(n67677), .I1(baudrate[12]), .I2(n25_adj_5122), 
            .I3(GND_net), .O(n66777));   // verilog/uart_rx.v(119[33:55])
    defparam i49761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51220_3_lut (.I0(n68283), .I1(baudrate[19]), .I2(n39_adj_5113), 
            .I3(GND_net), .O(n68236));   // verilog/uart_rx.v(119[33:55])
    defparam i51220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49111_4_lut (.I0(n43_adj_5124), .I1(n41_adj_5112), .I2(n39_adj_5113), 
            .I3(n68209), .O(n66127));
    defparam i49111_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i45701_1_lut_2_lut (.I0(baudrate[9]), .I1(n62689), .I2(GND_net), 
            .I3(GND_net), .O(n59329));
    defparam i45701_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i51145_4_lut (.I0(n66777), .I1(n67729), .I2(n45_adj_5123), 
            .I3(n66125), .O(n68161));   // verilog/uart_rx.v(119[33:55])
    defparam i51145_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49769_3_lut (.I0(n68236), .I1(baudrate[20]), .I2(n41_adj_5112), 
            .I3(GND_net), .O(n66785));   // verilog/uart_rx.v(119[33:55])
    defparam i49769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51299_3_lut (.I0(n68314), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n68315));   // verilog/uart_rx.v(119[33:55])
    defparam i51299_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51405_2_lut_3_lut_4_lut (.I0(baudrate[9]), .I1(n62689), .I2(n48_adj_5048), 
            .I3(baudrate[8]), .O(n294[16]));
    defparam i51405_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_3_lut_4_lut_adj_1076 (.I0(\r_Bit_Index[0] ), .I1(\r_SM_Main[1] ), 
            .I2(\r_SM_Main[2] ), .I3(r_SM_Main[0]), .O(n61572));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_4_lut_adj_1076.LUT_INIT = 16'hfff7;
    SB_LUT4 i3936_2_lut_4_lut (.I0(baudrate[2]), .I1(n805), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n9299));   // verilog/uart_rx.v(119[33:55])
    defparam i3936_2_lut_4_lut.LUT_INIT = 16'h0445;
    SB_LUT4 i51408_2_lut_3_lut (.I0(baudrate[9]), .I1(n62689), .I2(n48_adj_5044), 
            .I3(GND_net), .O(n294[15]));
    defparam i51408_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i45704_2_lut_3_lut_4_lut (.I0(baudrate[9]), .I1(n62689), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n62711));
    defparam i45704_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45703_1_lut_2_lut_3_lut (.I0(baudrate[9]), .I1(n62689), .I2(baudrate[8]), 
            .I3(GND_net), .O(n59333));
    defparam i45703_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n61114));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n7989[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51147_4_lut (.I0(n66785), .I1(n68161), .I2(n45_adj_5123), 
            .I3(n66127), .O(n68163));   // verilog/uart_rx.v(119[33:55])
    defparam i51147_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1078 (.I0(n62100), .I1(n61946), .I2(n61114), 
            .I3(n61944), .O(n61122));
    defparam i1_4_lut_adj_1078.LUT_INIT = 16'hfffe;
    SB_LUT4 i51547_4_lut (.I0(n61122), .I1(n68163), .I2(baudrate[23]), 
            .I3(n3253), .O(n60086));   // verilog/uart_rx.v(119[33:55])
    defparam i51547_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n7963[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51246_3_lut (.I0(n68315), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n68262));   // verilog/uart_rx.v(119[33:55])
    defparam i51246_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49709_3_lut (.I0(n68262), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam i49709_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45586_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n62593));
    defparam i45586_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45590_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n62597));
    defparam i45590_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i48991_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n66007));   // verilog/uart_rx.v(119[33:55])
    defparam i48991_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n7963[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1079 (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[1] ), .I3(\r_Bit_Index[0] ), .O(n61608));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_4_lut_adj_1079.LUT_INIT = 16'hffef;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n7963[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n7963[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49291_2_lut_3_lut (.I0(n25163), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n65498));   // verilog/uart_rx.v(119[33:55])
    defparam i49291_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_4_lut_adj_1080 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n62004));
    defparam i1_2_lut_4_lut_adj_1080.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1081 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n62002));
    defparam i1_2_lut_4_lut_adj_1081.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n7963[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n7963[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n7963[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48763_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5083), .I2(n25166), 
            .I3(GND_net), .O(n65779));   // verilog/uart_rx.v(119[33:55])
    defparam i48763_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51402_2_lut_4_lut (.I0(n68025), .I1(baudrate[6]), .I2(n1111), 
            .I3(n62711), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i51402_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n7963[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1082 (.I0(n68025), .I1(baudrate[6]), .I2(n1111), 
            .I3(n61156), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1082.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n7963[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n7703[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n7963[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n7963[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n7729[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n7963[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n7963[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n7963[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n7963[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n7729[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n7963[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n7963[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n7963[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n7963[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n7963[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n7963[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49412_3_lut_4_lut (.I0(n962), .I1(baudrate[1]), .I2(n48_adj_5098), 
            .I3(n25172), .O(n1115));
    defparam i49412_3_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n7729[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n62102));
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n62104));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1085 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n62100));
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(n62104), .I1(n62106), .I2(n61944), 
            .I3(n62102), .O(n25221));
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'hfffe;
    SB_LUT4 i49235_4_lut (.I0(n29_adj_5168), .I1(n17_adj_5166), .I2(n15_adj_5165), 
            .I3(n13_adj_5164), .O(n66251));
    defparam i49235_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50128_4_lut (.I0(n11_adj_5161), .I1(n9_adj_5159), .I2(n3171), 
            .I3(baudrate[2]), .O(n67144));
    defparam i50128_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50537_4_lut (.I0(n17_adj_5166), .I1(n15_adj_5165), .I2(n13_adj_5164), 
            .I3(n67144), .O(n67553));
    defparam i50537_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48904_4_lut (.I0(n33_adj_5167), .I1(n31_adj_5162), .I2(n29_adj_5160), 
            .I3(n27_adj_5169), .O(n65920));
    defparam i48904_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50533_4_lut (.I0(n23_adj_5158), .I1(n21_adj_5157), .I2(n19_adj_5163), 
            .I3(n67553), .O(n67549));
    defparam i50533_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49251_4_lut (.I0(n29_adj_5168), .I1(n27_adj_5156), .I2(n25_adj_5155), 
            .I3(n67549), .O(n66267));
    defparam i49251_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50666_3_lut (.I0(n6_adj_5170), .I1(baudrate[13]), .I2(n29_adj_5168), 
            .I3(GND_net), .O(n67682));   // verilog/uart_rx.v(119[33:55])
    defparam i50666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5084), .I1(baudrate[17]), 
            .I2(n37_adj_5153), .I3(GND_net), .O(n32_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50667_3_lut (.I0(n67682), .I1(baudrate[14]), .I2(n31_adj_5152), 
            .I3(GND_net), .O(n67683));   // verilog/uart_rx.v(119[33:55])
    defparam i50667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49229_4_lut (.I0(n35_adj_5154), .I1(n33_adj_5151), .I2(n31_adj_5152), 
            .I3(n66251), .O(n66245));
    defparam i49229_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51010_4_lut (.I0(n32_adj_5171), .I1(n12_adj_5082), .I2(n37_adj_5153), 
            .I3(n66243), .O(n68026));   // verilog/uart_rx.v(119[33:55])
    defparam i51010_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49749_3_lut (.I0(n67683), .I1(baudrate[15]), .I2(n33_adj_5151), 
            .I3(GND_net), .O(n66765));   // verilog/uart_rx.v(119[33:55])
    defparam i49749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50715_3_lut (.I0(n8_adj_5081), .I1(baudrate[10]), .I2(n23_adj_5158), 
            .I3(GND_net), .O(n67731));   // verilog/uart_rx.v(119[33:55])
    defparam i50715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50716_3_lut (.I0(n67731), .I1(baudrate[11]), .I2(n25_adj_5155), 
            .I3(GND_net), .O(n67732));   // verilog/uart_rx.v(119[33:55])
    defparam i50716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1087 (.I0(n57762), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main[1] ), .O(n61280));
    defparam i1_3_lut_4_lut_adj_1087.LUT_INIT = 16'hfdfc;
    SB_LUT4 i50110_4_lut (.I0(n25_adj_5155), .I1(n23_adj_5158), .I2(n21_adj_5157), 
            .I3(n66298), .O(n67126));
    defparam i50110_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50711_3_lut (.I0(n10_adj_5085), .I1(baudrate[9]), .I2(n21_adj_5157), 
            .I3(GND_net), .O(n67727));   // verilog/uart_rx.v(119[33:55])
    defparam i50711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49747_3_lut (.I0(n67732), .I1(baudrate[12]), .I2(n27_adj_5156), 
            .I3(GND_net), .O(n66763));   // verilog/uart_rx.v(119[33:55])
    defparam i49747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50885_4_lut (.I0(n35_adj_5154), .I1(n33_adj_5151), .I2(n31_adj_5152), 
            .I3(n66267), .O(n67901));
    defparam i50885_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30), .I1(baudrate[10]), 
            .I2(n41_adj_5172), .I3(GND_net), .O(n38_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51230_4_lut (.I0(n66765), .I1(n68026), .I2(n37_adj_5153), 
            .I3(n66245), .O(n68246));   // verilog/uart_rx.v(119[33:55])
    defparam i51230_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50953_4_lut (.I0(n66763), .I1(n67727), .I2(n27_adj_5156), 
            .I3(n67126), .O(n67969));   // verilog/uart_rx.v(119[33:55])
    defparam i50953_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51334_4_lut (.I0(n67969), .I1(n68246), .I2(n37_adj_5153), 
            .I3(n67901), .O(n68350));   // verilog/uart_rx.v(119[33:55])
    defparam i51334_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i23432_rep_3_2_lut (.I0(n7729[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n59314));   // verilog/uart_rx.v(119[33:55])
    defparam i23432_rep_3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51583_2_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(\r_SM_Main[2] ), .I3(r_SM_Main[0]), .O(n27292));
    defparam i51583_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i51335_3_lut (.I0(n68350), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n68351));   // verilog/uart_rx.v(119[33:55])
    defparam i51335_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n59314), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51223_3_lut (.I0(n68351), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n68239));   // verilog/uart_rx.v(119[33:55])
    defparam i51223_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50743_3_lut (.I0(n26_adj_5174), .I1(baudrate[6]), .I2(n33_adj_5167), 
            .I3(GND_net), .O(n67759));   // verilog/uart_rx.v(119[33:55])
    defparam i50743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51138_3_lut (.I0(n68239), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n68154));   // verilog/uart_rx.v(119[33:55])
    defparam i51138_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51139_3_lut (.I0(n68154), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n68155));   // verilog/uart_rx.v(119[33:55])
    defparam i51139_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50744_3_lut (.I0(n67759), .I1(baudrate[7]), .I2(n35_adj_5175), 
            .I3(GND_net), .O(n67760));   // verilog/uart_rx.v(119[33:55])
    defparam i50744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49759_3_lut (.I0(n68155), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam i49759_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n7937[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42330_1_lut (.I0(n25206), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59299));
    defparam i42330_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n7937[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n7937[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48894_4_lut (.I0(n39_adj_5176), .I1(n37_adj_5177), .I2(n35_adj_5175), 
            .I3(n65920), .O(n65910));
    defparam i48894_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n7937[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n7937[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n7937[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n7937[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51014_4_lut (.I0(n38_adj_5173), .I1(n28_adj_5080), .I2(n41_adj_5172), 
            .I3(n65904), .O(n68030));   // verilog/uart_rx.v(119[33:55])
    defparam i51014_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n7937[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n7937[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n7937[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n7937[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n7937[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n7937[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n7937[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n7937[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49711_3_lut (.I0(n67760), .I1(baudrate[8]), .I2(n37_adj_5177), 
            .I3(GND_net), .O(n66727));   // verilog/uart_rx.v(119[33:55])
    defparam i49711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51300_4_lut (.I0(n66727), .I1(n68030), .I2(n41_adj_5172), 
            .I3(n65910), .O(n68316));   // verilog/uart_rx.v(119[33:55])
    defparam i51300_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n7937[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n7937[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51301_3_lut (.I0(n68316), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n68317));   // verilog/uart_rx.v(119[33:55])
    defparam i51301_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n7937[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51244_3_lut (.I0(n68317), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n68260));   // verilog/uart_rx.v(119[33:55])
    defparam i51244_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n7937[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n7937[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49717_3_lut (.I0(n68260), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam i49717_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49351_4_lut (.I0(n31_adj_5193), .I1(n19_adj_5192), .I2(n17_adj_5191), 
            .I3(n15_adj_5189), .O(n66367));
    defparam i49351_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1088 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n61998));
    defparam i1_4_lut_adj_1088.LUT_INIT = 16'hfffe;
    SB_LUT4 i50208_4_lut (.I0(n13_adj_5187), .I1(n11_adj_5186), .I2(n3065), 
            .I3(baudrate[2]), .O(n67224));
    defparam i50208_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50575_4_lut (.I0(n19_adj_5192), .I1(n17_adj_5191), .I2(n15_adj_5189), 
            .I3(n67224), .O(n67591));
    defparam i50575_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50571_4_lut (.I0(n25_adj_5185), .I1(n23_adj_5184), .I2(n21_adj_5188), 
            .I3(n67591), .O(n67587));
    defparam i50571_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49353_4_lut (.I0(n31_adj_5193), .I1(n29_adj_5183), .I2(n27_adj_5182), 
            .I3(n67587), .O(n66369));
    defparam i49353_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_3_lut_adj_1089 (.I0(n61948), .I1(n61996), .I2(n61730), 
            .I3(GND_net), .O(n62006));
    defparam i1_3_lut_adj_1089.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(n62006), .I1(n62002), .I2(n62004), 
            .I3(n61998), .O(n25194));
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1091 (.I0(n25194), .I1(n48_adj_5190), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1091.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n7781[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50723_3_lut (.I0(n8_adj_5194), .I1(baudrate[13]), .I2(n31_adj_5193), 
            .I3(GND_net), .O(n67739));   // verilog/uart_rx.v(119[33:55])
    defparam i50723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50724_3_lut (.I0(n67739), .I1(baudrate[14]), .I2(n33_adj_5180), 
            .I3(GND_net), .O(n67740));   // verilog/uart_rx.v(119[33:55])
    defparam i50724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5077), .I1(baudrate[17]), 
            .I2(n39_adj_5178), .I3(GND_net), .O(n34_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48841_4_lut (.I0(n27_adj_5197), .I1(n25_adj_5198), .I2(n23_adj_5199), 
            .I3(n21_adj_5195), .O(n65857));
    defparam i48841_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48836_4_lut (.I0(n33_adj_5200), .I1(n31_adj_5201), .I2(n29_adj_5202), 
            .I3(n65857), .O(n65852));
    defparam i48836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49335_4_lut (.I0(n37_adj_5181), .I1(n35_adj_5179), .I2(n33_adj_5180), 
            .I3(n66367), .O(n66351));
    defparam i49335_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50988_4_lut (.I0(n34_adj_5196), .I1(n14_adj_5075), .I2(n39_adj_5178), 
            .I3(n66346), .O(n68004));   // verilog/uart_rx.v(119[33:55])
    defparam i50988_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i42326_1_lut (.I0(n25209), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n59295));
    defparam i42326_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49739_3_lut (.I0(n67740), .I1(baudrate[15]), .I2(n35_adj_5179), 
            .I3(GND_net), .O(n66755));   // verilog/uart_rx.v(119[33:55])
    defparam i49739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50725_3_lut (.I0(n10), .I1(baudrate[10]), .I2(n25_adj_5185), 
            .I3(GND_net), .O(n67741));   // verilog/uart_rx.v(119[33:55])
    defparam i50725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50726_3_lut (.I0(n67741), .I1(baudrate[11]), .I2(n27_adj_5182), 
            .I3(GND_net), .O(n67742));   // verilog/uart_rx.v(119[33:55])
    defparam i50726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50184_4_lut (.I0(n27_adj_5182), .I1(n25_adj_5185), .I2(n23_adj_5184), 
            .I3(n66402), .O(n67200));
    defparam i50184_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5078), .I1(baudrate[9]), 
            .I2(n23_adj_5184), .I3(GND_net), .O(n20_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49737_3_lut (.I0(n67742), .I1(baudrate[12]), .I2(n29_adj_5183), 
            .I3(GND_net), .O(n66753));   // verilog/uart_rx.v(119[33:55])
    defparam i49737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50897_4_lut (.I0(n37_adj_5181), .I1(n35_adj_5179), .I2(n33_adj_5180), 
            .I3(n66369), .O(n67913));
    defparam i50897_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51304_4_lut (.I0(n66755), .I1(n68004), .I2(n39_adj_5178), 
            .I3(n66351), .O(n68320));   // verilog/uart_rx.v(119[33:55])
    defparam i51304_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50707_4_lut (.I0(n66753), .I1(n20_adj_5203), .I2(n29_adj_5183), 
            .I3(n67200), .O(n67723));   // verilog/uart_rx.v(119[33:55])
    defparam i50707_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51332_4_lut (.I0(n67723), .I1(n68320), .I2(n39_adj_5178), 
            .I3(n67913), .O(n68348));   // verilog/uart_rx.v(119[33:55])
    defparam i51332_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51333_3_lut (.I0(n68348), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n68349));   // verilog/uart_rx.v(119[33:55])
    defparam i51333_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50779_3_lut (.I0(n68349), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n67795));   // verilog/uart_rx.v(119[33:55])
    defparam i50779_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50780_3_lut (.I0(n67795), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n67796));   // verilog/uart_rx.v(119[33:55])
    defparam i50780_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n7859[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4102_2_lut_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), 
            .I3(baudrate[1]), .O(n42_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam i4102_2_lut_4_lut.LUT_INIT = 16'hb2bb;
    SB_LUT4 i4100_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9463));   // verilog/uart_rx.v(119[33:55])
    defparam i4100_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i3931_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam i3931_2_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n7859[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5074), .I1(baudrate[7]), 
            .I2(n31_adj_5201), .I3(GND_net), .O(n28_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6047_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n21473));   // verilog/uart_rx.v(119[33:55])
    defparam i6047_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n7911[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n7859[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n7911[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n7911[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n7911[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n7911[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n7911[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n7911[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n7859[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n7911[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n7859[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n7859[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n7859[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5071), .I1(baudrate[9]), 
            .I2(n35_adj_5208), .I3(GND_net), .O(n32_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51228_4_lut (.I0(n32_adj_5209), .I1(n22_adj_5069), .I2(n35_adj_5208), 
            .I3(n65847), .O(n68244));   // verilog/uart_rx.v(119[33:55])
    defparam i51228_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n7859[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n7911[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51229_3_lut (.I0(n68244), .I1(baudrate[10]), .I2(n37_adj_5211), 
            .I3(GND_net), .O(n68245));   // verilog/uart_rx.v(119[33:55])
    defparam i51229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n7859[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n7911[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51227_3_lut (.I0(n68245), .I1(baudrate[11]), .I2(n39_adj_5213), 
            .I3(GND_net), .O(n68243));   // verilog/uart_rx.v(119[33:55])
    defparam i51227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50717_4_lut (.I0(n39_adj_5213), .I1(n37_adj_5211), .I2(n35_adj_5208), 
            .I3(n65852), .O(n67733));
    defparam i50717_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n7859[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n7911[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51169_4_lut (.I0(n28_adj_5204), .I1(n20_adj_5073), .I2(n31_adj_5201), 
            .I3(n65854), .O(n68185));   // verilog/uart_rx.v(119[33:55])
    defparam i51169_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n7859[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51141_3_lut (.I0(n68243), .I1(baudrate[12]), .I2(n41_adj_5215), 
            .I3(GND_net), .O(n40_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam i51141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51241_4_lut (.I0(n40_adj_5216), .I1(n68185), .I2(n41_adj_5215), 
            .I3(n67733), .O(n68257));   // verilog/uart_rx.v(119[33:55])
    defparam i51241_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n7911[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n7911[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51242_3_lut (.I0(n68257), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n68258));   // verilog/uart_rx.v(119[33:55])
    defparam i51242_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n7859[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1092 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n61608), .I3(GND_net), .O(n61610));
    defparam i1_2_lut_3_lut_adj_1092.LUT_INIT = 16'hf7f7;
    SB_LUT4 i51182_3_lut (.I0(n68258), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n68198));   // verilog/uart_rx.v(119[33:55])
    defparam i51182_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n7859[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n7859[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1093 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n61572), .I3(GND_net), .O(n61538));
    defparam i1_2_lut_3_lut_adj_1093.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n7911[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n7911[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n7911[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n7859[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51411_2_lut_4_lut (.I0(n67772), .I1(baudrate[9]), .I2(n1552), 
            .I3(n62689), .O(n294[14]));
    defparam i51411_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n7859[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n7833[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n7911[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n7833[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49011_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n66027));   // verilog/uart_rx.v(119[33:55])
    defparam i49011_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n7911[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50968_3_lut (.I0(n68198), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i50968_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n7911[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n7833[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n7833[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n7781[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n7833[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49450_4_lut (.I0(n33_adj_5225), .I1(n21_adj_5224), .I2(n19_adj_5223), 
            .I3(n17_adj_5222), .O(n66466));
    defparam i49450_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49499_4_lut (.I0(n15_adj_5221), .I1(n13_adj_5220), .I2(n2956), 
            .I3(baudrate[2]), .O(n66515));
    defparam i49499_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n7833[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n7833[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n7833[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50266_4_lut (.I0(n21_adj_5224), .I1(n19_adj_5223), .I2(n17_adj_5222), 
            .I3(n66515), .O(n67282));
    defparam i50266_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n7807[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50260_4_lut (.I0(n27_adj_5219), .I1(n25_adj_5218), .I2(n23_adj_5217), 
            .I3(n67282), .O(n67276));
    defparam i50260_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49452_4_lut (.I0(n33_adj_5225), .I1(n31_adj_5214), .I2(n29_adj_5212), 
            .I3(n67276), .O(n66468));
    defparam i49452_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n7833[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n7833[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5017));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5016));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50731_3_lut (.I0(n10_adj_5226), .I1(baudrate[13]), .I2(n33_adj_5225), 
            .I3(GND_net), .O(n67747));   // verilog/uart_rx.v(119[33:55])
    defparam i50731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n7833[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n7833[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50732_3_lut (.I0(n67747), .I1(baudrate[14]), .I2(n35_adj_5207), 
            .I3(GND_net), .O(n67748));   // verilog/uart_rx.v(119[33:55])
    defparam i50732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n7833[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n7833[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5015));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n7807[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5068), .I1(baudrate[17]), 
            .I2(n41_adj_5206), .I3(GND_net), .O(n36_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n7807[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49442_4_lut (.I0(n39_adj_5210), .I1(n37_adj_5205), .I2(n35_adj_5207), 
            .I3(n66466), .O(n66458));
    defparam i49442_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n7807[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n7807[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n7807[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50986_4_lut (.I0(n36_adj_5229), .I1(n16_adj_5067), .I2(n41_adj_5206), 
            .I3(n66456), .O(n68002));   // verilog/uart_rx.v(119[33:55])
    defparam i50986_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49727_3_lut (.I0(n67748), .I1(baudrate[15]), .I2(n37_adj_5205), 
            .I3(GND_net), .O(n66743));   // verilog/uart_rx.v(119[33:55])
    defparam i49727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n7807[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5066), .I1(baudrate[9]), 
            .I2(n25_adj_5218), .I3(GND_net), .O(n22_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n7807[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n7807[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n7807[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51179_4_lut (.I0(n22_adj_5233), .I1(n12), .I2(n25_adj_5218), 
            .I3(n65594), .O(n68195));   // verilog/uart_rx.v(119[33:55])
    defparam i51179_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51180_3_lut (.I0(n68195), .I1(baudrate[10]), .I2(n27_adj_5219), 
            .I3(GND_net), .O(n68196));   // verilog/uart_rx.v(119[33:55])
    defparam i51180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50993_3_lut (.I0(n68196), .I1(baudrate[11]), .I2(n29_adj_5212), 
            .I3(GND_net), .O(n68009));   // verilog/uart_rx.v(119[33:55])
    defparam i50993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50911_4_lut (.I0(n39_adj_5210), .I1(n37_adj_5205), .I2(n35_adj_5207), 
            .I3(n66468), .O(n67927));
    defparam i50911_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n7807[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n7807[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51302_4_lut (.I0(n66743), .I1(n68002), .I2(n41_adj_5206), 
            .I3(n66458), .O(n68318));   // verilog/uart_rx.v(119[33:55])
    defparam i51302_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49725_3_lut (.I0(n68009), .I1(baudrate[12]), .I2(n31_adj_5214), 
            .I3(GND_net), .O(n66741));   // verilog/uart_rx.v(119[33:55])
    defparam i49725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n7807[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n7807[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51338_4_lut (.I0(n66741), .I1(n68318), .I2(n41_adj_5206), 
            .I3(n67927), .O(n68354));   // verilog/uart_rx.v(119[33:55])
    defparam i51338_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51339_3_lut (.I0(n68354), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n68355));   // verilog/uart_rx.v(119[33:55])
    defparam i51339_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51337_3_lut (.I0(n68355), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n68353));   // verilog/uart_rx.v(119[33:55])
    defparam i51337_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n7807[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n7781[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n7781[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1094 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n61608), .I3(GND_net), .O(n61628));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1094.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1095 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n61572), .I3(GND_net), .O(n61574));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1095.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_3_lut_4_lut_adj_1096 (.I0(n61712), .I1(n62711), .I2(baudrate[0]), 
            .I3(n48_adj_5065), .O(n962));
    defparam i1_3_lut_4_lut_adj_1096.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n7781[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n7781[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1097 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n61608), .I3(GND_net), .O(n61592));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1097.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n7885[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n7781[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n7885[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n7885[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n7885[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1098 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n61572), .I3(GND_net), .O(n61646));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1098.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n7885[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n7781[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48713_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n65729));
    defparam i48713_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n7781[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n7755[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45512_2_lut (.I0(baudrate[17]), .I1(n25206), .I2(GND_net), 
            .I3(GND_net), .O(n62516));
    defparam i45512_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n7885[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n7885[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n7755[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n7755[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n7755[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n7755[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n7885[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n7885[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n7755[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n7755[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n7885[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n7885[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n7755[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n7885[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48880_4_lut (.I0(n29_adj_5253), .I1(n27_adj_5252), .I2(n25_adj_5251), 
            .I3(n23_adj_5258), .O(n65896));
    defparam i48880_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5259));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48871_4_lut (.I0(n35_adj_5257), .I1(n33_adj_5256), .I2(n31_adj_5254), 
            .I3(n65896), .O(n65887));
    defparam i48871_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5064), .I1(baudrate[7]), 
            .I2(n33_adj_5256), .I3(GND_net), .O(n30_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5063), .I1(baudrate[9]), 
            .I2(n37_adj_5250), .I3(GND_net), .O(n34_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50767_4_lut (.I0(n34_adj_5264), .I1(n24_adj_5062), .I2(n37_adj_5250), 
            .I3(n65882), .O(n67783));   // verilog/uart_rx.v(119[33:55])
    defparam i50767_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n7885[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48781_4_lut (.I0(n25_adj_5227), .I1(n23_adj_5240), .I2(n21_adj_5239), 
            .I3(n19_adj_5261), .O(n65797));
    defparam i48781_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n7885[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48775_4_lut (.I0(n31_adj_5238), .I1(n29_adj_5237), .I2(n27_adj_5228), 
            .I3(n65797), .O(n65791));
    defparam i48775_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50656_4_lut (.I0(n37_adj_5236), .I1(n35_adj_5235), .I2(n33_adj_5234), 
            .I3(n65791), .O(n67672));
    defparam i50656_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50799_3_lut (.I0(n18_adj_5060), .I1(baudrate[13]), .I2(n41_adj_5232), 
            .I3(GND_net), .O(n67815));   // verilog/uart_rx.v(119[33:55])
    defparam i50799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50768_3_lut (.I0(n67783), .I1(baudrate[10]), .I2(n39_adj_5246), 
            .I3(GND_net), .O(n67784));   // verilog/uart_rx.v(119[33:55])
    defparam i50768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50738_3_lut (.I0(n67784), .I1(baudrate[11]), .I2(n41_adj_5247), 
            .I3(GND_net), .O(n67754));   // verilog/uart_rx.v(119[33:55])
    defparam i50738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50733_4_lut (.I0(n41_adj_5247), .I1(n39_adj_5246), .I2(n37_adj_5250), 
            .I3(n65887), .O(n67749));
    defparam i50733_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n7885[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50800_3_lut (.I0(n67815), .I1(baudrate[14]), .I2(n43_adj_5231), 
            .I3(GND_net), .O(n67816));   // verilog/uart_rx.v(119[33:55])
    defparam i50800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50809_4_lut (.I0(n30_adj_5263), .I1(n22_adj_5262), .I2(n33_adj_5256), 
            .I3(n65893), .O(n67825));   // verilog/uart_rx.v(119[33:55])
    defparam i50809_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49721_3_lut (.I0(n67754), .I1(baudrate[12]), .I2(n43_adj_5245), 
            .I3(GND_net), .O(n66737));   // verilog/uart_rx.v(119[33:55])
    defparam i49721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51004_4_lut (.I0(n66737), .I1(n67825), .I2(n43_adj_5245), 
            .I3(n67749), .O(n68020));   // verilog/uart_rx.v(119[33:55])
    defparam i51004_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51005_3_lut (.I0(n68020), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n68021));   // verilog/uart_rx.v(119[33:55])
    defparam i51005_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50964_3_lut (.I0(n68021), .I1(baudrate[14]), .I2(n2227), 
            .I3(GND_net), .O(n48_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam i50964_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(n61164), .I1(n48_adj_5072), .I2(GND_net), 
            .I3(GND_net), .O(n2367));
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n7755[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n7885[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n7755[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n7781[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n7755[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n7781[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n7781[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n7885[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n7885[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1100 (.I0(n62659), .I1(n48_adj_5150), .I2(n7729[11]), 
            .I3(GND_net), .O(n2110));
    defparam i1_3_lut_adj_1100.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n7755[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49605_4_lut (.I0(n43_adj_5231), .I1(n41_adj_5232), .I2(n29_adj_5237), 
            .I3(n65795), .O(n66621));
    defparam i49605_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n7755[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n7781[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n7781[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48617_4_lut (.I0(n35_adj_5270), .I1(n23_adj_5269), .I2(n21_adj_5268), 
            .I3(n19_adj_5267), .O(n65633));
    defparam i48617_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49533_4_lut (.I0(n17_adj_5266), .I1(n15_adj_5265), .I2(n2844), 
            .I3(baudrate[2]), .O(n66549));
    defparam i49533_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24), .I1(baudrate[7]), 
            .I2(n29_adj_5237), .I3(GND_net), .O(n26_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n61730));
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'heeee;
    SB_LUT4 i50282_4_lut (.I0(n23_adj_5269), .I1(n21_adj_5268), .I2(n19_adj_5267), 
            .I3(n66549), .O(n67298));
    defparam i50282_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50280_4_lut (.I0(n29_adj_5260), .I1(n27_adj_5259), .I2(n25_adj_5255), 
            .I3(n67298), .O(n67296));
    defparam i50280_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48619_4_lut (.I0(n35_adj_5270), .I1(n33_adj_5249), .I2(n31_adj_5248), 
            .I3(n67296), .O(n65635));
    defparam i48619_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n7729[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n7729[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n7729[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n7729[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n7729[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50783_3_lut (.I0(n12_adj_5272), .I1(baudrate[13]), .I2(n35_adj_5270), 
            .I3(GND_net), .O(n67799));   // verilog/uart_rx.v(119[33:55])
    defparam i50783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n7729[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n7729[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50689_3_lut (.I0(n67816), .I1(baudrate[15]), .I2(n45), .I3(GND_net), 
            .O(n42_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam i50689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n7729[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5059), .I1(baudrate[17]), 
            .I2(n43_adj_5242), .I3(GND_net), .O(n38_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n7729[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n7703[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n7703[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n7703[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n7703[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50784_3_lut (.I0(n67799), .I1(baudrate[14]), .I2(n37_adj_5243), 
            .I3(GND_net), .O(n67800));   // verilog/uart_rx.v(119[33:55])
    defparam i50784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48611_4_lut (.I0(n41_adj_5244), .I1(n39_adj_5241), .I2(n37_adj_5243), 
            .I3(n65633), .O(n65627));
    defparam i48611_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50781_4_lut (.I0(n38_adj_5274), .I1(n18_adj_5057), .I2(n43_adj_5242), 
            .I3(n65625), .O(n67797));   // verilog/uart_rx.v(119[33:55])
    defparam i50781_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50704_3_lut (.I0(n67800), .I1(baudrate[15]), .I2(n39_adj_5241), 
            .I3(GND_net), .O(n67720));   // verilog/uart_rx.v(119[33:55])
    defparam i50704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48721_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n65737));
    defparam i48721_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n7703[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n61162), .I1(n48_adj_5090), .I2(GND_net), 
            .I3(GND_net), .O(n1977));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n7703[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n7703[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5056), .I1(baudrate[9]), 
            .I2(n27_adj_5259), .I3(GND_net), .O(n24_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51177_4_lut (.I0(n24_adj_5275), .I1(n14_adj_5055), .I2(n27_adj_5259), 
            .I3(n65643), .O(n68193));   // verilog/uart_rx.v(119[33:55])
    defparam i51177_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n7703[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n7703[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51178_3_lut (.I0(n68193), .I1(baudrate[10]), .I2(n29_adj_5260), 
            .I3(GND_net), .O(n68194));   // verilog/uart_rx.v(119[33:55])
    defparam i51178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50995_3_lut (.I0(n68194), .I1(baudrate[11]), .I2(n31_adj_5248), 
            .I3(GND_net), .O(n68011));   // verilog/uart_rx.v(119[33:55])
    defparam i50995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5058), .I1(baudrate[9]), 
            .I2(n33_adj_5234), .I3(GND_net), .O(n30_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50611_4_lut (.I0(n41_adj_5244), .I1(n39_adj_5241), .I2(n37_adj_5243), 
            .I3(n65635), .O(n67627));
    defparam i50611_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51149_4_lut (.I0(n67720), .I1(n67797), .I2(n43_adj_5242), 
            .I3(n65627), .O(n68165));   // verilog/uart_rx.v(119[33:55])
    defparam i51149_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50979_3_lut (.I0(n68011), .I1(baudrate[12]), .I2(n33_adj_5249), 
            .I3(GND_net), .O(n67995));   // verilog/uart_rx.v(119[33:55])
    defparam i50979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51310_4_lut (.I0(n67995), .I1(n68165), .I2(n43_adj_5242), 
            .I3(n67627), .O(n68326));   // verilog/uart_rx.v(119[33:55])
    defparam i51310_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51311_3_lut (.I0(n68326), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n68327));   // verilog/uart_rx.v(119[33:55])
    defparam i51311_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51171_4_lut (.I0(n30_adj_5276), .I1(n20_adj_5054), .I2(n33_adj_5234), 
            .I3(n65789), .O(n68187));   // verilog/uart_rx.v(119[33:55])
    defparam i51171_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48674_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n65690));
    defparam i48674_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1103 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n61148));
    defparam i1_3_lut_4_lut_adj_1103.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48643_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n65659));
    defparam i48643_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n61944));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'heeee;
    SB_LUT4 i51172_3_lut (.I0(n68187), .I1(baudrate[10]), .I2(n35_adj_5235), 
            .I3(GND_net), .O(n68188));   // verilog/uart_rx.v(119[33:55])
    defparam i51172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1105 (.I0(n61988), .I1(n61944), .I2(n61946), 
            .I3(baudrate[11]), .O(n61974));
    defparam i1_4_lut_adj_1105.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1106 (.I0(n61974), .I1(n61976), .I2(n61964), 
            .I3(n61904), .O(n25185));
    defparam i1_4_lut_adj_1106.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i23400_rep_4_2_lut (.I0(n7651[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n59323));   // verilog/uart_rx.v(119[33:55])
    defparam i23400_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n59323), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51001_3_lut (.I0(n68188), .I1(baudrate[11]), .I2(n37_adj_5236), 
            .I3(GND_net), .O(n68017));   // verilog/uart_rx.v(119[33:55])
    defparam i51001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49607_4_lut (.I0(n43_adj_5231), .I1(n41_adj_5232), .I2(n39_adj_5230), 
            .I3(n67672), .O(n66623));
    defparam i49607_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50753_3_lut (.I0(n32_adj_5281), .I1(baudrate[6]), .I2(n39_adj_5279), 
            .I3(GND_net), .O(n67769));   // verilog/uart_rx.v(119[33:55])
    defparam i50753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50340_4_lut (.I0(n42_adj_5273), .I1(n26_adj_5271), .I2(n45), 
            .I3(n66621), .O(n67356));   // verilog/uart_rx.v(119[33:55])
    defparam i50340_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50754_3_lut (.I0(n67769), .I1(baudrate[7]), .I2(n41_adj_5280), 
            .I3(GND_net), .O(n67770));   // verilog/uart_rx.v(119[33:55])
    defparam i50754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49874_4_lut (.I0(n41_adj_5280), .I1(n39_adj_5279), .I2(n37_adj_5278), 
            .I3(n65985), .O(n66890));
    defparam i49874_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50674_3_lut (.I0(n34_adj_5108), .I1(baudrate[5]), .I2(n37_adj_5278), 
            .I3(GND_net), .O(n67690));   // verilog/uart_rx.v(119[33:55])
    defparam i50674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49698_3_lut (.I0(n67770), .I1(baudrate[8]), .I2(n43_adj_5277), 
            .I3(GND_net), .O(n66714));   // verilog/uart_rx.v(119[33:55])
    defparam i49698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50751_4_lut (.I0(n66714), .I1(n67690), .I2(n43_adj_5277), 
            .I3(n66890), .O(n67767));   // verilog/uart_rx.v(119[33:55])
    defparam i50751_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50752_3_lut (.I0(n67767), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n67768));   // verilog/uart_rx.v(119[33:55])
    defparam i50752_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1107 (.I0(n67993), .I1(baudrate[18]), .I2(n2713), 
            .I3(n61172), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1107.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n67768), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50970_3_lut (.I0(n68017), .I1(baudrate[12]), .I2(n39_adj_5230), 
            .I3(GND_net), .O(n67986));   // verilog/uart_rx.v(119[33:55])
    defparam i50970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5007));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7651[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n7677[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51501_2_lut_4_lut (.I0(n67993), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25209), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i51501_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7651[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n7677[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7651[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n7677[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, enable_slow_N_4211, ready_prev, clk16MHz, n5753, 
            \state[2] , \state[0] , \state[1] , n58096, data, ID, 
            n25014, \state[0]_adj_3 , baudrate, n29123, n29122, n29121, 
            n29120, n29119, n29118, n29117, n29116, n39313, n29033, 
            rw, n57558, data_ready, n57286, n57342, n38869, \state_7__N_3916[0] , 
            n4, n25133, n60892, VCC_net, scl_enable, \state_7__N_4108[0] , 
            n6388, n29039, \saved_addr[0] , sda_enable, scl, n4_adj_4, 
            n29920, n29919, n29918, n29917, n29916, n29915, n29914, 
            n4_adj_5, n29647, n38965, n8, \state_7__N_4124[3] , n10, 
            n6, n38852, sda_out, n25136, n25119) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output enable_slow_N_4211;
    output ready_prev;
    input clk16MHz;
    output [0:0]n5753;
    output \state[2] ;
    output \state[0] ;
    output \state[1] ;
    output n58096;
    output [7:0]data;
    output [7:0]ID;
    output n25014;
    output \state[0]_adj_3 ;
    output [31:0]baudrate;
    input n29123;
    input n29122;
    input n29121;
    input n29120;
    input n29119;
    input n29118;
    input n29117;
    input n29116;
    output n39313;
    input n29033;
    output rw;
    input n57558;
    output data_ready;
    input n57286;
    input n57342;
    output n38869;
    input \state_7__N_3916[0] ;
    output n4;
    output n25133;
    output n60892;
    input VCC_net;
    output scl_enable;
    output \state_7__N_4108[0] ;
    output n6388;
    input n29039;
    output \saved_addr[0] ;
    output sda_enable;
    output scl;
    output n4_adj_4;
    input n29920;
    input n29919;
    input n29918;
    input n29917;
    input n29916;
    input n29915;
    input n29914;
    output n4_adj_5;
    input n29647;
    output n38965;
    input n8;
    input \state_7__N_4124[3] ;
    output n10;
    output n6;
    output n38852;
    output sda_out;
    output n25136;
    output n25119;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n4_c, enable, n52416, n59048;
    wire [15:0]delay_counter_15__N_3954;
    
    wire n27261;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n28717, n6_c, n58104, n4_adj_4996, n6642, n6644, n6645, 
        n6646, n6647, n6648, n29027, n29148, n29149, n29150, n14, 
        n13, n14_adj_4997, n15, n29151;
    wire [7:0]state_7__N_3883;
    
    wire n60689, n29152, n29153, n53272, n27551, n28952, n29154;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    wire [2:0]n17;
    
    wire n29147, n29146, n29145, n29144, n29143, n29142, n29141, 
        n29140, n29139, n29138, n29137, n29136, n29135, n29134, 
        n29133, n29132, n29131, n29130, n29129, n29128, n29127, 
        n29126, n29125, n29124;
    wire [15:0]n5040;
    
    wire n51421, n51420, n51419, n51418, n51417, n51416, n39114, 
        n51415, n51414, n51413, n51412, n51411, n51410, n51409, 
        n51408, n51407, n62537, n7, n4_adj_5001, n65588;
    
    SB_LUT4 equal_327_i4_2_lut (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));   // verilog/eeprom.v(66[9:28])
    defparam equal_327_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4211));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5753[0]), .R(\state[2] ));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i42080_2_lut (.I0(n52416), .I1(byte_counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n59048));
    defparam i42080_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27261), 
            .D(delay_counter_15__N_3954[1]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27261), 
            .D(delay_counter_15__N_3954[2]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27261), 
            .D(delay_counter_15__N_3954[3]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i4_4_lut (.I0(ready_prev), .I1(n58096), .I2(\state[2] ), .I3(n6_c), 
            .O(n52416));
    defparam i4_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_977 (.I0(byte_counter[0]), .I1(n52416), .I2(GND_net), 
            .I3(GND_net), .O(n58104));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_adj_977.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_329_i4_2_lut (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4996));   // verilog/eeprom.v(66[9:28])
    defparam equal_329_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27261), 
            .D(n6642), .S(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27261), 
            .D(delay_counter_15__N_3954[5]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27261), 
            .D(n6644), .S(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27261), 
            .D(n6645), .S(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27261), 
            .D(n6646), .S(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27261), 
            .D(n6647), .S(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27261), .D(n6648), .S(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13284_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[0]), 
            .I3(ID[0]), .O(n29027));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21969_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[7]), 
            .I3(ID[7]), .O(n29148));   // verilog/eeprom.v(35[8] 81[4])
    defparam i21969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27261), .D(delay_counter_15__N_3954[11]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27261), .D(delay_counter_15__N_3954[12]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27261), .D(delay_counter_15__N_3954[13]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27261), .D(delay_counter_15__N_3954[14]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13406_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[6]), 
            .I3(ID[6]), .O(n29149));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13407_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[5]), 
            .I3(ID[5]), .O(n29150));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut (.I0(delay_counter[7]), .I1(delay_counter[1]), .I2(delay_counter[3]), 
            .I3(delay_counter[15]), .O(n14));   // verilog/eeprom.v(55[12:28])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27261), .D(delay_counter_15__N_3954[15]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i5_4_lut (.I0(delay_counter[13]), .I1(delay_counter[11]), .I2(delay_counter[9]), 
            .I3(delay_counter[14]), .O(n13));   // verilog/eeprom.v(55[12:28])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_978 (.I0(delay_counter[6]), .I1(delay_counter[4]), 
            .I2(n13), .I3(n14), .O(n14_adj_4997));   // verilog/eeprom.v(55[12:28])
    defparam i5_4_lut_adj_978.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_979 (.I0(delay_counter[0]), .I1(delay_counter[8]), 
            .I2(delay_counter[5]), .I3(delay_counter[2]), .O(n15));   // verilog/eeprom.v(55[12:28])
    defparam i6_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(delay_counter[12]), .I2(n14_adj_4997), 
            .I3(delay_counter[10]), .O(n25014));   // verilog/eeprom.v(55[12:28])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1438_Mux_0_i3_4_lut (.I0(\state[0] ), .I1(enable_slow_N_4211), 
            .I2(\state[1] ), .I3(n25014), .O(n5753[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1438_Mux_0_i3_4_lut.LUT_INIT = 16'h0a4a;
    SB_LUT4 i13408_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[4]), 
            .I3(ID[4]), .O(n29151));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(n60689), .D(state_7__N_3883[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13409_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[3]), 
            .I3(ID[3]), .O(n29152));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13410_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[2]), 
            .I3(ID[2]), .O(n29153));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_counter_1938__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27551), .D(n53272), .R(n28952));   // verilog/eeprom.v(68[25:39])
    SB_LUT4 i13411_3_lut_4_lut (.I0(n4_adj_4996), .I1(n58104), .I2(data[1]), 
            .I3(ID[1]), .O(n29154));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0]_adj_3 ), .I1(state[3]), .I2(state[2]), 
            .I3(state[1]), .O(n58096));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35373_2_lut_3_lut_4_lut (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i35373_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_DFFESR byte_counter_1938__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27551), .D(n17[2]), .R(n28952));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1938__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27551), .D(n17[1]), .R(n28952));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n29154));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n29153));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n29152));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n29151));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n29150));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n29149));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n29148));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n29147));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n29146));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n29145));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n29144));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n29143));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n29142));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n29141));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n29140));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n29139));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n29138));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n29137));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n29136));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n29135));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n29134));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n29133));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n29132));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n29131));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n29130));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n29129));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n29128));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n29127));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n29126));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n29125));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n29124));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n29123));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n29122));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n29121));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n29120));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n29119));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n29118));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n29117));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n29116));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(n39313), .O(n28717));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1012;
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n29033));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n57558));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29027));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27261), 
            .D(delay_counter_15__N_3954[0]), .R(n28717));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13397_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[7]), 
            .I3(baudrate[7]), .O(n29140));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13397_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13398_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[6]), 
            .I3(baudrate[6]), .O(n29141));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13398_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13399_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[5]), 
            .I3(baudrate[5]), .O(n29142));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13399_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13400_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[4]), 
            .I3(baudrate[4]), .O(n29143));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13400_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF state_i2 (.Q(\state[2] ), .C(clk16MHz), .D(n57286));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i0 (.Q(\state[0] ), .C(clk16MHz), .D(n57342));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13401_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[3]), 
            .I3(baudrate[3]), .O(n29144));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13401_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i51396_3_lut_4_lut_4_lut (.I0(\state[2] ), .I1(n39313), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n27261));
    defparam i51396_3_lut_4_lut_4_lut.LUT_INIT = 16'h0552;
    SB_LUT4 i13402_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[2]), 
            .I3(baudrate[2]), .O(n29145));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13402_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13403_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[1]), 
            .I3(baudrate[1]), .O(n29146));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13403_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13404_3_lut_4_lut (.I0(n4_adj_4996), .I1(n59048), .I2(data[0]), 
            .I3(baudrate[0]), .O(n29147));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13404_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13389_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[7]), 
            .I3(baudrate[15]), .O(n29132));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13390_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[6]), 
            .I3(baudrate[14]), .O(n29133));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13391_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[5]), 
            .I3(baudrate[13]), .O(n29134));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i51377_2_lut (.I0(n25014), .I1(enable_slow_N_4211), .I2(GND_net), 
            .I3(GND_net), .O(n5040[1]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i51377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13392_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[4]), 
            .I3(baudrate[12]), .O(n29135));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13393_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[3]), 
            .I3(baudrate[11]), .O(n29136));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13394_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[2]), 
            .I3(baudrate[10]), .O(n29137));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_1087_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5040[1]), 
            .I3(n51421), .O(delay_counter_15__N_3954[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1087_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5040[1]), 
            .I3(n51420), .O(delay_counter_15__N_3954[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_16 (.CI(n51420), .I0(delay_counter[14]), .I1(n5040[1]), 
            .CO(n51421));
    SB_LUT4 add_1087_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5040[1]), 
            .I3(n51419), .O(delay_counter_15__N_3954[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_15 (.CI(n51419), .I0(delay_counter[13]), .I1(n5040[1]), 
            .CO(n51420));
    SB_LUT4 add_1087_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5040[1]), 
            .I3(n51418), .O(delay_counter_15__N_3954[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_14 (.CI(n51418), .I0(delay_counter[12]), .I1(n5040[1]), 
            .CO(n51419));
    SB_LUT4 add_1087_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5040[1]), 
            .I3(n51417), .O(delay_counter_15__N_3954[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_13 (.CI(n51417), .I0(delay_counter[11]), .I1(n5040[1]), 
            .CO(n51418));
    SB_LUT4 add_1087_12_lut (.I0(n39114), .I1(delay_counter[10]), .I2(n5040[1]), 
            .I3(n51416), .O(n6648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1087_12 (.CI(n51416), .I0(delay_counter[10]), .I1(n5040[1]), 
            .CO(n51417));
    SB_LUT4 add_1087_11_lut (.I0(n39114), .I1(delay_counter[9]), .I2(n5040[1]), 
            .I3(n51415), .O(n6647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1087_11 (.CI(n51415), .I0(delay_counter[9]), .I1(n5040[1]), 
            .CO(n51416));
    SB_LUT4 add_1087_10_lut (.I0(n39114), .I1(delay_counter[8]), .I2(n5040[1]), 
            .I3(n51414), .O(n6646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1087_10 (.CI(n51414), .I0(delay_counter[8]), .I1(n5040[1]), 
            .CO(n51415));
    SB_LUT4 add_1087_9_lut (.I0(n39114), .I1(delay_counter[7]), .I2(n5040[1]), 
            .I3(n51413), .O(n6645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1087_9 (.CI(n51413), .I0(delay_counter[7]), .I1(n5040[1]), 
            .CO(n51414));
    SB_LUT4 add_1087_8_lut (.I0(n39114), .I1(delay_counter[6]), .I2(n5040[1]), 
            .I3(n51412), .O(n6644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1087_8 (.CI(n51412), .I0(delay_counter[6]), .I1(n5040[1]), 
            .CO(n51413));
    SB_LUT4 add_1087_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5040[1]), 
            .I3(n51411), .O(delay_counter_15__N_3954[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_7 (.CI(n51411), .I0(delay_counter[5]), .I1(n5040[1]), 
            .CO(n51412));
    SB_LUT4 add_1087_6_lut (.I0(n39114), .I1(delay_counter[4]), .I2(n5040[1]), 
            .I3(n51410), .O(n6642)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1087_6 (.CI(n51410), .I0(delay_counter[4]), .I1(n5040[1]), 
            .CO(n51411));
    SB_LUT4 add_1087_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5040[1]), 
            .I3(n51409), .O(delay_counter_15__N_3954[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_5 (.CI(n51409), .I0(delay_counter[3]), .I1(n5040[1]), 
            .CO(n51410));
    SB_LUT4 add_1087_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5040[1]), 
            .I3(n51408), .O(delay_counter_15__N_3954[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_4 (.CI(n51408), .I0(delay_counter[2]), .I1(n5040[1]), 
            .CO(n51409));
    SB_LUT4 add_1087_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5040[1]), 
            .I3(n51407), .O(delay_counter_15__N_3954[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_3 (.CI(n51407), .I0(delay_counter[1]), .I1(n5040[1]), 
            .CO(n51408));
    SB_LUT4 add_1087_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5040[1]), 
            .I3(GND_net), .O(delay_counter_15__N_3954[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1087_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1087_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5040[1]), 
            .CO(n51407));
    SB_LUT4 i13395_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[1]), 
            .I3(baudrate[9]), .O(n29138));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13396_3_lut_4_lut (.I0(n4_c), .I1(n58104), .I2(data[0]), 
            .I3(baudrate[8]), .O(n29139));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i45530_2_lut_3_lut (.I0(\state[0]_adj_3 ), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n62537));
    defparam i45530_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable_slow_N_4211), .I1(ready_prev), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n53272));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i23223_2_lut (.I0(enable_slow_N_4211), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n38869));
    defparam i23223_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(55[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(\state_7__N_3916[0] ), 
            .I3(\state[0] ), .O(n4_adj_5001));
    defparam i1_4_lut.LUT_INIT = 16'hbbba;
    SB_LUT4 i49418_4_lut (.I0(n62537), .I1(n25014), .I2(\state[1] ), .I3(state[3]), 
            .O(n65588));
    defparam i49418_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n65588), .I1(n4_adj_5001), .I2(n38869), .I3(\state[0] ), 
            .O(n60689));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i6842_4_lut (.I0(\state[1] ), .I1(n39313), .I2(\state[2] ), 
            .I3(\state[0] ), .O(state_7__N_3883[1]));   // verilog/eeprom.v(38[3] 80[10])
    defparam i6842_4_lut.LUT_INIT = 16'ha5ba;
    SB_LUT4 i23468_1_lut_2_lut (.I0(\state[2] ), .I1(n39313), .I2(GND_net), 
            .I3(GND_net), .O(n39114));
    defparam i23468_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state[0]_adj_3 ), .I1(state[3]), 
            .I2(state[1]), .I3(state[2]), .O(n4));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_980 (.I0(\state_7__N_3916[0] ), .I1(\state[0] ), 
            .I2(\state[1] ), .I3(\state[2] ), .O(n28952));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut_adj_980.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state_7__N_3916[0] ), .I1(\state[0] ), 
            .I2(\state[1] ), .I3(\state[2] ), .O(n27551));   // verilog/eeprom.v(68[25:39])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h00c2;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n25133));   // verilog/eeprom.v(71[5:15])
    defparam i1_2_lut_adj_981.LUT_INIT = 16'heeee;
    SB_LUT4 i23664_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n39313));
    defparam i23664_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13381_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[7]), 
            .I3(baudrate[23]), .O(n29124));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13381_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13382_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[6]), 
            .I3(baudrate[22]), .O(n29125));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13382_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13383_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[5]), 
            .I3(baudrate[21]), .O(n29126));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13383_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13384_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[4]), 
            .I3(baudrate[20]), .O(n29127));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13384_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13385_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[3]), 
            .I3(baudrate[19]), .O(n29128));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13385_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i35380_3_lut_4_lut (.I0(n38869), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i35380_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i13386_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[2]), 
            .I3(baudrate[18]), .O(n29129));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13386_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13387_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[1]), 
            .I3(baudrate[17]), .O(n29130));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13387_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13388_3_lut_4_lut (.I0(n4_c), .I1(n59048), .I2(data[0]), 
            .I3(baudrate[16]), .O(n29131));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13388_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_982 (.I0(byte_counter[1]), .I1(byte_counter[0]), 
            .I2(n52416), .I3(byte_counter[2]), .O(n60892));   // verilog/eeprom.v(35[8] 81[4])
    defparam i2_3_lut_4_lut_adj_982.LUT_INIT = 16'hefff;
    i2c_controller i2c (.GND_net(GND_net), .VCC_net(VCC_net), .\state[0] (\state[0]_adj_3 ), 
            .\state[1] (state[1]), .\state[3] (state[3]), .\state[2] (state[2]), 
            .enable_slow_N_4211(enable_slow_N_4211), .clk16MHz(clk16MHz), 
            .scl_enable(scl_enable), .\state_7__N_4108[0] (\state_7__N_4108[0] ), 
            .n6388(n6388), .n29039(n29039), .\saved_addr[0] (\saved_addr[0] ), 
            .sda_enable(sda_enable), .scl(scl), .n4(n4_adj_4), .n29920(n29920), 
            .data({data}), .n29919(n29919), .n29918(n29918), .n29917(n29917), 
            .n29916(n29916), .n29915(n29915), .n29914(n29914), .n4_adj_2(n4_adj_5), 
            .n29647(n29647), .n38965(n38965), .n8(n8), .enable(enable), 
            .n7(n7), .\state_7__N_4124[3] (\state_7__N_4124[3] ), .n10(n10), 
            .n6(n6), .n38852(n38852), .sda_out(sda_out), .n25136(n25136), 
            .n25119(n25119)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (GND_net, VCC_net, \state[0] , \state[1] , \state[3] , 
            \state[2] , enable_slow_N_4211, clk16MHz, scl_enable, \state_7__N_4108[0] , 
            n6388, n29039, \saved_addr[0] , sda_enable, scl, n4, 
            n29920, data, n29919, n29918, n29917, n29916, n29915, 
            n29914, n4_adj_2, n29647, n38965, n8, enable, n7, 
            \state_7__N_4124[3] , n10, n6, n38852, sda_out, n25136, 
            n25119) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    output \state[0] ;
    output \state[1] ;
    output \state[3] ;
    output \state[2] ;
    output enable_slow_N_4211;
    input clk16MHz;
    output scl_enable;
    output \state_7__N_4108[0] ;
    output n6388;
    input n29039;
    output \saved_addr[0] ;
    output sda_enable;
    output scl;
    output n4;
    input n29920;
    output [7:0]data;
    input n29919;
    input n29918;
    input n29917;
    input n29916;
    input n29915;
    input n29914;
    output n4_adj_2;
    input n29647;
    output n38965;
    input n8;
    input enable;
    input n7;
    input \state_7__N_4124[3] ;
    output n10;
    output n6;
    output n38852;
    output sda_out;
    output n25136;
    output n25119;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n52187, n52186, n52185, n52184, n52183;
    wire [1:0]n6452;
    
    wire n60097, n15, n6719, i2c_clk_N_4197, scl_enable_N_4198, enable_slow_N_4210, 
        n27321, n10_c, n28716, n5, n39131, n39147, n39322, n60949, 
        n59974;
    wire [7:0]n119;
    
    wire n27306;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n28702, n60911, n27315, n57398, n27313, sda_out_adj_4986, 
        n11, n6381, n4_adj_4988, n65586, n11_adj_4989, n4_adj_4990, 
        n51428, n51427, n51426, n51425, n51424, n51423, n51422, 
        n9, n10_adj_4991, n12, n11_adj_4993, n11_adj_4994, state_7__N_4107, 
        n11_adj_4995, n28, n68386, n59054;
    
    SB_LUT4 counter2_1947_1948_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n52187), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1947_1948_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1947_1948_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n52186), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1947_1948_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1947_1948_add_4_6 (.CI(n52186), .I0(GND_net), .I1(counter2[4]), 
            .CO(n52187));
    SB_LUT4 counter2_1947_1948_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n52185), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1947_1948_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1947_1948_add_4_5 (.CI(n52185), .I0(GND_net), .I1(counter2[3]), 
            .CO(n52186));
    SB_LUT4 counter2_1947_1948_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n52184), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1947_1948_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1947_1948_add_4_4 (.CI(n52184), .I0(GND_net), .I1(counter2[2]), 
            .CO(n52185));
    SB_LUT4 counter2_1947_1948_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n52183), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1947_1948_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1947_1948_add_4_3 (.CI(n52183), .I0(GND_net), .I1(counter2[1]), 
            .CO(n52184));
    SB_LUT4 counter2_1947_1948_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1947_1948_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1947_1948_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n52183));
    SB_LUT4 i51454_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(enable_slow_N_4211));   // verilog/i2c_controller.v(44[32:47])
    defparam i51454_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6452[1]), 
            .I3(\state[1] ), .O(n60097));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 equal_280_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n15));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam equal_280_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n6719));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4197));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4198));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4108[0] ), .C(clk16MHz), .E(n27321), 
            .D(enable_slow_N_4210));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n28716));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n28716), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4197));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR counter2_1947_1948__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n28716));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6388), .D(n5), 
            .S(n39131));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6388), .D(n39147), 
            .S(n39322));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6388), .D(n60949), 
            .S(n59974));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27306), .D(n119[1]), 
            .S(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27306), .D(n119[2]), 
            .S(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27306), .D(n119[3]), 
            .R(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27306), .D(n119[4]), 
            .R(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27306), .D(n119[5]), 
            .R(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27306), .D(n119[6]), 
            .R(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27306), .D(n119[7]), 
            .R(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29039));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27315), 
            .D(n60911), .S(n57398));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4986), .C(i2c_clk), .E(n27313), 
            .D(n60097), .S(n57398));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27306), .D(n119[0]), 
            .S(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_1505_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));
    defparam equal_1505_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_3_lut_4_lut_adj_967 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n60911));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_967.LUT_INIT = 16'h1110;
    SB_LUT4 i23243_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i23243_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_359_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_359_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29920));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29919));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29918));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29917));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29916));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29915));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29914));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_357_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_357_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29647));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i23319_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n38965));
    defparam i23319_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_4108[0] ), .I2(enable_slow_N_4211), 
            .I3(GND_net), .O(n27321));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_DFFSR counter2_1947_1948__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n28716));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1947_1948__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n28716));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1947_1948__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n28716));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1947_1948__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n28716));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1947_1948__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n28716));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i1_2_lut_adj_968 (.I0(\state[3] ), .I1(n6381), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4988));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'hbbbb;
    SB_LUT4 i49394_4_lut (.I0(n7), .I1(n4_adj_4988), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n65586));
    defparam i49394_4_lut.LUT_INIT = 16'hfcdd;
    SB_LUT4 i14_4_lut (.I0(n65586), .I1(n15), .I2(n6719), .I3(\state_7__N_4124[3] ), 
            .O(n27306));
    defparam i14_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i1_4_lut (.I0(\state_7__N_4124[3] ), .I1(n11_adj_4989), .I2(n11), 
            .I3(enable), .O(n4_adj_4990));
    defparam i1_4_lut.LUT_INIT = 16'h2a2f;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n51428), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n51427), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n51427), .I0(counter[6]), .I1(VCC_net), 
            .CO(n51428));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n51426), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n51426), .I0(counter[5]), .I1(VCC_net), 
            .CO(n51427));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n51425), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n51425), .I0(counter[4]), .I1(VCC_net), 
            .CO(n51426));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n51424), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n51424), .I0(counter[3]), .I1(VCC_net), 
            .CO(n51425));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n51423), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n51423), .I0(counter[2]), .I1(VCC_net), 
            .CO(n51424));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n51422), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n51422), .I0(counter[1]), .I1(VCC_net), 
            .CO(n51423));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n51422));
    SB_LUT4 i51556_2_lut (.I0(\state_7__N_4124[3] ), .I1(n11_adj_4989), 
            .I2(GND_net), .I3(GND_net), .O(n39147));
    defparam i51556_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_139_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_139_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_141_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4991));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_141_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6381));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_969 (.I0(n11_adj_4993), .I1(n11_adj_4994), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut_adj_969.LUT_INIT = 16'h8888;
    SB_LUT4 i51553_4_lut (.I0(n6388), .I1(\state[0] ), .I2(n11_adj_4993), 
            .I3(n7), .O(n39131));
    defparam i51553_4_lut.LUT_INIT = 16'h0a8a;
    SB_LUT4 i51386_4_lut (.I0(state_7__N_4107), .I1(n6381), .I2(n11_adj_4993), 
            .I3(n38852), .O(n6388));
    defparam i51386_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_970 (.I0(n11_adj_4995), .I1(n11_adj_4989), .I2(\state_7__N_4124[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_970.LUT_INIT = 16'h5755;
    SB_LUT4 i23550_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n38852));
    defparam i23550_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i51550_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6388), .O(n59974));
    defparam i51550_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i12964_2_lut_4_lut (.I0(n27306), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n28702));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i12964_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i2418_2_lut (.I0(sda_out_adj_4986), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51426_2_lut (.I0(\state_7__N_4108[0] ), .I1(enable_slow_N_4211), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4210));   // verilog/i2c_controller.v(62[6:32])
    defparam i51426_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4995));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut_adj_971 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut_adj_971.LUT_INIT = 16'h5110;
    SB_LUT4 i51370_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n68386));
    defparam i51370_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_972 (.I0(n11), .I1(n68386), .I2(n28), .I3(n59054), 
            .O(n27313));
    defparam i1_4_lut_adj_972.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1722_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6452[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1722_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i42086_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n59054));
    defparam i42086_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[0] ), .I1(n7), .I2(\state[3] ), .I3(n11), 
            .O(n57398));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_973 (.I0(n11), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n59054), .O(n27315));
    defparam i1_4_lut_adj_973.LUT_INIT = 16'h0a22;
    SB_LUT4 i23656_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_4107));
    defparam i23656_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n11_adj_4989));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_adj_974 (.I0(n9), .I1(n10_adj_4991), .I2(counter[0]), 
            .I3(GND_net), .O(n25136));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_974.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_975 (.I0(n9), .I1(n10_adj_4991), .I2(counter[0]), 
            .I3(GND_net), .O(n25119));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_975.LUT_INIT = 16'hefef;
    SB_LUT4 i51552_3_lut_4_lut (.I0(n9), .I1(n10_adj_4991), .I2(n11_adj_4994), 
            .I3(n6388), .O(n39322));   // verilog/i2c_controller.v(151[5:14])
    defparam i51552_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n11_adj_4994));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_976 (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_adj_4990), 
            .I3(n9), .O(n60949));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut_adj_976.LUT_INIT = 16'hf0f4;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4993));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i23651_3_lut_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(scl_enable_N_4198));   // verilog/i2c_controller.v(44[32:47])
    defparam i23651_3_lut_4_lut_4_lut.LUT_INIT = 16'hfefc;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_setpoint, GND_net, n39, n3014, pwm_out, clk32MHz, 
            \pwm_counter[19] , reset, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input [23:0]pwm_setpoint;
    input GND_net;
    input n39;
    input n3014;
    output pwm_out;
    input clk32MHz;
    output \pwm_counter[19] ;
    input reset;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n41, n45, n43, n37, n23, n25, n29, n31, n35, n9, 
        n17, n19, n21, n33, n11, n13, n15, n27, n66224, n66181, 
        n12, n30, n66296, n67130, n67102, n68086, n67503, n68207, 
        n6, n67861, n67862, n16, n24, n66111, n8, n66108, n67642, 
        n66604, n4, n67863, n67864, n66158, n10, n66141, n68171, 
        n66600, n68308, n68309, n68273, n66115, n68134, n67645, 
        n68231, pwm_out_N_577, n56754, n52023, n48, n56776, n52022, 
        n56796, n52021, n56816, n52020, n56838, n52019, n56860, 
        n52018, n56888, n52017, n56910, n52016, n56952, n52015, 
        n56992, n52014, n57610, n57024, n52013, n57058, n52012, 
        n57102, n52011, n57144, n52010, n57174, n52009, n57206, 
        n52008, n57242, n52007, n57284, n52006, n57368, n52005, 
        n57528, n52004, n57626, n52003, n57624, n52002, n57622, 
        n52001, n60886, n22, n15_adj_4983, n20, n24_adj_4984, n19_adj_4985;
    
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49208_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n66224));
    defparam i49208_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49165_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n66181));
    defparam i49165_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50114_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n66296), 
            .O(n67130));
    defparam i50114_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50086_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n67130), 
            .O(n67102));
    defparam i50086_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51070_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n67102), 
            .O(n68086));
    defparam i51070_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50487_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n68086), 
            .O(n67503));
    defparam i50487_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51191_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67503), 
            .O(n68207));
    defparam i51191_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50845_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n67861));   // verilog/pwm.v(21[8:24])
    defparam i50845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50846_3_lut (.I0(n67861), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n67862));   // verilog/pwm.v(21[8:24])
    defparam i50846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49095_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n66224), 
            .O(n66111));
    defparam i49095_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50626_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n66108), 
            .O(n67642));   // verilog/pwm.v(21[8:24])
    defparam i50626_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49588_3_lut (.I0(n67862), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n66604));   // verilog/pwm.v(21[8:24])
    defparam i49588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50847_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n67863));   // verilog/pwm.v(21[8:24])
    defparam i50847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50848_3_lut (.I0(n67863), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n67864));   // verilog/pwm.v(21[8:24])
    defparam i50848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49142_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n66181), 
            .O(n66158));
    defparam i49142_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51155_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n66141), 
            .O(n68171));   // verilog/pwm.v(21[8:24])
    defparam i51155_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49584_3_lut (.I0(n67864), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n66600));   // verilog/pwm.v(21[8:24])
    defparam i49584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51292_4_lut (.I0(n66600), .I1(n68171), .I2(n35), .I3(n66158), 
            .O(n68308));   // verilog/pwm.v(21[8:24])
    defparam i51292_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51293_3_lut (.I0(n68308), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n68309));   // verilog/pwm.v(21[8:24])
    defparam i51293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51257_3_lut (.I0(n68309), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n68273));   // verilog/pwm.v(21[8:24])
    defparam i51257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49099_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n68207), 
            .O(n66115));
    defparam i49099_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51118_4_lut (.I0(n66604), .I1(n67642), .I2(n45), .I3(n66111), 
            .O(n68134));   // verilog/pwm.v(21[8:24])
    defparam i51118_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50629_3_lut (.I0(n68273), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n67645));   // verilog/pwm.v(21[8:24])
    defparam i50629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51215_4_lut (.I0(n67645), .I1(n68134), .I2(n45), .I3(n66115), 
            .O(n68231));   // verilog/pwm.v(21[8:24])
    defparam i51215_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51216_3_lut (.I0(n68231), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i51216_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n3014), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_1931_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n52023), .O(n56754)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1931_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n52022), .O(n56776)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_24 (.CI(n52022), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n52023));
    SB_LUT4 pwm_counter_1931_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n52021), .O(n56796)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_23 (.CI(n52021), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n52022));
    SB_LUT4 pwm_counter_1931_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n52020), .O(n56816)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_22 (.CI(n52020), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n52021));
    SB_LUT4 pwm_counter_1931_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[19] ), 
            .I3(n52019), .O(n56838)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_21 (.CI(n52019), .I0(GND_net), .I1(\pwm_counter[19] ), 
            .CO(n52020));
    SB_LUT4 pwm_counter_1931_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n52018), .O(n56860)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_20 (.CI(n52018), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n52019));
    SB_LUT4 pwm_counter_1931_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n52017), .O(n56888)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_19 (.CI(n52017), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n52018));
    SB_LUT4 pwm_counter_1931_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n52016), .O(n56910)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_18 (.CI(n52016), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n52017));
    SB_LUT4 pwm_counter_1931_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n52015), .O(n56952)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_17 (.CI(n52015), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n52016));
    SB_LUT4 pwm_counter_1931_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n52014), .O(n56992)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_DFFR pwm_counter_1931__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n57610), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_1931_add_4_16 (.CI(n52014), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n52015));
    SB_LUT4 pwm_counter_1931_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n52013), .O(n57024)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_15 (.CI(n52013), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n52014));
    SB_LUT4 pwm_counter_1931_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n52012), .O(n57058)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_14 (.CI(n52012), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n52013));
    SB_LUT4 pwm_counter_1931_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n52011), .O(n57102)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_13 (.CI(n52011), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n52012));
    SB_LUT4 pwm_counter_1931_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n52010), .O(n57144)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_12 (.CI(n52010), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n52011));
    SB_LUT4 pwm_counter_1931_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n52009), .O(n57174)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_11 (.CI(n52009), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n52010));
    SB_LUT4 pwm_counter_1931_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n52008), .O(n57206)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_10 (.CI(n52008), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n52009));
    SB_LUT4 pwm_counter_1931_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n52007), .O(n57242)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_9 (.CI(n52007), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n52008));
    SB_LUT4 pwm_counter_1931_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n52006), .O(n57284)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_8 (.CI(n52006), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n52007));
    SB_LUT4 pwm_counter_1931_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n52005), .O(n57368)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_7 (.CI(n52005), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n52006));
    SB_LUT4 pwm_counter_1931_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n52004), .O(n57528)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_6 (.CI(n52004), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n52005));
    SB_LUT4 pwm_counter_1931_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n52003), .O(n57626)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_5 (.CI(n52003), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n52004));
    SB_LUT4 pwm_counter_1931_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n52002), .O(n57624)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_4 (.CI(n52002), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n52003));
    SB_LUT4 pwm_counter_1931_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n52001), .O(n57622)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_3 (.CI(n52001), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n52002));
    SB_LUT4 pwm_counter_1931_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n57610)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1931_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1931_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n52001));
    SB_DFFR pwm_counter_1931__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n57622), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n57624), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n57626), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n57528), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n57368), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n57284), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n57242), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n57206), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n57174), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n57144), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n57102), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n57058), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n57024), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n56992), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n56952), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n56910), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n56888), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n56860), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i19 (.Q(\pwm_counter[19] ), .C(clk32MHz), 
            .D(n56838), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n56816), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n56796), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n56776), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1931__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n56754), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n60886));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[15]), .I1(\pwm_counter[19] ), .I2(pwm_counter[16]), 
            .I3(pwm_counter[14]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n60886), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4983));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[20]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4983), .I1(n22), .I2(pwm_counter[22]), 
            .I3(pwm_counter[18]), .O(n24_adj_4984));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[17]), .I1(pwm_counter[13]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4985));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4985), .I2(n24_adj_4984), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49092_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n66108));
    defparam i49092_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49125_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n66141));
    defparam i49125_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49280_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n66296));   // verilog/pwm.v(21[8:24])
    defparam i49280_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, control_update, duty, clk16MHz, reset, 
            VCC_net, \Kp[4] , \Kp[5] , n363, \Kp[2] , \Kp[0] , \Kp[1] , 
            \Kp[6] , \Kp[3] , IntegralLimit, \PID_CONTROLLER.integral_23__N_3715 , 
            \Ki[1] , \Ki[0] , \Kp[11] , PWMLimit, \Ki[2] , \Kp[12] , 
            \Ki[3] , deadband, \Ki[4] , \Ki[11] , \Ki[5] , \Ki[6] , 
            \Ki[7] , \Ki[8] , n29183, \PID_CONTROLLER.integral , n29182, 
            n29181, n29180, n29179, n29178, n29177, n29176, n29175, 
            n29174, n29173, n29172, n29171, n29170, n29169, n29168, 
            n29164, n29160, n29159, n29158, n29157, n29156, n29155, 
            \Ki[9] , \Ki[10] , \Ki[12] , \Kp[13] , n29023, \Kp[14] , 
            \Kp[15] , \Kp[7] , \Kp[8] , \Kp[9] , \Kp[10] , n35, 
            \Ki[13] , \Ki[14] , \Ki[15] , setpoint, \motor_state[23] , 
            \motor_state[22] , \motor_state[21] , \motor_state[20] , \motor_state[19] , 
            n14, \motor_state[17] , \motor_state[16] , \encoder1_position_scaled[0] , 
            n15, n65364, n15_adj_1, \motor_state[15] , \motor_state[14] , 
            \encoder1_position_scaled[1] , n65475, \motor_state[13] , 
            \encoder1_position_scaled[2] , n65474, \motor_state[12] , 
            \motor_state[11] , \motor_state[10] , n38106, \motor_state[8] , 
            \motor_state[7] , \motor_state[6] , \motor_state[5] , \motor_state[4] , 
            \motor_state[3] , n25) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input VCC_net;
    input \Kp[4] ;
    input \Kp[5] ;
    output n363;
    input \Kp[2] ;
    input \Kp[0] ;
    input \Kp[1] ;
    input \Kp[6] ;
    input \Kp[3] ;
    input [23:0]IntegralLimit;
    output [23:0]\PID_CONTROLLER.integral_23__N_3715 ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Kp[11] ;
    input [23:0]PWMLimit;
    input \Ki[2] ;
    input \Kp[12] ;
    input \Ki[3] ;
    input [23:0]deadband;
    input \Ki[4] ;
    input \Ki[11] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input n29183;
    output [23:0]\PID_CONTROLLER.integral ;
    input n29182;
    input n29181;
    input n29180;
    input n29179;
    input n29178;
    input n29177;
    input n29176;
    input n29175;
    input n29174;
    input n29173;
    input n29172;
    input n29171;
    input n29170;
    input n29169;
    input n29168;
    input n29164;
    input n29160;
    input n29159;
    input n29158;
    input n29157;
    input n29156;
    input n29155;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[12] ;
    input \Kp[13] ;
    input n29023;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input n35;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]setpoint;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input n14;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \encoder1_position_scaled[0] ;
    input n15;
    input n65364;
    input n15_adj_1;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \encoder1_position_scaled[1] ;
    input n65475;
    input \motor_state[13] ;
    input \encoder1_position_scaled[2] ;
    input n65474;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input n38106;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    output n25;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n67853;
    wire [23:0]n356;
    
    wire n29, n67854;
    wire [16:0]n17045;
    wire [15:0]n17626;
    
    wire n165, n52274, n51760;
    wire [15:0]n17338;
    
    wire n822, n51761;
    wire [23:0]n382;
    
    wire n66412;
    wire [16:0]n16722;
    
    wire n749, n51759, n67214;
    wire [23:0]n1;
    
    wire n69092, n52275, n676, n51758, n23, n92, n67176, n603, 
        n51757, n530, n51756;
    wire [23:0]n436;
    wire [23:0]n1_adj_4980;
    
    wire n51347;
    wire [14:0]n18151;
    
    wire n52273, n457, n51755, n51346, n1117, n52272, n384, n51754, 
        n69086, n311, n51753, n51345, n1044, n52271, n971, n52270, 
        n238, n51752, n165_adj_4428, n51751, n66395, n51344, n898, 
        n52269, n23_adj_4429, n92_adj_4430, n51343, n825, n52268, 
        n51342, n51341, n752, n52267, n51340, n51339, n679, n52266, 
        n51338, n606, n52265, n51337, n51336, n533, n52264, n460, 
        n52263, n387, n52262, n314, n52261, n241, n52260, n51335, 
        n51334, n168, n52259, n51333;
    wire [14:0]n17896;
    
    wire n51732, n51332, n26, n95, n1117_adj_4431, n51731, n51331, 
        n1044_adj_4432, n51730, n51330;
    wire [13:0]n18600;
    
    wire n1120, n52258, n971_adj_4433, n51729, n51329, n1047, n52257, 
        n898_adj_4434, n51728, n51328, n825_adj_4435, n51727, n51327, 
        n974, n52256, n752_adj_4437, n51726, n679_adj_4438, n51725, 
        n51326, n901, n52255, n606_adj_4440, n51724, n533_adj_4441, 
        n51723, n51325, n828, n52254, n460_adj_4442, n51722, n387_adj_4443, 
        n51721, n755, n52253, n314_adj_4445, n51720, n241_adj_4446, 
        n51719, n67202, n47;
    wire [23:0]n1_adj_4981;
    
    wire n51324, n51323, n682, n52252, n168_adj_4450, n51718, n51322, 
        n26_adj_4452, n95_adj_4453, n51321, n609, n52251, n51320, 
        n51319, n536, n52250, n51318, n51317, n463, n52249, n51316, 
        n390_adj_4461, n52248, n317, n52247, n244, n52246, n171, 
        n52245, n51315, n29_adj_4463, n98, n51314, n51313;
    wire [6:0]n20280;
    wire [5:0]n20392;
    
    wire n560, n52244, n51312, n487, n52243;
    wire [7:0]n20216;
    wire [6:0]n20343;
    
    wire n630, n51700, n557, n51699, n51311, n484, n51698, n414, 
        n52242, n411, n51697, n51310, n338, n51696, n341, n52241, 
        n265, n51695, n51309, n192, n51694, n268, n52240, n50, 
        n119, n51308;
    wire [13:0]n18376;
    
    wire n1120_adj_4471, n51693, n195, n52239, n1047_adj_4472, n51692, 
        n51307, n974_adj_4474, n51691, n51306, n53, n122, n901_adj_4476, 
        n51690, n828_adj_4477, n51689, n51305;
    wire [12:0]n18991;
    
    wire n1050, n52238, n755_adj_4479, n51688, n51304, n977, n52237, 
        n682_adj_4481, n51687, n51303, n609_adj_4483, n51686, n904, 
        n52236, n536_adj_4484, n51685, n51302, n831, n52235, n758, 
        n52234, n685, n52233, n612, n52232, n539, n52231, n466, 
        n52230, n393_adj_4486, n52229, n320, n52228, n247, n52227, 
        n174, n52226, n32, n101;
    wire [11:0]n19328;
    
    wire n980, n52225, n907, n52224, n834, n52223, n69107, n761, 
        n52222, n688, n52221, n615, n52220, n542, n52219, n469, 
        n52218, n396_adj_4487, n52217, n323, n52216, n250, n52215, 
        n177, n52214, n35_c, n104, n60196, n490, n52213;
    wire [4:0]n20476;
    
    wire n417, n52212, n344, n52211, n271, n52210, n198, n52209, 
        n56, n125;
    wire [10:0]n19615;
    
    wire n910, n52208, n837, n52207, n764, n52206, n67196, n691, 
        n52205, n618, n52204, n545, n52203, n472, n52202, n399_adj_4488, 
        n52201, n326, n52200, n253, n52199, n180, n52198, n38, 
        n107, n69102;
    wire [9:0]n19856;
    
    wire n840, n52197, n16_adj_4489, n767, n52196, n694, n52195, 
        n621, n52194, n548, n52193, n475, n52192, n402_adj_4490, 
        n52191, n329, n52190, n256, n52189, n183, n52188, n41, 
        n110, n65413, n39319, n463_adj_4492, n51684, n390_adj_4493, 
        n51683, n317_adj_4494, n51682, n244_adj_4495, n51681, n171_adj_4496, 
        n51680;
    wire [23:0]n182;
    wire [23:0]n1_adj_4982;
    
    wire n51301, n29_adj_4499, n98_adj_4500, n51300;
    wire [12:0]n18796;
    
    wire n1050_adj_4502, n51679, n977_adj_4503, n51678, n904_adj_4504, 
        n51677, n51299, n831_adj_4506, n51676, n758_adj_4507, n51675, 
        n685_adj_4508, n51674, n612_adj_4509, n51673, n539_adj_4510, 
        n51672, n51298, n466_adj_4512, n51671, n51297, n393_adj_4514, 
        n51670, n51296, n320_adj_4516, n51669, n247_adj_4517, n51668, 
        n51295, n174_adj_4519, n51667, n66262, n51294, n32_adj_4521, 
        n101_adj_4522, n51293;
    wire [23:0]n130;
    
    wire n43, n51292, n51291, n51290, n51289, n33, n31, n66460, 
        n66447, n51288, n51287, n51286, n51285;
    wire [5:0]n20440;
    
    wire n560_adj_4535, n51650, n51284, n487_adj_4537, n51649, n51283, 
        n414_adj_4539, n51648, n51282, n341_adj_4541, n51647, n51281, 
        n268_adj_4543, n51646, n195_adj_4544, n51645, n53_adj_4545, 
        n122_adj_4546;
    wire [11:0]n19160;
    
    wire n980_adj_4547, n51644, n907_adj_4548, n51643, n8_adj_4549, 
        n834_adj_4550, n51642, n761_adj_4551, n51641, n51280, n688_adj_4553, 
        n51640, n51279, n615_adj_4555, n51639, n542_adj_4557, n51638, 
        n469_adj_4558, n51637, n396_adj_4559, n51636, n323_adj_4560, 
        n51635, n250_adj_4561, n51634, n177_adj_4562, n51633, n35_adj_4563, 
        n104_adj_4564, n24_adj_4565, n30, n10_adj_4566, n35_adj_4567, 
        n66444, n68169, n66420, n69100, n66418, n41_adj_4568, n69128, 
        n67589, n69125, n67206, n67915;
    wire [23:0]n49;
    
    wire n344_adj_4569, n417_adj_4570;
    wire [3:0]n20560;
    
    wire n6_adj_4571;
    wire [4:0]n20511;
    wire [31:0]n51;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    
    wire n52123, n52122, counter_31__N_3714, n66362, n52121, n52120;
    wire [10:0]n19472;
    
    wire n910_adj_4574, n51617, n837_adj_4575, n51616, n52119, n764_adj_4576, 
        n51615, n52118, n691_adj_4577, n51614, n69090, n52117, n618_adj_4578, 
        n51613, n67571, n69118, n52116, n545_adj_4579, n51612, n52115, 
        n472_adj_4580, n51611, n68106, n399_adj_4581, n51610, n52114, 
        n69081, n39, n326_adj_4583, n51609, n52113, n68292, n66638, 
        n253_adj_4584, n51608, n52112, n52111, n68304, n45, n69078, 
        n180_adj_4585, n51607, n52110, n38_adj_4586, n107_adj_4587, 
        n60592, n490_adj_4588, n51606, n27, n15_adj_4589, n13_adj_4590, 
        n11_adj_4591, n52109, n12_adj_4592, n52108, n52107, n51605, 
        n52106, n52105, n52104, n52103, n51604, n37, n271_adj_4594, 
        n51603, n52102, n198_adj_4595, n51602, n52101, n56_adj_4596, 
        n125_adj_4597, n52100, n52099, n52098, n52097, n37_adj_4598, 
        n68305, n52096, n52095, n52094, n52093, n204_adj_4600;
    wire [1:0]n20608;
    
    wire n131, n62, n62070, n62072, n210, n62076, n50901, n62080, 
        n8_adj_4602, n6_adj_4603, n4_adj_4604, n39_adj_4605, n68277, 
        n181;
    wire [23:0]n207;
    
    wire n155_adj_4607, n9_adj_4608, n65598, n67278, n43_adj_4609, 
        n41_adj_4610, n68219, n66436, n19_adj_4611, n17_adj_4612, 
        n67272, n25_adj_4613, n23_adj_4614, n21_adj_4615, n68124, 
        n67607, n6_adj_4616, n67855, n16_adj_4617, n8_adj_4618, n45_adj_4619, 
        n24_adj_4620, n66475, n67856, n66432, n66426, n67662, n66636, 
        n12_adj_4621, n4_adj_4622, n67847, n67848, n66329, n69113, 
        n10_adj_4623, n30_adj_4624;
    wire [9:0]n19736;
    
    wire n840_adj_4625, n51587, n767_adj_4626, n51586, n694_adj_4627, 
        n51585, n66331, n621_adj_4628, n51584, n548_adj_4630, n51583, 
        n475_adj_4631, n51582, n402_adj_4632, n51581, n68138, n329_adj_4633, 
        n51580, n256_adj_4634, n51579, n68173, n183_adj_4636, n51578, 
        n41_adj_4637, n110_adj_4638;
    wire [0:0]n10755;
    wire [0:0]n10161;
    
    wire n51247;
    wire [47:0]n257;
    wire [47:0]n306;
    
    wire n51246, n66648, n51245, n66644, n51244, n31_adj_4639, n51243, 
        n68306, n51242, n68307, n68140, n51241, n35_adj_4643, n21_adj_4644, 
        n19_adj_4645, n17_adj_4646, n9_adj_4647, n65870, n27_adj_4648, 
        n15_adj_4649, n13_adj_4650, n11_adj_4651, n65700, n33_adj_4652, 
        n12_adj_4653, n6_adj_4654, n51240, n67849, n10_adj_4656, n30_adj_4658, 
        n67850, n51239, n65914, n66830;
    wire [8:0]n19956;
    
    wire n770, n51565, n697, n51564, n51238, n624, n51563, n551, 
        n51562, n51237, n66806, n25_adj_4661, n23_adj_4662, n67973, 
        n66654, n68142, n69076, n66285, n68144, n29_adj_4663, n67310, 
        n66282, n478, n51561, n405_adj_4665, n51560, n62056, n61055, 
        n68128, n16_adj_4666, n6_adj_4667, n67835, n67836, n8_adj_4668, 
        n24_adj_4669, n332_adj_4670, n51559, n51236, n259, n51558, 
        n65609, n65600, n67660, n67655, n4_adj_4672, n67833, n51235, 
        n51234, n186_adj_4674, n51557, n67834, n65661, n65647, n68167, 
        n67657, n68324, n44, n113, n68325, n68250, n65611, n67961, 
        n40, n67963, n51029, n67664;
    wire [2:0]n20591;
    
    wire n66646, n51233, n51232, n68275, n51231, n51230, n4_adj_4678, 
        n4_adj_4679, n50826, n51229, n65916, n51228, n4_adj_4681, 
        n12_adj_4682, n51227, n11_adj_4683, n8_adj_4684, n18_adj_4685, 
        n10_adj_4686, n16_adj_4687, n15_adj_4688, n24_adj_4689, n23_adj_4690, 
        n25_adj_4691, n51226, n65950, n51225, n51224, n51223;
    wire [21:0]n10731;
    
    wire n51983, n68148, n9647, n15_adj_4693, n41_adj_4694, n39_adj_4695, 
        n45_adj_4696, n51982, n19_adj_4697, n17_adj_4698;
    wire [3:0]n20536;
    
    wire n9_adj_4699, n11_adj_4700, n13_adj_4701, n15_adj_4702, n9_adj_4703, 
        n11_adj_4704, n13_adj_4705, n9_adj_4706, n11_adj_4707, n13_adj_4708, 
        n15_adj_4709, n21_adj_4711, n19_adj_4712, n17_adj_4714, n23_adj_4716, 
        n25_adj_4717, n27_adj_4719, n51981, n51222, n51980, n51979, 
        n51978, n51977, n51976, n1096, n51975, n1023, n51974, 
        n51221, n51220, n950, n51973, n877, n51972, n804, n51971, 
        n731, n51970, n658, n51969, n51219, n585, n51968, n51218, 
        n512, n51967;
    wire [7:0]n20136;
    
    wire n700, n51515, n51217, n439_adj_4730, n51966, n33_adj_4731, 
        n627, n51514, n51216, n554, n51513, n366_adj_4733, n51965, 
        n51215, n293_adj_4734, n51964, n481, n51512, n37_adj_4735, 
        n21_adj_4736, n23_adj_4737, n238_adj_4738, n25_adj_4739, n311_adj_4740, 
        n384_adj_4741, n43_adj_4742, n457_adj_4743, n530_adj_4744, n603_adj_4745, 
        n676_adj_4746, n749_adj_4747, n822_adj_4748, n895, n968, n51214, 
        n408, n51511, n220, n51963, n335_adj_4749, n51510, n262, 
        n51509, n1041, n1114, n89, n147_adj_4750, n51962, n189_adj_4751, 
        n51508, n47_adj_4752, n116, n20_adj_4753, n51213, n162_adj_4755, 
        n235, n27_adj_4756, n5_adj_4757, n74, n308, n51212, n381, 
        n454_adj_4758, n51211, n527, n600, n29_adj_4759, n673, n746, 
        n819, n892;
    wire [20:0]n12441;
    
    wire n51961, n965, n1038, n51960, n31_adj_4760, n66230, n1111, 
        n86, n66213, n17_adj_4761, n159_adj_4762, n51210, n232, 
        n12_adj_4764, n305_adj_4765, n378_adj_4766, n51959, n51958, 
        n451_adj_4767, n524, n597, n51957, n51209, n670, n743, 
        n10_adj_4768, n816, n51208, n889, n962, n51956, n1035, 
        n1108, n83, n14_adj_4770, n51207, n156_adj_4771, n229_adj_4772, 
        n302_adj_4773, n30_adj_4775, n375_adj_4776, n448_adj_4777, n51955, 
        n66259, n67114, n521, n594, n667, n740, n1099, n51954, 
        n813, n886, n67100, n959, n1032, n1026, n51953, n1105, 
        n80, n11_adj_4778, n153_adj_4779, n953, n51952, n68088, 
        n226_adj_4780, n880, n51951, n299_adj_4781, n372_adj_4782, 
        n67519, n445_adj_4783, n518, n591, n664, n737, n810, n68211, 
        n883, n956, n807, n51950, n1029, n734, n51949, n51206, 
        n661, n51948, n588, n51947, n515, n51946, n1102, n77, 
        n442_adj_4784, n51945, n369_adj_4785, n51944, n296_adj_4786, 
        n51943, n8_adj_4787, n150_adj_4788, n223, n51942, n223_adj_4789, 
        n296_adj_4790, n150_adj_4791, n51941, n369_adj_4792, n442_adj_4793, 
        n8_adj_4794, n77_adj_4795, n515_adj_4796;
    wire [19:0]n13743;
    
    wire n51940, n588_adj_4797, n661_adj_4798, n51939, n734_adj_4799, 
        n807_adj_4800, n880_adj_4801, n953_adj_4802, n51938, n1026_adj_4803, 
        n1099_adj_4804, n74_adj_4805, n5_adj_4806, n147_adj_4807, n51937, 
        n51936, n220_adj_4808, n51935, n1102_adj_4809, n51934, n293_adj_4810, 
        n1029_adj_4811, n51933, n366_adj_4812, n956_adj_4813, n51932, 
        n883_adj_4814, n51931, n439_adj_4815, n810_adj_4816, n51930, 
        n737_adj_4817, n51929, n512_adj_4818, n585_adj_4819, n51205, 
        n16_adj_4820, n658_adj_4821, n731_adj_4822, n664_adj_4823, n51928, 
        n591_adj_4824, n51927, n518_adj_4825, n51926, n804_adj_4826, 
        n877_adj_4827, n950_adj_4828, n1023_adj_4829, n1096_adj_4830, 
        n119_adj_4831, n50_adj_4832, n192_adj_4833, n265_adj_4834, n338_adj_4835, 
        n411_adj_4836, n484_adj_4837, n557_adj_4838, n630_adj_4839, 
        n445_adj_4840, n51925, n895_adj_4841, n968_adj_4842, n1041_adj_4843, 
        n6_adj_4844, n67841, n1114_adj_4845, n372_adj_4846, n51924, 
        n299_adj_4847, n51923, n51204, n226_adj_4848, n51922, n153_adj_4849, 
        n51921, n11_adj_4850, n80_adj_4851, n116_adj_4852, n47_adj_4853, 
        n189_adj_4854;
    wire [18:0]n14896;
    
    wire n51920, n51919, n262_adj_4855, n335_adj_4856, n408_adj_4857, 
        n67842, n481_adj_4858, n554_adj_4859, n627_adj_4860, n51203, 
        n700_adj_4861, n51202, n51918, n89_adj_4862, n20_adj_4863, 
        n162_adj_4864, n51917, n51916, n1105_adj_4865, n51915, n1032_adj_4866, 
        n51914, n235_adj_4867, n308_adj_4868, n959_adj_4869, n51913, 
        n886_adj_4870, n51912, n813_adj_4871, n51911, n381_adj_4872, 
        n454_adj_4873, n527_adj_4874, n51201, n8_adj_4875, n600_adj_4876, 
        n51200, n673_adj_4877, n740_adj_4878, n51910, n746_adj_4879, 
        n667_adj_4880, n51909, n819_adj_4881, n892_adj_4882, n965_adj_4883, 
        n1038_adj_4884, n1111_adj_4885, n594_adj_4886, n51908, n521_adj_4887, 
        n51907, n448_adj_4888, n51906, n375_adj_4889, n51905, n302_adj_4890, 
        n51904, n229_adj_4891, n51903, n156_adj_4892, n51902, n14_adj_4893, 
        n83_adj_4894;
    wire [8:0]n20055;
    
    wire n770_adj_4895, n51901, n697_adj_4896, n51900, n624_adj_4897, 
        n51899, n51199, n51198, n551_adj_4898, n51898, n478_adj_4899, 
        n51897, n405_adj_4900, n51896, n332_adj_4901, n51895, n259_adj_4902, 
        n51894, n186_adj_4903, n51893, n44_adj_4904, n113_adj_4905, 
        n51197, n51196, n51195, n51194;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n86_adj_4909, n17_adj_4910, n159_adj_4911, n51193, n51192, 
        n232_adj_4912, n305_adj_4913, n51191, n378_adj_4914, n51190, 
        n51189, n451_adj_4915, n524_adj_4916, n597_adj_4917, n24_adj_4918, 
        n670_adj_4919, n743_adj_4920, n66183, n66177, n67666, n816_adj_4921, 
        n889_adj_4922, n962_adj_4923, n66656, n51188, n51187, n1035_adj_4924, 
        n1108_adj_4925, n51186, n4_adj_4926, n51185, n67839, n67840;
    wire [17:0]n15911;
    
    wire n51869, n51868, n51867, n51184, n51866, n51865, n51183, 
        n51864, n51182, n66207, n51863, n51862, n51861, n51181, 
        n51860, n51859, n51858, n51857, n51856, n51855, n51180, 
        n51854, n51853, n51179, n51852, n66205, n68175, n66658, 
        n68310, n51810, n51809, n51808, n51807, n51806, n51805, 
        n51804, n51803, n51802, n51801, n51800, n51799, n51798, 
        n51797, n51796, n51795, n51794, n51793, n51792, n51791, 
        n51790, n51789, n51788, n51787, n51786, n68311, n51766, 
        n51765, n51764, n51763, n51762, n68269, n66187, n68146, 
        n66664, n66082, n409, n41_adj_4927, n66119, n52413, n52412, 
        n52411, n52410, n52409, n52408, n52407;
    wire [21:0]n11262;
    
    wire n52406, n52405, n52404, n39_adj_4928, n52403, n52402, n52401, 
        n52400, n52399, n52398, n52397, n52396, n52395, n52394, 
        n52393, n52392, n52391, n52390, n52389, n52388, n52387, 
        n52386, n52385;
    wire [20:0]n12924;
    
    wire n52384, n52383, n52382, n52381, n52380, n52379, n52378, 
        n52377, n52376, n52375, n52374, n52373, n52372, n52371, 
        n52370, n52369, n52368, n45_adj_4929, n52367, n52366, n52365, 
        n52364;
    wire [19:0]n14183;
    
    wire n52363, n52362, n52361, n52360, n52359, n52358, n52357, 
        n52356, n52355, n52354, n52353, n52352, n52351, n52350, 
        n52349, n52348, n52347, n52346, n52345, n52344;
    wire [18:0]n15295;
    
    wire n52343, n52342, n52341, n52340, n52339, n52338, n52337, 
        n17_adj_4930, n52336, n52335, n52334, n52333, n52332, n52331, 
        n52330, n19_adj_4931, n52329, n52328, n52327, n52326, n52325;
    wire [17:0]n16271;
    
    wire n52324, n52323, n52322, n52321, n52320, n52319, n52318, 
        n52317, n52316, n52315, n52314, n52313, n52312, n52311, 
        n52310, n52309, n52308, n52307, n52306, n52305, n52304, 
        n43_adj_4932, n52303, n52302, n52301, n52300, n52299, n52298, 
        n52297, n52296, n52295, n52294, n52293, n52292, n52291, 
        n52290, n52289, n52288, n52287, n52286, n52285, n52284, 
        n52283, n52282, n52281, n52280, n52279, n52278, n52277, 
        n52276, n33_adj_4933, n35_adj_4934, n37_adj_4935, n27_adj_4936, 
        n29_adj_4937, n31_adj_4938, n21_adj_4939, n23_adj_4940, n25_adj_4941, 
        n66143, n66131, n12_adj_4942, n10_adj_4943, n30_adj_4944, 
        n9649, n27546, n66173, n67038, n27541, n27536, n27531, 
        n27526, n67028, n68072, n67481, n27521, n68205, n6_adj_4945, 
        n67829, n16_adj_4946, n27516, n27511, n8_adj_4947, n27506, 
        n27501, n24_adj_4948, n67830, n27496, n66088, n27219, n67668, 
        n27491, n27486, n66666, n27481, n4_adj_4949, n27476, n27471, 
        n27466, n67827, n27461, n67828, n66123, n27456, n27451, 
        n68177, n66668, n68312, n27446, n68313, n27441, n68267, 
        n66092, n27436, n68150, n66674, n68152, n68153;
    wire [1:0]n20600;
    
    wire n50810, n4_adj_4951, n6_adj_4952, n50958, n4_adj_4953;
    wire [2:0]n20576;
    
    wire n6_adj_4954, n62_adj_4955, n131_adj_4956, n204_adj_4957, n50876, 
        n62030, n62034, n62032, n62040, n4_adj_4960, n8_adj_4961, 
        n41_adj_4962, n43_adj_4963, n39_adj_4964, n37_adj_4965, n45_adj_4966, 
        n29_adj_4967, n31_adj_4968, n33_adj_4969, n35_adj_4970, n65987, 
        n65964, n12_adj_4972, n10_adj_4973, n30_adj_4974, n66033, 
        n6_adj_4975, n66926, n66918, n68050, n67415, n68199, n16_adj_4976, 
        n67441, n67442, n8_adj_4977, n24_adj_4978, n65918, n67652, 
        n66626, n4_adj_4979, n67439, n67440, n65954, n68028, n66628, 
        n68270, n68271, n68204, n65927, n67957, n66634, n68136;
    
    SB_LUT4 i50838_3_lut (.I0(n67853), .I1(n356[14]), .I2(n29), .I3(GND_net), 
            .O(n67854));   // verilog/motorControl.v(51[12:29])
    defparam i50838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4941_3_lut (.I0(GND_net), .I1(n17626[0]), .I2(n165), .I3(n52274), 
            .O(n17045[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_12 (.CI(n51760), .I0(n17338[9]), .I1(n822), .CO(n51761));
    SB_LUT4 i49396_4_lut (.I0(n356[6]), .I1(n356[5]), .I2(n382[6]), .I3(n382[5]), 
            .O(n66412));
    defparam i49396_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 add_4924_11_lut (.I0(GND_net), .I1(n17338[8]), .I2(n749), 
            .I3(n51759), .O(n16722[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50198_3_lut (.I0(n356[7]), .I1(n66412), .I2(n382[7]), .I3(GND_net), 
            .O(n67214));
    defparam i50198_3_lut.LUT_INIT = 16'hdede;
    SB_DFFER result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n1[0]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 LessThan_21_i27_rep_75_2_lut (.I0(n356[13]), .I1(n382[13]), 
            .I2(GND_net), .I3(GND_net), .O(n69092));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i27_rep_75_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4941_3 (.CI(n52274), .I0(n17626[0]), .I1(n165), .CO(n52275));
    SB_CARRY add_4924_11 (.CI(n51759), .I0(n17338[8]), .I1(n749), .CO(n51760));
    SB_LUT4 add_4924_10_lut (.I0(GND_net), .I1(n17338[7]), .I2(n676), 
            .I3(n51758), .O(n16722[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4941_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n17045[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_10 (.CI(n51758), .I0(n17338[7]), .I1(n676), .CO(n51759));
    SB_LUT4 i50160_4_lut (.I0(n356[14]), .I1(n69092), .I2(n382[14]), .I3(n67214), 
            .O(n67176));
    defparam i50160_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_4924_9_lut (.I0(GND_net), .I1(n17338[6]), .I2(n603), .I3(n51757), 
            .O(n16722[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n52274));
    SB_CARRY add_4924_9 (.CI(n51757), .I0(n17338[6]), .I1(n603), .CO(n51758));
    SB_LUT4 add_4924_8_lut (.I0(GND_net), .I1(n17338[5]), .I2(n530), .I3(n51756), 
            .O(n16722[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[23]), 
            .I3(n51347), .O(n436[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4975_17_lut (.I0(GND_net), .I1(n18151[14]), .I2(GND_net), 
            .I3(n52273), .O(n17626[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_8 (.CI(n51756), .I0(n17338[5]), .I1(n530), .CO(n51757));
    SB_LUT4 add_4924_7_lut (.I0(GND_net), .I1(n17338[4]), .I2(n457), .I3(n51755), 
            .O(n16722[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[22]), 
            .I3(n51346), .O(n436[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4975_16_lut (.I0(GND_net), .I1(n18151[13]), .I2(n1117), 
            .I3(n52272), .O(n17626[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_7 (.CI(n51755), .I0(n17338[4]), .I1(n457), .CO(n51756));
    SB_LUT4 add_4924_6_lut (.I0(GND_net), .I1(n17338[3]), .I2(n384), .I3(n51754), 
            .O(n16722[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_24 (.CI(n51346), .I0(GND_net), .I1(n1_adj_4980[22]), 
            .CO(n51347));
    SB_CARRY add_4975_16 (.CI(n52272), .I0(n18151[13]), .I1(n1117), .CO(n52273));
    SB_LUT4 LessThan_21_i31_rep_69_2_lut (.I0(n356[15]), .I1(n382[15]), 
            .I2(GND_net), .I3(GND_net), .O(n69086));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i31_rep_69_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4924_6 (.CI(n51754), .I0(n17338[3]), .I1(n384), .CO(n51755));
    SB_LUT4 add_4924_5_lut (.I0(GND_net), .I1(n17338[2]), .I2(n311), .I3(n51753), 
            .O(n16722[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[21]), 
            .I3(n51345), .O(n436[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4975_15_lut (.I0(GND_net), .I1(n18151[12]), .I2(n1044), 
            .I3(n52271), .O(n17626[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_15 (.CI(n52271), .I0(n18151[12]), .I1(n1044), .CO(n52272));
    SB_LUT4 add_4975_14_lut (.I0(GND_net), .I1(n18151[11]), .I2(n971), 
            .I3(n52270), .O(n17626[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_5 (.CI(n51753), .I0(n17338[2]), .I1(n311), .CO(n51754));
    SB_LUT4 add_4924_4_lut (.I0(GND_net), .I1(n17338[1]), .I2(n238), .I3(n51752), 
            .O(n16722[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_23 (.CI(n51345), .I0(GND_net), .I1(n1_adj_4980[21]), 
            .CO(n51346));
    SB_CARRY add_4924_4 (.CI(n51752), .I0(n17338[1]), .I1(n238), .CO(n51753));
    SB_LUT4 add_4924_3_lut (.I0(GND_net), .I1(n17338[0]), .I2(n165_adj_4428), 
            .I3(n51751), .O(n16722[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49379_4_lut (.I0(n356[8]), .I1(n356[4]), .I2(n382[8]), .I3(n382[4]), 
            .O(n66395));
    defparam i49379_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[20]), 
            .I3(n51344), .O(n436[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_14 (.CI(n52270), .I0(n18151[11]), .I1(n971), .CO(n52271));
    SB_CARRY add_4924_3 (.CI(n51751), .I0(n17338[0]), .I1(n165_adj_4428), 
            .CO(n51752));
    SB_CARRY unary_minus_26_add_3_22 (.CI(n51344), .I0(GND_net), .I1(n1_adj_4980[20]), 
            .CO(n51345));
    SB_LUT4 add_4975_13_lut (.I0(GND_net), .I1(n18151[10]), .I2(n898), 
            .I3(n52269), .O(n17626[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_13 (.CI(n52269), .I0(n18151[10]), .I1(n898), .CO(n52270));
    SB_LUT4 add_4924_2_lut (.I0(GND_net), .I1(n23_adj_4429), .I2(n92_adj_4430), 
            .I3(GND_net), .O(n16722[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_2 (.CI(GND_net), .I0(n23_adj_4429), .I1(n92_adj_4430), 
            .CO(n51751));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[19]), 
            .I3(n51343), .O(n436[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_21 (.CI(n51343), .I0(GND_net), .I1(n1_adj_4980[19]), 
            .CO(n51344));
    SB_LUT4 add_4975_12_lut (.I0(GND_net), .I1(n18151[9]), .I2(n825), 
            .I3(n52268), .O(n17626[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[18]), 
            .I3(n51342), .O(n436[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_20 (.CI(n51342), .I0(GND_net), .I1(n1_adj_4980[18]), 
            .CO(n51343));
    SB_CARRY add_4975_12 (.CI(n52268), .I0(n18151[9]), .I1(n825), .CO(n52269));
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[17]), 
            .I3(n51341), .O(n436[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_19 (.CI(n51341), .I0(GND_net), .I1(n1_adj_4980[17]), 
            .CO(n51342));
    SB_LUT4 add_4975_11_lut (.I0(GND_net), .I1(n18151[8]), .I2(n752), 
            .I3(n52267), .O(n17626[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[16]), 
            .I3(n51340), .O(n436[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_18 (.CI(n51340), .I0(GND_net), .I1(n1_adj_4980[16]), 
            .CO(n51341));
    SB_CARRY add_4975_11 (.CI(n52267), .I0(n18151[8]), .I1(n752), .CO(n52268));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[15]), 
            .I3(n51339), .O(n436[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_17 (.CI(n51339), .I0(GND_net), .I1(n1_adj_4980[15]), 
            .CO(n51340));
    SB_LUT4 add_4975_10_lut (.I0(GND_net), .I1(n18151[7]), .I2(n679), 
            .I3(n52266), .O(n17626[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_10 (.CI(n52266), .I0(n18151[7]), .I1(n679), .CO(n52267));
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[14]), 
            .I3(n51338), .O(n436[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_16 (.CI(n51338), .I0(GND_net), .I1(n1_adj_4980[14]), 
            .CO(n51339));
    SB_LUT4 add_4975_9_lut (.I0(GND_net), .I1(n18151[6]), .I2(n606), .I3(n52265), 
            .O(n17626[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[13]), 
            .I3(n51337), .O(n436[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_15 (.CI(n51337), .I0(GND_net), .I1(n1_adj_4980[13]), 
            .CO(n51338));
    SB_CARRY add_4975_9 (.CI(n52265), .I0(n18151[6]), .I1(n606), .CO(n52266));
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[12]), 
            .I3(n51336), .O(n436[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_14 (.CI(n51336), .I0(GND_net), .I1(n1_adj_4980[12]), 
            .CO(n51337));
    SB_LUT4 add_4975_8_lut (.I0(GND_net), .I1(n18151[5]), .I2(n533), .I3(n52264), 
            .O(n17626[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_8 (.CI(n52264), .I0(n18151[5]), .I1(n533), .CO(n52265));
    SB_LUT4 add_4975_7_lut (.I0(GND_net), .I1(n18151[4]), .I2(n460), .I3(n52263), 
            .O(n17626[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_7 (.CI(n52263), .I0(n18151[4]), .I1(n460), .CO(n52264));
    SB_LUT4 add_4975_6_lut (.I0(GND_net), .I1(n18151[3]), .I2(n387), .I3(n52262), 
            .O(n17626[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_6 (.CI(n52262), .I0(n18151[3]), .I1(n387), .CO(n52263));
    SB_LUT4 add_4975_5_lut (.I0(GND_net), .I1(n18151[2]), .I2(n314), .I3(n52261), 
            .O(n17626[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4975_5 (.CI(n52261), .I0(n18151[2]), .I1(n314), .CO(n52262));
    SB_LUT4 add_4975_4_lut (.I0(GND_net), .I1(n18151[1]), .I2(n241), .I3(n52260), 
            .O(n17626[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[11]), 
            .I3(n51335), .O(n436[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n51335), .I0(GND_net), .I1(n1_adj_4980[11]), 
            .CO(n51336));
    SB_CARRY add_4975_4 (.CI(n52260), .I0(n18151[1]), .I1(n241), .CO(n52261));
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[10]), 
            .I3(n51334), .O(n436[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_12 (.CI(n51334), .I0(GND_net), .I1(n1_adj_4980[10]), 
            .CO(n51335));
    SB_LUT4 add_4975_3_lut (.I0(GND_net), .I1(n18151[0]), .I2(n168), .I3(n52259), 
            .O(n17626[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[9]), 
            .I3(n51333), .O(n436[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_11 (.CI(n51333), .I0(GND_net), .I1(n1_adj_4980[9]), 
            .CO(n51334));
    SB_CARRY add_4975_3 (.CI(n52259), .I0(n18151[0]), .I1(n168), .CO(n52260));
    SB_LUT4 add_4959_17_lut (.I0(GND_net), .I1(n17896[14]), .I2(GND_net), 
            .I3(n51732), .O(n17338[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[8]), 
            .I3(n51332), .O(n436[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n51332), .I0(GND_net), .I1(n1_adj_4980[8]), 
            .CO(n51333));
    SB_LUT4 add_4975_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n17626[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4975_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_16_lut (.I0(GND_net), .I1(n17896[13]), .I2(n1117_adj_4431), 
            .I3(n51731), .O(n17338[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_16 (.CI(n51731), .I0(n17896[13]), .I1(n1117_adj_4431), 
            .CO(n51732));
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[7]), 
            .I3(n51331), .O(n436[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_9 (.CI(n51331), .I0(GND_net), .I1(n1_adj_4980[7]), 
            .CO(n51332));
    SB_CARRY add_4975_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n52259));
    SB_LUT4 add_4959_15_lut (.I0(GND_net), .I1(n17896[12]), .I2(n1044_adj_4432), 
            .I3(n51730), .O(n17338[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_15 (.CI(n51730), .I0(n17896[12]), .I1(n1044_adj_4432), 
            .CO(n51731));
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[6]), 
            .I3(n51330), .O(n436[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_8 (.CI(n51330), .I0(GND_net), .I1(n1_adj_4980[6]), 
            .CO(n51331));
    SB_LUT4 add_5005_16_lut (.I0(GND_net), .I1(n18600[13]), .I2(n1120), 
            .I3(n52258), .O(n18151[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_14_lut (.I0(GND_net), .I1(n17896[11]), .I2(n971_adj_4433), 
            .I3(n51729), .O(n17338[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_14 (.CI(n51729), .I0(n17896[11]), .I1(n971_adj_4433), 
            .CO(n51730));
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[5]), 
            .I3(n51329), .O(n436[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n51329), .I0(GND_net), .I1(n1_adj_4980[5]), 
            .CO(n51330));
    SB_LUT4 add_5005_15_lut (.I0(GND_net), .I1(n18600[12]), .I2(n1047), 
            .I3(n52257), .O(n18151[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_13_lut (.I0(GND_net), .I1(n17896[10]), .I2(n898_adj_4434), 
            .I3(n51728), .O(n17338[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_13 (.CI(n51728), .I0(n17896[10]), .I1(n898_adj_4434), 
            .CO(n51729));
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[4]), 
            .I3(n51328), .O(n436[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_6 (.CI(n51328), .I0(GND_net), .I1(n1_adj_4980[4]), 
            .CO(n51329));
    SB_CARRY add_5005_15 (.CI(n52257), .I0(n18600[12]), .I1(n1047), .CO(n52258));
    SB_LUT4 add_4959_12_lut (.I0(GND_net), .I1(n17896[9]), .I2(n825_adj_4435), 
            .I3(n51727), .O(n17338[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_12 (.CI(n51727), .I0(n17896[9]), .I1(n825_adj_4435), 
            .CO(n51728));
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[3]), 
            .I3(n51327), .O(n436[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_14_lut (.I0(GND_net), .I1(n18600[11]), .I2(n974), 
            .I3(n52256), .O(n18151[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_11_lut (.I0(GND_net), .I1(n17896[8]), .I2(n752_adj_4437), 
            .I3(n51726), .O(n17338[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_11 (.CI(n51726), .I0(n17896[8]), .I1(n752_adj_4437), 
            .CO(n51727));
    SB_CARRY unary_minus_26_add_3_5 (.CI(n51327), .I0(GND_net), .I1(n1_adj_4980[3]), 
            .CO(n51328));
    SB_CARRY add_5005_14 (.CI(n52256), .I0(n18600[11]), .I1(n974), .CO(n52257));
    SB_LUT4 add_4959_10_lut (.I0(GND_net), .I1(n17896[7]), .I2(n679_adj_4438), 
            .I3(n51725), .O(n17338[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_10 (.CI(n51725), .I0(n17896[7]), .I1(n679_adj_4438), 
            .CO(n51726));
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[2]), 
            .I3(n51326), .O(n436[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_13_lut (.I0(GND_net), .I1(n18600[10]), .I2(n901), 
            .I3(n52255), .O(n18151[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_9_lut (.I0(GND_net), .I1(n17896[6]), .I2(n606_adj_4440), 
            .I3(n51724), .O(n17338[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_9 (.CI(n51724), .I0(n17896[6]), .I1(n606_adj_4440), 
            .CO(n51725));
    SB_CARRY unary_minus_26_add_3_4 (.CI(n51326), .I0(GND_net), .I1(n1_adj_4980[2]), 
            .CO(n51327));
    SB_CARRY add_5005_13 (.CI(n52255), .I0(n18600[10]), .I1(n901), .CO(n52256));
    SB_LUT4 add_4959_8_lut (.I0(GND_net), .I1(n17896[5]), .I2(n533_adj_4441), 
            .I3(n51723), .O(n17338[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_8 (.CI(n51723), .I0(n17896[5]), .I1(n533_adj_4441), 
            .CO(n51724));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[1]), 
            .I3(n51325), .O(n436[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_12_lut (.I0(GND_net), .I1(n18600[9]), .I2(n828), 
            .I3(n52254), .O(n18151[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_7_lut (.I0(GND_net), .I1(n17896[4]), .I2(n460_adj_4442), 
            .I3(n51722), .O(n17338[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_7 (.CI(n51722), .I0(n17896[4]), .I1(n460_adj_4442), 
            .CO(n51723));
    SB_CARRY unary_minus_26_add_3_3 (.CI(n51325), .I0(GND_net), .I1(n1_adj_4980[1]), 
            .CO(n51326));
    SB_CARRY add_5005_12 (.CI(n52254), .I0(n18600[9]), .I1(n828), .CO(n52255));
    SB_LUT4 add_4959_6_lut (.I0(GND_net), .I1(n17896[3]), .I2(n387_adj_4443), 
            .I3(n51721), .O(n17338[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_6 (.CI(n51721), .I0(n17896[3]), .I1(n387_adj_4443), 
            .CO(n51722));
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4980[0]), 
            .I3(VCC_net), .O(n436[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_11_lut (.I0(GND_net), .I1(n18600[8]), .I2(n755), 
            .I3(n52253), .O(n18151[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_5_lut (.I0(GND_net), .I1(n17896[2]), .I2(n314_adj_4445), 
            .I3(n51720), .O(n17338[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_5 (.CI(n51720), .I0(n17896[2]), .I1(n314_adj_4445), 
            .CO(n51721));
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4980[0]), 
            .CO(n51325));
    SB_CARRY add_5005_11 (.CI(n52253), .I0(n18600[8]), .I1(n755), .CO(n52254));
    SB_LUT4 add_4959_4_lut (.I0(GND_net), .I1(n17896[1]), .I2(n241_adj_4446), 
            .I3(n51719), .O(n17338[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_4 (.CI(n51719), .I0(n17896[1]), .I1(n241_adj_4446), 
            .CO(n51720));
    SB_LUT4 i50186_3_lut (.I0(n356[9]), .I1(n66395), .I2(n382[9]), .I3(GND_net), 
            .O(n67202));
    defparam i50186_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n356[23]), .I1(GND_net), .I2(n1_adj_4981[23]), 
            .I3(n51324), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[22]), 
            .I3(n51323), .O(n382[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_10_lut (.I0(GND_net), .I1(n18600[7]), .I2(n682), 
            .I3(n52252), .O(n18151[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4959_3_lut (.I0(GND_net), .I1(n17896[0]), .I2(n168_adj_4450), 
            .I3(n51718), .O(n17338[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_3 (.CI(n51718), .I0(n17896[0]), .I1(n168_adj_4450), 
            .CO(n51719));
    SB_CARRY unary_minus_20_add_3_24 (.CI(n51323), .I0(GND_net), .I1(n1_adj_4981[22]), 
            .CO(n51324));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[21]), 
            .I3(n51322), .O(n382[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_10 (.CI(n52252), .I0(n18600[7]), .I1(n682), .CO(n52253));
    SB_LUT4 add_4959_2_lut (.I0(GND_net), .I1(n26_adj_4452), .I2(n95_adj_4453), 
            .I3(GND_net), .O(n17338[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4959_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4959_2 (.CI(GND_net), .I0(n26_adj_4452), .I1(n95_adj_4453), 
            .CO(n51718));
    SB_CARRY unary_minus_20_add_3_23 (.CI(n51322), .I0(GND_net), .I1(n1_adj_4981[21]), 
            .CO(n51323));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[20]), 
            .I3(n51321), .O(n382[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_9_lut (.I0(GND_net), .I1(n18600[6]), .I2(n609), .I3(n52251), 
            .O(n18151[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n51321), .I0(GND_net), .I1(n1_adj_4981[20]), 
            .CO(n51322));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[19]), 
            .I3(n51320), .O(n382[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_9 (.CI(n52251), .I0(n18600[6]), .I1(n609), .CO(n52252));
    SB_CARRY unary_minus_20_add_3_21 (.CI(n51320), .I0(GND_net), .I1(n1_adj_4981[19]), 
            .CO(n51321));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[18]), 
            .I3(n51319), .O(n382[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_8_lut (.I0(GND_net), .I1(n18600[5]), .I2(n536), .I3(n52250), 
            .O(n18151[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n51319), .I0(GND_net), .I1(n1_adj_4981[18]), 
            .CO(n51320));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[17]), 
            .I3(n51318), .O(n382[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_8 (.CI(n52250), .I0(n18600[5]), .I1(n536), .CO(n52251));
    SB_CARRY unary_minus_20_add_3_19 (.CI(n51318), .I0(GND_net), .I1(n1_adj_4981[17]), 
            .CO(n51319));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[16]), 
            .I3(n51317), .O(n382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5005_7_lut (.I0(GND_net), .I1(n18600[4]), .I2(n463), .I3(n52249), 
            .O(n18151[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n51317), .I0(GND_net), .I1(n1_adj_4981[16]), 
            .CO(n51318));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[15]), 
            .I3(n51316), .O(n382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_7 (.CI(n52249), .I0(n18600[4]), .I1(n463), .CO(n52250));
    SB_LUT4 add_5005_6_lut (.I0(GND_net), .I1(n18600[3]), .I2(n390_adj_4461), 
            .I3(n52248), .O(n18151[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_6 (.CI(n52248), .I0(n18600[3]), .I1(n390_adj_4461), 
            .CO(n52249));
    SB_LUT4 add_5005_5_lut (.I0(GND_net), .I1(n18600[2]), .I2(n317), .I3(n52247), 
            .O(n18151[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_5 (.CI(n52247), .I0(n18600[2]), .I1(n317), .CO(n52248));
    SB_LUT4 add_5005_4_lut (.I0(GND_net), .I1(n18600[1]), .I2(n244), .I3(n52246), 
            .O(n18151[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_4 (.CI(n52246), .I0(n18600[1]), .I1(n244), .CO(n52247));
    SB_LUT4 add_5005_3_lut (.I0(GND_net), .I1(n18600[0]), .I2(n171), .I3(n52245), 
            .O(n18151[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n51316), .I0(GND_net), .I1(n1_adj_4981[15]), 
            .CO(n51317));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[14]), 
            .I3(n51315), .O(n382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5005_3 (.CI(n52245), .I0(n18600[0]), .I1(n171), .CO(n52246));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n51315), .I0(GND_net), .I1(n1_adj_4981[14]), 
            .CO(n51316));
    SB_LUT4 add_5005_2_lut (.I0(GND_net), .I1(n29_adj_4463), .I2(n98), 
            .I3(GND_net), .O(n18151[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5005_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[13]), 
            .I3(n51314), .O(n382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n51314), .I0(GND_net), .I1(n1_adj_4981[13]), 
            .CO(n51315));
    SB_CARRY add_5005_2 (.CI(GND_net), .I0(n29_adj_4463), .I1(n98), .CO(n52245));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[12]), 
            .I3(n51313), .O(n382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5166_8_lut (.I0(GND_net), .I1(n20392[5]), .I2(n560), .I3(n52244), 
            .O(n20280[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n51313), .I0(GND_net), .I1(n1_adj_4981[12]), 
            .CO(n51314));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[11]), 
            .I3(n51312), .O(n382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5166_7_lut (.I0(GND_net), .I1(n20392[4]), .I2(n487), .I3(n52243), 
            .O(n20280[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_9_lut (.I0(GND_net), .I1(n20343[6]), .I2(n630), .I3(n51700), 
            .O(n20216[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n51312), .I0(GND_net), .I1(n1_adj_4981[11]), 
            .CO(n51313));
    SB_CARRY add_5166_7 (.CI(n52243), .I0(n20392[4]), .I1(n487), .CO(n52244));
    SB_LUT4 add_5159_8_lut (.I0(GND_net), .I1(n20343[5]), .I2(n557), .I3(n51699), 
            .O(n20216[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_8 (.CI(n51699), .I0(n20343[5]), .I1(n557), .CO(n51700));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[10]), 
            .I3(n51311), .O(n382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n51311), .I0(GND_net), .I1(n1_adj_4981[10]), 
            .CO(n51312));
    SB_LUT4 add_5159_7_lut (.I0(GND_net), .I1(n20343[4]), .I2(n484), .I3(n51698), 
            .O(n20216[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5166_6_lut (.I0(GND_net), .I1(n20392[3]), .I2(n414), .I3(n52242), 
            .O(n20280[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_7 (.CI(n51698), .I0(n20343[4]), .I1(n484), .CO(n51699));
    SB_LUT4 add_5159_6_lut (.I0(GND_net), .I1(n20343[3]), .I2(n411), .I3(n51697), 
            .O(n20216[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[9]), 
            .I3(n51310), .O(n382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_6 (.CI(n52242), .I0(n20392[3]), .I1(n414), .CO(n52243));
    SB_CARRY add_5159_6 (.CI(n51697), .I0(n20343[3]), .I1(n411), .CO(n51698));
    SB_LUT4 add_5159_5_lut (.I0(GND_net), .I1(n20343[2]), .I2(n338), .I3(n51696), 
            .O(n20216[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n51310), .I0(GND_net), .I1(n1_adj_4981[9]), 
            .CO(n51311));
    SB_LUT4 add_5166_5_lut (.I0(GND_net), .I1(n20392[2]), .I2(n341), .I3(n52241), 
            .O(n20280[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_5 (.CI(n51696), .I0(n20343[2]), .I1(n338), .CO(n51697));
    SB_LUT4 add_5159_4_lut (.I0(GND_net), .I1(n20343[1]), .I2(n265), .I3(n51695), 
            .O(n20216[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[8]), 
            .I3(n51309), .O(n382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_5 (.CI(n52241), .I0(n20392[2]), .I1(n341), .CO(n52242));
    SB_CARRY add_5159_4 (.CI(n51695), .I0(n20343[1]), .I1(n265), .CO(n51696));
    SB_LUT4 add_5159_3_lut (.I0(GND_net), .I1(n20343[0]), .I2(n192), .I3(n51694), 
            .O(n20216[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n51309), .I0(GND_net), .I1(n1_adj_4981[8]), 
            .CO(n51310));
    SB_LUT4 add_5166_4_lut (.I0(GND_net), .I1(n20392[1]), .I2(n268), .I3(n52240), 
            .O(n20280[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_3 (.CI(n51694), .I0(n20343[0]), .I1(n192), .CO(n51695));
    SB_LUT4 add_5159_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n20216[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[7]), 
            .I3(n51308), .O(n382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_4 (.CI(n52240), .I0(n20392[1]), .I1(n268), .CO(n52241));
    SB_CARRY add_5159_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n51694));
    SB_LUT4 add_4990_16_lut (.I0(GND_net), .I1(n18376[13]), .I2(n1120_adj_4471), 
            .I3(n51693), .O(n17896[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n51308), .I0(GND_net), .I1(n1_adj_4981[7]), 
            .CO(n51309));
    SB_LUT4 add_5166_3_lut (.I0(GND_net), .I1(n20392[0]), .I2(n195), .I3(n52239), 
            .O(n20280[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4990_15_lut (.I0(GND_net), .I1(n18376[12]), .I2(n1047_adj_4472), 
            .I3(n51692), .O(n17896[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_15 (.CI(n51692), .I0(n18376[12]), .I1(n1047_adj_4472), 
            .CO(n51693));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[6]), 
            .I3(n51307), .O(n382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_3 (.CI(n52239), .I0(n20392[0]), .I1(n195), .CO(n52240));
    SB_LUT4 add_4990_14_lut (.I0(GND_net), .I1(n18376[11]), .I2(n974_adj_4474), 
            .I3(n51691), .O(n17896[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_14 (.CI(n51691), .I0(n18376[11]), .I1(n974_adj_4474), 
            .CO(n51692));
    SB_CARRY unary_minus_20_add_3_8 (.CI(n51307), .I0(GND_net), .I1(n1_adj_4981[6]), 
            .CO(n51308));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[5]), 
            .I3(n51306), .O(n382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5166_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20280[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4990_13_lut (.I0(GND_net), .I1(n18376[10]), .I2(n901_adj_4476), 
            .I3(n51690), .O(n17896[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_13 (.CI(n51690), .I0(n18376[10]), .I1(n901_adj_4476), 
            .CO(n51691));
    SB_CARRY unary_minus_20_add_3_7 (.CI(n51306), .I0(GND_net), .I1(n1_adj_4981[5]), 
            .CO(n51307));
    SB_CARRY add_5166_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n52239));
    SB_LUT4 add_4990_12_lut (.I0(GND_net), .I1(n18376[9]), .I2(n828_adj_4477), 
            .I3(n51689), .O(n17896[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_12 (.CI(n51689), .I0(n18376[9]), .I1(n828_adj_4477), 
            .CO(n51690));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[4]), 
            .I3(n51305), .O(n382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n51305), .I0(GND_net), .I1(n1_adj_4981[4]), 
            .CO(n51306));
    SB_LUT4 add_5033_15_lut (.I0(GND_net), .I1(n18991[12]), .I2(n1050), 
            .I3(n52238), .O(n18600[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4990_11_lut (.I0(GND_net), .I1(n18376[8]), .I2(n755_adj_4479), 
            .I3(n51688), .O(n17896[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_11 (.CI(n51688), .I0(n18376[8]), .I1(n755_adj_4479), 
            .CO(n51689));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[3]), 
            .I3(n51304), .O(n382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5033_14_lut (.I0(GND_net), .I1(n18991[11]), .I2(n977), 
            .I3(n52237), .O(n18600[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4990_10_lut (.I0(GND_net), .I1(n18376[7]), .I2(n682_adj_4481), 
            .I3(n51687), .O(n17896[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_10 (.CI(n51687), .I0(n18376[7]), .I1(n682_adj_4481), 
            .CO(n51688));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n51304), .I0(GND_net), .I1(n1_adj_4981[3]), 
            .CO(n51305));
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[2]), 
            .I3(n51303), .O(n382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_14 (.CI(n52237), .I0(n18991[11]), .I1(n977), .CO(n52238));
    SB_LUT4 add_4990_9_lut (.I0(GND_net), .I1(n18376[6]), .I2(n609_adj_4483), 
            .I3(n51686), .O(n17896[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_9 (.CI(n51686), .I0(n18376[6]), .I1(n609_adj_4483), 
            .CO(n51687));
    SB_CARRY unary_minus_20_add_3_4 (.CI(n51303), .I0(GND_net), .I1(n1_adj_4981[2]), 
            .CO(n51304));
    SB_LUT4 add_5033_13_lut (.I0(GND_net), .I1(n18991[10]), .I2(n904), 
            .I3(n52236), .O(n18600[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4990_8_lut (.I0(GND_net), .I1(n18376[5]), .I2(n536_adj_4484), 
            .I3(n51685), .O(n17896[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_8 (.CI(n51685), .I0(n18376[5]), .I1(n536_adj_4484), 
            .CO(n51686));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4981[1]), 
            .I3(n51302), .O(n382[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n51302), .I0(GND_net), .I1(n1_adj_4981[1]), 
            .CO(n51303));
    SB_CARRY add_5033_13 (.CI(n52236), .I0(n18991[10]), .I1(n904), .CO(n52237));
    SB_LUT4 add_5033_12_lut (.I0(GND_net), .I1(n18991[9]), .I2(n831), 
            .I3(n52235), .O(n18600[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_12 (.CI(n52235), .I0(n18991[9]), .I1(n831), .CO(n52236));
    SB_LUT4 add_5033_11_lut (.I0(GND_net), .I1(n18991[8]), .I2(n758), 
            .I3(n52234), .O(n18600[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_11 (.CI(n52234), .I0(n18991[8]), .I1(n758), .CO(n52235));
    SB_LUT4 add_5033_10_lut (.I0(GND_net), .I1(n18991[7]), .I2(n685), 
            .I3(n52233), .O(n18600[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_10 (.CI(n52233), .I0(n18991[7]), .I1(n685), .CO(n52234));
    SB_LUT4 add_5033_9_lut (.I0(GND_net), .I1(n18991[6]), .I2(n612), .I3(n52232), 
            .O(n18600[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_9 (.CI(n52232), .I0(n18991[6]), .I1(n612), .CO(n52233));
    SB_LUT4 add_5033_8_lut (.I0(GND_net), .I1(n18991[5]), .I2(n539), .I3(n52231), 
            .O(n18600[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_8 (.CI(n52231), .I0(n18991[5]), .I1(n539), .CO(n52232));
    SB_LUT4 add_5033_7_lut (.I0(GND_net), .I1(n18991[4]), .I2(n466), .I3(n52230), 
            .O(n18600[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_7 (.CI(n52230), .I0(n18991[4]), .I1(n466), .CO(n52231));
    SB_LUT4 add_5033_6_lut (.I0(GND_net), .I1(n18991[3]), .I2(n393_adj_4486), 
            .I3(n52229), .O(n18600[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_6 (.CI(n52229), .I0(n18991[3]), .I1(n393_adj_4486), 
            .CO(n52230));
    SB_LUT4 add_5033_5_lut (.I0(GND_net), .I1(n18991[2]), .I2(n320), .I3(n52228), 
            .O(n18600[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_5 (.CI(n52228), .I0(n18991[2]), .I1(n320), .CO(n52229));
    SB_LUT4 add_5033_4_lut (.I0(GND_net), .I1(n18991[1]), .I2(n247), .I3(n52227), 
            .O(n18600[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_4 (.CI(n52227), .I0(n18991[1]), .I1(n247), .CO(n52228));
    SB_LUT4 add_5033_3_lut (.I0(GND_net), .I1(n18991[0]), .I2(n174), .I3(n52226), 
            .O(n18600[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_3 (.CI(n52226), .I0(n18991[0]), .I1(n174), .CO(n52227));
    SB_LUT4 add_5033_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n18600[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n52226));
    SB_LUT4 add_5059_14_lut (.I0(GND_net), .I1(n19328[11]), .I2(n980), 
            .I3(n52225), .O(n18991[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5059_13_lut (.I0(GND_net), .I1(n19328[10]), .I2(n907), 
            .I3(n52224), .O(n18991[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_13 (.CI(n52224), .I0(n19328[10]), .I1(n907), .CO(n52225));
    SB_LUT4 add_5059_12_lut (.I0(GND_net), .I1(n19328[9]), .I2(n834), 
            .I3(n52223), .O(n18991[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_12 (.CI(n52223), .I0(n19328[9]), .I1(n834), .CO(n52224));
    SB_LUT4 LessThan_21_i21_rep_90_2_lut (.I0(n356[10]), .I1(n382[10]), 
            .I2(GND_net), .I3(GND_net), .O(n69107));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i21_rep_90_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5059_11_lut (.I0(GND_net), .I1(n19328[8]), .I2(n761), 
            .I3(n52222), .O(n18991[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_11 (.CI(n52222), .I0(n19328[8]), .I1(n761), .CO(n52223));
    SB_LUT4 add_5059_10_lut (.I0(GND_net), .I1(n19328[7]), .I2(n688), 
            .I3(n52221), .O(n18991[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_10 (.CI(n52221), .I0(n19328[7]), .I1(n688), .CO(n52222));
    SB_LUT4 add_5059_9_lut (.I0(GND_net), .I1(n19328[6]), .I2(n615), .I3(n52220), 
            .O(n18991[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_9 (.CI(n52220), .I0(n19328[6]), .I1(n615), .CO(n52221));
    SB_LUT4 add_5059_8_lut (.I0(GND_net), .I1(n19328[5]), .I2(n542), .I3(n52219), 
            .O(n18991[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_8 (.CI(n52219), .I0(n19328[5]), .I1(n542), .CO(n52220));
    SB_LUT4 add_5059_7_lut (.I0(GND_net), .I1(n19328[4]), .I2(n469), .I3(n52218), 
            .O(n18991[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_7 (.CI(n52218), .I0(n19328[4]), .I1(n469), .CO(n52219));
    SB_LUT4 add_5059_6_lut (.I0(GND_net), .I1(n19328[3]), .I2(n396_adj_4487), 
            .I3(n52217), .O(n18991[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_6 (.CI(n52217), .I0(n19328[3]), .I1(n396_adj_4487), 
            .CO(n52218));
    SB_LUT4 add_5059_5_lut (.I0(GND_net), .I1(n19328[2]), .I2(n323), .I3(n52216), 
            .O(n18991[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_5 (.CI(n52216), .I0(n19328[2]), .I1(n323), .CO(n52217));
    SB_LUT4 add_5059_4_lut (.I0(GND_net), .I1(n19328[1]), .I2(n250), .I3(n52215), 
            .O(n18991[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_4 (.CI(n52215), .I0(n19328[1]), .I1(n250), .CO(n52216));
    SB_LUT4 add_5059_3_lut (.I0(GND_net), .I1(n19328[0]), .I2(n177), .I3(n52214), 
            .O(n18991[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_3 (.CI(n52214), .I0(n19328[0]), .I1(n177), .CO(n52215));
    SB_LUT4 add_5059_2_lut (.I0(GND_net), .I1(n35_c), .I2(n104), .I3(GND_net), 
            .O(n18991[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_2 (.CI(GND_net), .I0(n35_c), .I1(n104), .CO(n52214));
    SB_LUT4 add_5179_7_lut (.I0(GND_net), .I1(n60196), .I2(n490), .I3(n52213), 
            .O(n20392[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_6_lut (.I0(GND_net), .I1(n20476[3]), .I2(n417), .I3(n52212), 
            .O(n20392[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_6 (.CI(n52212), .I0(n20476[3]), .I1(n417), .CO(n52213));
    SB_LUT4 add_5179_5_lut (.I0(GND_net), .I1(n20476[2]), .I2(n344), .I3(n52211), 
            .O(n20392[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_5 (.CI(n52211), .I0(n20476[2]), .I1(n344), .CO(n52212));
    SB_LUT4 add_5179_4_lut (.I0(GND_net), .I1(n20476[1]), .I2(n271), .I3(n52210), 
            .O(n20392[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_4 (.CI(n52210), .I0(n20476[1]), .I1(n271), .CO(n52211));
    SB_LUT4 add_5179_3_lut (.I0(GND_net), .I1(n20476[0]), .I2(n198), .I3(n52209), 
            .O(n20392[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_3 (.CI(n52209), .I0(n20476[0]), .I1(n198), .CO(n52210));
    SB_LUT4 add_5179_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20392[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n52209));
    SB_LUT4 add_5083_13_lut (.I0(GND_net), .I1(n19615[10]), .I2(n910), 
            .I3(n52208), .O(n19328[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_12_lut (.I0(GND_net), .I1(n19615[9]), .I2(n837), 
            .I3(n52207), .O(n19328[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_12 (.CI(n52207), .I0(n19615[9]), .I1(n837), .CO(n52208));
    SB_LUT4 add_5083_11_lut (.I0(GND_net), .I1(n19615[8]), .I2(n764), 
            .I3(n52206), .O(n19328[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_11 (.CI(n52206), .I0(n19615[8]), .I1(n764), .CO(n52207));
    SB_LUT4 i50180_4_lut (.I0(n356[11]), .I1(n69107), .I2(n382[11]), .I3(n67202), 
            .O(n67196));
    defparam i50180_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_5083_10_lut (.I0(GND_net), .I1(n19615[7]), .I2(n691), 
            .I3(n52205), .O(n19328[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_10 (.CI(n52205), .I0(n19615[7]), .I1(n691), .CO(n52206));
    SB_LUT4 add_5083_9_lut (.I0(GND_net), .I1(n19615[6]), .I2(n618), .I3(n52204), 
            .O(n19328[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_9 (.CI(n52204), .I0(n19615[6]), .I1(n618), .CO(n52205));
    SB_LUT4 add_5083_8_lut (.I0(GND_net), .I1(n19615[5]), .I2(n545), .I3(n52203), 
            .O(n19328[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_8 (.CI(n52203), .I0(n19615[5]), .I1(n545), .CO(n52204));
    SB_LUT4 add_5083_7_lut (.I0(GND_net), .I1(n19615[4]), .I2(n472), .I3(n52202), 
            .O(n19328[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_7 (.CI(n52202), .I0(n19615[4]), .I1(n472), .CO(n52203));
    SB_LUT4 add_5083_6_lut (.I0(GND_net), .I1(n19615[3]), .I2(n399_adj_4488), 
            .I3(n52201), .O(n19328[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_6 (.CI(n52201), .I0(n19615[3]), .I1(n399_adj_4488), 
            .CO(n52202));
    SB_LUT4 add_5083_5_lut (.I0(GND_net), .I1(n19615[2]), .I2(n326), .I3(n52200), 
            .O(n19328[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_5 (.CI(n52200), .I0(n19615[2]), .I1(n326), .CO(n52201));
    SB_LUT4 add_5083_4_lut (.I0(GND_net), .I1(n19615[1]), .I2(n253), .I3(n52199), 
            .O(n19328[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_4 (.CI(n52199), .I0(n19615[1]), .I1(n253), .CO(n52200));
    SB_LUT4 add_5083_3_lut (.I0(GND_net), .I1(n19615[0]), .I2(n180), .I3(n52198), 
            .O(n19328[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_3 (.CI(n52198), .I0(n19615[0]), .I1(n180), .CO(n52199));
    SB_LUT4 add_5083_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n19328[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i25_rep_85_2_lut (.I0(n356[12]), .I1(n382[12]), 
            .I2(GND_net), .I3(GND_net), .O(n69102));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i25_rep_85_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5083_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n52198));
    SB_LUT4 add_5105_12_lut (.I0(GND_net), .I1(n19856[9]), .I2(n840), 
            .I3(n52197), .O(n19615[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n382[9]), .I1(n382[21]), .I2(n356[21]), 
            .I3(GND_net), .O(n16_adj_4489));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5105_11_lut (.I0(GND_net), .I1(n19856[8]), .I2(n767), 
            .I3(n52196), .O(n19615[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_11 (.CI(n52196), .I0(n19856[8]), .I1(n767), .CO(n52197));
    SB_LUT4 add_5105_10_lut (.I0(GND_net), .I1(n19856[7]), .I2(n694), 
            .I3(n52195), .O(n19615[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_10 (.CI(n52195), .I0(n19856[7]), .I1(n694), .CO(n52196));
    SB_LUT4 add_5105_9_lut (.I0(GND_net), .I1(n19856[6]), .I2(n621), .I3(n52194), 
            .O(n19615[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_9 (.CI(n52194), .I0(n19856[6]), .I1(n621), .CO(n52195));
    SB_LUT4 add_5105_8_lut (.I0(GND_net), .I1(n19856[5]), .I2(n548), .I3(n52193), 
            .O(n19615[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_8 (.CI(n52193), .I0(n19856[5]), .I1(n548), .CO(n52194));
    SB_LUT4 add_5105_7_lut (.I0(GND_net), .I1(n19856[4]), .I2(n475), .I3(n52192), 
            .O(n19615[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_7 (.CI(n52192), .I0(n19856[4]), .I1(n475), .CO(n52193));
    SB_LUT4 add_5105_6_lut (.I0(GND_net), .I1(n19856[3]), .I2(n402_adj_4490), 
            .I3(n52191), .O(n19615[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_6 (.CI(n52191), .I0(n19856[3]), .I1(n402_adj_4490), 
            .CO(n52192));
    SB_LUT4 add_5105_5_lut (.I0(GND_net), .I1(n19856[2]), .I2(n329), .I3(n52190), 
            .O(n19615[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_5 (.CI(n52190), .I0(n19856[2]), .I1(n329), .CO(n52191));
    SB_LUT4 add_5105_4_lut (.I0(GND_net), .I1(n19856[1]), .I2(n256), .I3(n52189), 
            .O(n19615[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_4 (.CI(n52189), .I0(n19856[1]), .I1(n256), .CO(n52190));
    SB_LUT4 add_5105_3_lut (.I0(GND_net), .I1(n19856[0]), .I2(n183), .I3(n52188), 
            .O(n19615[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_3 (.CI(n52188), .I0(n19856[0]), .I1(n183), .CO(n52189));
    SB_LUT4 add_5105_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n19615[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n52188));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n39319), .I1(GND_net), .I2(n1_adj_4981[0]), 
            .I3(VCC_net), .O(n65413)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4981[0]), 
            .CO(n51302));
    SB_LUT4 add_4990_7_lut (.I0(GND_net), .I1(n18376[4]), .I2(n463_adj_4492), 
            .I3(n51684), .O(n17896[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_7 (.CI(n51684), .I0(n18376[4]), .I1(n463_adj_4492), 
            .CO(n51685));
    SB_LUT4 add_4990_6_lut (.I0(GND_net), .I1(n18376[3]), .I2(n390_adj_4493), 
            .I3(n51683), .O(n17896[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_6 (.CI(n51683), .I0(n18376[3]), .I1(n390_adj_4493), 
            .CO(n51684));
    SB_LUT4 add_4990_5_lut (.I0(GND_net), .I1(n18376[2]), .I2(n317_adj_4494), 
            .I3(n51682), .O(n17896[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_5 (.CI(n51682), .I0(n18376[2]), .I1(n317_adj_4494), 
            .CO(n51683));
    SB_LUT4 add_4990_4_lut (.I0(GND_net), .I1(n18376[1]), .I2(n244_adj_4495), 
            .I3(n51681), .O(n17896[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_4 (.CI(n51681), .I0(n18376[1]), .I1(n244_adj_4495), 
            .CO(n51682));
    SB_LUT4 add_4990_3_lut (.I0(GND_net), .I1(n18376[0]), .I2(n171_adj_4496), 
            .I3(n51680), .O(n17896[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_3 (.CI(n51680), .I0(n18376[0]), .I1(n171_adj_4496), 
            .CO(n51681));
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[23]), 
            .I3(n51301), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4990_2_lut (.I0(GND_net), .I1(n29_adj_4499), .I2(n98_adj_4500), 
            .I3(GND_net), .O(n17896[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4990_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4990_2 (.CI(GND_net), .I0(n29_adj_4499), .I1(n98_adj_4500), 
            .CO(n51680));
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[22]), 
            .I3(n51300), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_15_lut (.I0(GND_net), .I1(n18796[12]), .I2(n1050_adj_4502), 
            .I3(n51679), .O(n18376[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_14_lut (.I0(GND_net), .I1(n18796[11]), .I2(n977_adj_4503), 
            .I3(n51678), .O(n18376[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_24 (.CI(n51300), .I0(GND_net), .I1(n1_adj_4982[22]), 
            .CO(n51301));
    SB_CARRY add_5019_14 (.CI(n51678), .I0(n18796[11]), .I1(n977_adj_4503), 
            .CO(n51679));
    SB_LUT4 add_5019_13_lut (.I0(GND_net), .I1(n18796[10]), .I2(n904_adj_4504), 
            .I3(n51677), .O(n18376[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[21]), 
            .I3(n51299), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_13 (.CI(n51677), .I0(n18796[10]), .I1(n904_adj_4504), 
            .CO(n51678));
    SB_LUT4 add_5019_12_lut (.I0(GND_net), .I1(n18796[9]), .I2(n831_adj_4506), 
            .I3(n51676), .O(n18376[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_12 (.CI(n51676), .I0(n18796[9]), .I1(n831_adj_4506), 
            .CO(n51677));
    SB_LUT4 add_5019_11_lut (.I0(GND_net), .I1(n18796[8]), .I2(n758_adj_4507), 
            .I3(n51675), .O(n18376[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_11 (.CI(n51675), .I0(n18796[8]), .I1(n758_adj_4507), 
            .CO(n51676));
    SB_LUT4 add_5019_10_lut (.I0(GND_net), .I1(n18796[7]), .I2(n685_adj_4508), 
            .I3(n51674), .O(n18376[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_10 (.CI(n51674), .I0(n18796[7]), .I1(n685_adj_4508), 
            .CO(n51675));
    SB_LUT4 add_5019_9_lut (.I0(GND_net), .I1(n18796[6]), .I2(n612_adj_4509), 
            .I3(n51673), .O(n18376[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_9 (.CI(n51673), .I0(n18796[6]), .I1(n612_adj_4509), 
            .CO(n51674));
    SB_CARRY unary_minus_13_add_3_23 (.CI(n51299), .I0(GND_net), .I1(n1_adj_4982[21]), 
            .CO(n51300));
    SB_LUT4 add_5019_8_lut (.I0(GND_net), .I1(n18796[5]), .I2(n539_adj_4510), 
            .I3(n51672), .O(n18376[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_8 (.CI(n51672), .I0(n18796[5]), .I1(n539_adj_4510), 
            .CO(n51673));
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[20]), 
            .I3(n51298), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_22 (.CI(n51298), .I0(GND_net), .I1(n1_adj_4982[20]), 
            .CO(n51299));
    SB_LUT4 add_5019_7_lut (.I0(GND_net), .I1(n18796[4]), .I2(n466_adj_4512), 
            .I3(n51671), .O(n18376[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_7 (.CI(n51671), .I0(n18796[4]), .I1(n466_adj_4512), 
            .CO(n51672));
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[19]), 
            .I3(n51297), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_6_lut (.I0(GND_net), .I1(n18796[3]), .I2(n393_adj_4514), 
            .I3(n51670), .O(n18376[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_6 (.CI(n51670), .I0(n18796[3]), .I1(n393_adj_4514), 
            .CO(n51671));
    SB_CARRY unary_minus_13_add_3_21 (.CI(n51297), .I0(GND_net), .I1(n1_adj_4982[19]), 
            .CO(n51298));
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[18]), 
            .I3(n51296), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_5_lut (.I0(GND_net), .I1(n18796[2]), .I2(n320_adj_4516), 
            .I3(n51669), .O(n18376[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_5 (.CI(n51669), .I0(n18796[2]), .I1(n320_adj_4516), 
            .CO(n51670));
    SB_CARRY unary_minus_13_add_3_20 (.CI(n51296), .I0(GND_net), .I1(n1_adj_4982[18]), 
            .CO(n51297));
    SB_LUT4 add_5019_4_lut (.I0(GND_net), .I1(n18796[1]), .I2(n247_adj_4517), 
            .I3(n51668), .O(n18376[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_4 (.CI(n51668), .I0(n18796[1]), .I1(n247_adj_4517), 
            .CO(n51669));
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[17]), 
            .I3(n51295), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n51295), .I0(GND_net), .I1(n1_adj_4982[17]), 
            .CO(n51296));
    SB_LUT4 add_5019_3_lut (.I0(GND_net), .I1(n18796[0]), .I2(n174_adj_4519), 
            .I3(n51667), .O(n18376[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_3 (.CI(n51667), .I0(n18796[0]), .I1(n174_adj_4519), 
            .CO(n51668));
    SB_LUT4 i49246_4_lut (.I0(n356[21]), .I1(n356[9]), .I2(n382[21]), 
            .I3(n382[9]), .O(n66262));
    defparam i49246_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[16]), 
            .I3(n51294), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_2_lut (.I0(GND_net), .I1(n32_adj_4521), .I2(n101_adj_4522), 
            .I3(GND_net), .O(n18376[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_2 (.CI(GND_net), .I0(n32_adj_4521), .I1(n101_adj_4522), 
            .CO(n51667));
    SB_CARRY unary_minus_13_add_3_18 (.CI(n51294), .I0(GND_net), .I1(n1_adj_4982[16]), 
            .CO(n51295));
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[15]), 
            .I3(n51293), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n51293), .I0(GND_net), .I1(n1_adj_4982[15]), 
            .CO(n51294));
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[14]), 
            .I3(n51292), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_16 (.CI(n51292), .I0(GND_net), .I1(n1_adj_4982[14]), 
            .CO(n51293));
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[13]), 
            .I3(n51291), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n51291), .I0(GND_net), .I1(n1_adj_4982[13]), 
            .CO(n51292));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[12]), 
            .I3(n51290), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n51290), .I0(GND_net), .I1(n1_adj_4982[12]), 
            .CO(n51291));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[11]), 
            .I3(n51289), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49431_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n66460), 
            .O(n66447));
    defparam i49431_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_13_add_3_13 (.CI(n51289), .I0(GND_net), .I1(n1_adj_4982[11]), 
            .CO(n51290));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[10]), 
            .I3(n51288), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n51288), .I0(GND_net), .I1(n1_adj_4982[10]), 
            .CO(n51289));
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[9]), 
            .I3(n51287), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n51287), .I0(GND_net), .I1(n1_adj_4982[9]), 
            .CO(n51288));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[8]), 
            .I3(n51286), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_10 (.CI(n51286), .I0(GND_net), .I1(n1_adj_4982[8]), 
            .CO(n51287));
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[7]), 
            .I3(n51285), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5173_8_lut (.I0(GND_net), .I1(n20440[5]), .I2(n560_adj_4535), 
            .I3(n51650), .O(n20343[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n51285), .I0(GND_net), .I1(n1_adj_4982[7]), 
            .CO(n51286));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[6]), 
            .I3(n51284), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5173_7_lut (.I0(GND_net), .I1(n20440[4]), .I2(n487_adj_4537), 
            .I3(n51649), .O(n20343[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5173_7 (.CI(n51649), .I0(n20440[4]), .I1(n487_adj_4537), 
            .CO(n51650));
    SB_CARRY unary_minus_13_add_3_8 (.CI(n51284), .I0(GND_net), .I1(n1_adj_4982[6]), 
            .CO(n51285));
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[5]), 
            .I3(n51283), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5173_6_lut (.I0(GND_net), .I1(n20440[3]), .I2(n414_adj_4539), 
            .I3(n51648), .O(n20343[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5173_6 (.CI(n51648), .I0(n20440[3]), .I1(n414_adj_4539), 
            .CO(n51649));
    SB_CARRY unary_minus_13_add_3_7 (.CI(n51283), .I0(GND_net), .I1(n1_adj_4982[5]), 
            .CO(n51284));
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[4]), 
            .I3(n51282), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5173_5_lut (.I0(GND_net), .I1(n20440[2]), .I2(n341_adj_4541), 
            .I3(n51647), .O(n20343[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5173_5 (.CI(n51647), .I0(n20440[2]), .I1(n341_adj_4541), 
            .CO(n51648));
    SB_CARRY unary_minus_13_add_3_6 (.CI(n51282), .I0(GND_net), .I1(n1_adj_4982[4]), 
            .CO(n51283));
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[3]), 
            .I3(n51281), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5173_4_lut (.I0(GND_net), .I1(n20440[1]), .I2(n268_adj_4543), 
            .I3(n51646), .O(n20343[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5173_4 (.CI(n51646), .I0(n20440[1]), .I1(n268_adj_4543), 
            .CO(n51647));
    SB_LUT4 add_5173_3_lut (.I0(GND_net), .I1(n20440[0]), .I2(n195_adj_4544), 
            .I3(n51645), .O(n20343[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5173_3 (.CI(n51645), .I0(n20440[0]), .I1(n195_adj_4544), 
            .CO(n51646));
    SB_LUT4 add_5173_2_lut (.I0(GND_net), .I1(n53_adj_4545), .I2(n122_adj_4546), 
            .I3(GND_net), .O(n20343[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5173_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5173_2 (.CI(GND_net), .I0(n53_adj_4545), .I1(n122_adj_4546), 
            .CO(n51645));
    SB_LUT4 add_5046_14_lut (.I0(GND_net), .I1(n19160[11]), .I2(n980_adj_4547), 
            .I3(n51644), .O(n18796[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5046_13_lut (.I0(GND_net), .I1(n19160[10]), .I2(n907_adj_4548), 
            .I3(n51643), .O(n18796[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_13 (.CI(n51643), .I0(n19160[10]), .I1(n907_adj_4548), 
            .CO(n51644));
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n382[4]), .I1(n382[8]), .I2(n356[8]), 
            .I3(GND_net), .O(n8_adj_4549));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5046_12_lut (.I0(GND_net), .I1(n19160[9]), .I2(n834_adj_4550), 
            .I3(n51642), .O(n18796[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_12 (.CI(n51642), .I0(n19160[9]), .I1(n834_adj_4550), 
            .CO(n51643));
    SB_CARRY unary_minus_13_add_3_5 (.CI(n51281), .I0(GND_net), .I1(n1_adj_4982[3]), 
            .CO(n51282));
    SB_LUT4 add_5046_11_lut (.I0(GND_net), .I1(n19160[8]), .I2(n761_adj_4551), 
            .I3(n51641), .O(n18796[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[2]), 
            .I3(n51280), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_11 (.CI(n51641), .I0(n19160[8]), .I1(n761_adj_4551), 
            .CO(n51642));
    SB_CARRY unary_minus_13_add_3_4 (.CI(n51280), .I0(GND_net), .I1(n1_adj_4982[2]), 
            .CO(n51281));
    SB_LUT4 add_5046_10_lut (.I0(GND_net), .I1(n19160[7]), .I2(n688_adj_4553), 
            .I3(n51640), .O(n18796[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[1]), 
            .I3(n51279), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_10 (.CI(n51640), .I0(n19160[7]), .I1(n688_adj_4553), 
            .CO(n51641));
    SB_CARRY unary_minus_13_add_3_3 (.CI(n51279), .I0(GND_net), .I1(n1_adj_4982[1]), 
            .CO(n51280));
    SB_LUT4 add_5046_9_lut (.I0(GND_net), .I1(n19160[6]), .I2(n615_adj_4555), 
            .I3(n51639), .O(n18796[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4982[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_9 (.CI(n51639), .I0(n19160[6]), .I1(n615_adj_4555), 
            .CO(n51640));
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4982[0]), 
            .CO(n51279));
    SB_LUT4 add_5046_8_lut (.I0(GND_net), .I1(n19160[5]), .I2(n542_adj_4557), 
            .I3(n51638), .O(n18796[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_8 (.CI(n51638), .I0(n19160[5]), .I1(n542_adj_4557), 
            .CO(n51639));
    SB_LUT4 add_5046_7_lut (.I0(GND_net), .I1(n19160[4]), .I2(n469_adj_4558), 
            .I3(n51637), .O(n18796[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_7 (.CI(n51637), .I0(n19160[4]), .I1(n469_adj_4558), 
            .CO(n51638));
    SB_LUT4 add_5046_6_lut (.I0(GND_net), .I1(n19160[3]), .I2(n396_adj_4559), 
            .I3(n51636), .O(n18796[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_6 (.CI(n51636), .I0(n19160[3]), .I1(n396_adj_4559), 
            .CO(n51637));
    SB_LUT4 add_5046_5_lut (.I0(GND_net), .I1(n19160[2]), .I2(n323_adj_4560), 
            .I3(n51635), .O(n18796[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_5 (.CI(n51635), .I0(n19160[2]), .I1(n323_adj_4560), 
            .CO(n51636));
    SB_LUT4 add_5046_4_lut (.I0(GND_net), .I1(n19160[1]), .I2(n250_adj_4561), 
            .I3(n51634), .O(n18796[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_4 (.CI(n51634), .I0(n19160[1]), .I1(n250_adj_4561), 
            .CO(n51635));
    SB_LUT4 add_5046_3_lut (.I0(GND_net), .I1(n19160[0]), .I2(n177_adj_4562), 
            .I3(n51633), .O(n18796[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_3 (.CI(n51633), .I0(n19160[0]), .I1(n177_adj_4562), 
            .CO(n51634));
    SB_LUT4 add_5046_2_lut (.I0(GND_net), .I1(n35_adj_4563), .I2(n104_adj_4564), 
            .I3(GND_net), .O(n18796[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_4489), .I1(n382[22]), .I2(n356[22]), 
            .I3(GND_net), .O(n24_adj_4565));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5046_2 (.CI(GND_net), .I0(n35_adj_4563), .I1(n104_adj_4564), 
            .CO(n51633));
    SB_LUT4 i51153_4_lut (.I0(n30), .I1(n10_adj_4566), .I2(n35_adj_4567), 
            .I3(n66444), .O(n68169));   // verilog/motorControl.v(51[12:29])
    defparam i51153_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49404_4_lut (.I0(n356[3]), .I1(n356[2]), .I2(n382[3]), .I3(n382[2]), 
            .O(n66420));
    defparam i49404_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i9_rep_83_2_lut (.I0(n356[4]), .I1(n382[4]), .I2(GND_net), 
            .I3(GND_net), .O(n69100));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i9_rep_83_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49402_4_lut (.I0(n356[5]), .I1(n69100), .I2(n382[5]), .I3(n66420), 
            .O(n66418));
    defparam i49402_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4568));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i13_rep_111_2_lut (.I0(n356[6]), .I1(n382[6]), .I2(GND_net), 
            .I3(GND_net), .O(n69128));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i13_rep_111_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50573_4_lut (.I0(n356[7]), .I1(n69128), .I2(n382[7]), .I3(n66418), 
            .O(n67589));
    defparam i50573_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i17_rep_108_2_lut (.I0(n356[8]), .I1(n382[8]), .I2(GND_net), 
            .I3(GND_net), .O(n69125));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i17_rep_108_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50190_4_lut (.I0(n356[9]), .I1(n69125), .I2(n382[9]), .I3(n67589), 
            .O(n67206));
    defparam i50190_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i50899_4_lut (.I0(n356[11]), .I1(n69107), .I2(n382[11]), .I3(n67206), 
            .O(n67915));
    defparam i50899_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4569));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4570));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n20560[2]), .I1(n6_adj_4571), .I2(\Kp[4] ), 
            .I3(n49[18]), .O(n20511[3]));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 counter_1936_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n52123), .O(n51[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n52122), .O(n51[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(23[10] 30[6])
    SB_LUT4 i49346_4_lut (.I0(n356[13]), .I1(n69102), .I2(n382[13]), .I3(n67915), 
            .O(n66362));
    defparam i49346_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY counter_1936_add_4_32 (.CI(n52122), .I0(GND_net), .I1(counter[30]), 
            .CO(n52123));
    SB_LUT4 counter_1936_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n52121), .O(n51[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_31 (.CI(n52121), .I0(GND_net), .I1(counter[29]), 
            .CO(n52122));
    SB_LUT4 counter_1936_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n52120), .O(n51[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5071_13_lut (.I0(GND_net), .I1(n19472[10]), .I2(n910_adj_4574), 
            .I3(n51617), .O(n19160[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5071_12_lut (.I0(GND_net), .I1(n19472[9]), .I2(n837_adj_4575), 
            .I3(n51616), .O(n19160[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_30 (.CI(n52120), .I0(GND_net), .I1(counter[28]), 
            .CO(n52121));
    SB_LUT4 counter_1936_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n52119), .O(n51[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_29 (.CI(n52119), .I0(GND_net), .I1(counter[27]), 
            .CO(n52120));
    SB_CARRY add_5071_12 (.CI(n51616), .I0(n19472[9]), .I1(n837_adj_4575), 
            .CO(n51617));
    SB_LUT4 add_5071_11_lut (.I0(GND_net), .I1(n19472[8]), .I2(n764_adj_4576), 
            .I3(n51615), .O(n19160[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n52118), .O(n51[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_11 (.CI(n51615), .I0(n19472[8]), .I1(n764_adj_4576), 
            .CO(n51616));
    SB_CARRY counter_1936_add_4_28 (.CI(n52118), .I0(GND_net), .I1(counter[26]), 
            .CO(n52119));
    SB_LUT4 add_5071_10_lut (.I0(GND_net), .I1(n19472[7]), .I2(n691_adj_4577), 
            .I3(n51614), .O(n19160[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i29_rep_73_2_lut (.I0(n356[14]), .I1(n382[14]), 
            .I2(GND_net), .I3(GND_net), .O(n69090));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i29_rep_73_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 counter_1936_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n52117), .O(n51[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_10 (.CI(n51614), .I0(n19472[7]), .I1(n691_adj_4577), 
            .CO(n51615));
    SB_LUT4 add_5071_9_lut (.I0(GND_net), .I1(n19472[6]), .I2(n618_adj_4578), 
            .I3(n51613), .O(n19160[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50555_4_lut (.I0(n356[15]), .I1(n69090), .I2(n382[15]), .I3(n66362), 
            .O(n67571));
    defparam i50555_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY counter_1936_add_4_27 (.CI(n52117), .I0(GND_net), .I1(counter[25]), 
            .CO(n52118));
    SB_LUT4 LessThan_21_i33_rep_101_2_lut (.I0(n356[16]), .I1(n382[16]), 
            .I2(GND_net), .I3(GND_net), .O(n69118));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i33_rep_101_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5071_9 (.CI(n51613), .I0(n19472[6]), .I1(n618_adj_4578), 
            .CO(n51614));
    SB_LUT4 counter_1936_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n52116), .O(n51[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5071_8_lut (.I0(GND_net), .I1(n19472[5]), .I2(n545_adj_4579), 
            .I3(n51612), .O(n19160[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_26 (.CI(n52116), .I0(GND_net), .I1(counter[24]), 
            .CO(n52117));
    SB_CARRY add_5071_8 (.CI(n51612), .I0(n19472[5]), .I1(n545_adj_4579), 
            .CO(n51613));
    SB_LUT4 counter_1936_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n52115), .O(n51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5071_7_lut (.I0(GND_net), .I1(n19472[4]), .I2(n472_adj_4580), 
            .I3(n51611), .O(n19160[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_7 (.CI(n51611), .I0(n19472[4]), .I1(n472_adj_4580), 
            .CO(n51612));
    SB_LUT4 i51090_4_lut (.I0(n363), .I1(n69118), .I2(n382[17]), .I3(n67571), 
            .O(n68106));
    defparam i51090_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY counter_1936_add_4_25 (.CI(n52115), .I0(GND_net), .I1(counter[23]), 
            .CO(n52116));
    SB_LUT4 add_5071_6_lut (.I0(GND_net), .I1(n19472[3]), .I2(n399_adj_4581), 
            .I3(n51610), .O(n19160[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n52114), .O(n51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_24 (.CI(n52114), .I0(GND_net), .I1(counter[22]), 
            .CO(n52115));
    SB_LUT4 LessThan_21_i37_rep_64_2_lut (.I0(n356[18]), .I1(n382[18]), 
            .I2(GND_net), .I3(GND_net), .O(n69081));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i37_rep_64_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5071_6 (.CI(n51610), .I0(n19472[3]), .I1(n399_adj_4581), 
            .CO(n51611));
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5071_5_lut (.I0(GND_net), .I1(n19472[2]), .I2(n326_adj_4583), 
            .I3(n51609), .O(n19160[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n52113), .O(n51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_5 (.CI(n51609), .I0(n19472[2]), .I1(n326_adj_4583), 
            .CO(n51610));
    SB_LUT4 i51276_4_lut (.I0(n356[19]), .I1(n69081), .I2(n382[19]), .I3(n68106), 
            .O(n68292));
    defparam i51276_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i49622_3_lut (.I0(n67854), .I1(n356[15]), .I2(n31), .I3(GND_net), 
            .O(n66638));   // verilog/motorControl.v(51[12:29])
    defparam i49622_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1936_add_4_23 (.CI(n52113), .I0(GND_net), .I1(counter[21]), 
            .CO(n52114));
    SB_LUT4 add_5071_4_lut (.I0(GND_net), .I1(n19472[1]), .I2(n253_adj_4584), 
            .I3(n51608), .O(n19160[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n52112), .O(n51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_4 (.CI(n51608), .I0(n19472[1]), .I1(n253_adj_4584), 
            .CO(n51609));
    SB_CARRY counter_1936_add_4_22 (.CI(n52112), .I0(GND_net), .I1(counter[20]), 
            .CO(n52113));
    SB_LUT4 counter_1936_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n52111), .O(n51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51288_4_lut (.I0(n66638), .I1(n68169), .I2(n35_adj_4567), 
            .I3(n66447), .O(n68304));   // verilog/motorControl.v(51[12:29])
    defparam i51288_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i41_rep_61_2_lut (.I0(n356[20]), .I1(n382[20]), 
            .I2(GND_net), .I3(GND_net), .O(n69078));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i41_rep_61_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5071_3_lut (.I0(GND_net), .I1(n19472[0]), .I2(n180_adj_4585), 
            .I3(n51607), .O(n19160[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_21 (.CI(n52111), .I0(GND_net), .I1(counter[19]), 
            .CO(n52112));
    SB_LUT4 counter_1936_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n52110), .O(n51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_3 (.CI(n51607), .I0(n19472[0]), .I1(n180_adj_4585), 
            .CO(n51608));
    SB_CARRY counter_1936_add_4_20 (.CI(n52110), .I0(GND_net), .I1(counter[18]), 
            .CO(n52111));
    SB_LUT4 add_5071_2_lut (.I0(GND_net), .I1(n38_adj_4586), .I2(n107_adj_4587), 
            .I3(GND_net), .O(n19160[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_2 (.CI(GND_net), .I0(n38_adj_4586), .I1(n107_adj_4587), 
            .CO(n51607));
    SB_LUT4 add_5185_7_lut (.I0(GND_net), .I1(n60592), .I2(n490_adj_4588), 
            .I3(n51606), .O(n20440[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49444_4_lut (.I0(n27), .I1(n15_adj_4589), .I2(n13_adj_4590), 
            .I3(n11_adj_4591), .O(n66460));
    defparam i49444_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 counter_1936_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n52109), .O(n51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_19 (.CI(n52109), .I0(GND_net), .I1(counter[17]), 
            .CO(n52110));
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4592));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_1936_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n52108), .O(n51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_18 (.CI(n52108), .I0(GND_net), .I1(counter[16]), 
            .CO(n52109));
    SB_LUT4 counter_1936_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n52107), .O(n51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_17 (.CI(n52107), .I0(GND_net), .I1(counter[15]), 
            .CO(n52108));
    SB_LUT4 add_5185_6_lut (.I0(GND_net), .I1(n20511[3]), .I2(n417_adj_4570), 
            .I3(n51605), .O(n20440[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n52106), .O(n51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_16 (.CI(n52106), .I0(GND_net), .I1(counter[14]), 
            .CO(n52107));
    SB_LUT4 counter_1936_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n52105), .O(n51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_6 (.CI(n51605), .I0(n20511[3]), .I1(n417_adj_4570), 
            .CO(n51606));
    SB_CARRY counter_1936_add_4_15 (.CI(n52105), .I0(GND_net), .I1(counter[13]), 
            .CO(n52106));
    SB_LUT4 counter_1936_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n52104), .O(n51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_14 (.CI(n52104), .I0(GND_net), .I1(counter[12]), 
            .CO(n52105));
    SB_LUT4 counter_1936_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n52103), .O(n51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5185_5_lut (.I0(GND_net), .I1(n20511[2]), .I2(n344_adj_4569), 
            .I3(n51604), .O(n20440[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY counter_1936_add_4_13 (.CI(n52103), .I0(GND_net), .I1(counter[11]), 
            .CO(n52104));
    SB_CARRY add_5185_5 (.CI(n51604), .I0(n20511[2]), .I1(n344_adj_4569), 
            .CO(n51605));
    SB_LUT4 add_5185_4_lut (.I0(GND_net), .I1(n20511[1]), .I2(n271_adj_4594), 
            .I3(n51603), .O(n20440[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n52102), .O(n51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_4 (.CI(n51603), .I0(n20511[1]), .I1(n271_adj_4594), 
            .CO(n51604));
    SB_LUT4 add_5185_3_lut (.I0(GND_net), .I1(n20511[0]), .I2(n198_adj_4595), 
            .I3(n51602), .O(n20440[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_12 (.CI(n52102), .I0(GND_net), .I1(counter[10]), 
            .CO(n52103));
    SB_LUT4 counter_1936_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n52101), .O(n51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_3 (.CI(n51602), .I0(n20511[0]), .I1(n198_adj_4595), 
            .CO(n51603));
    SB_CARRY counter_1936_add_4_11 (.CI(n52101), .I0(GND_net), .I1(counter[9]), 
            .CO(n52102));
    SB_LUT4 add_5185_2_lut (.I0(GND_net), .I1(n56_adj_4596), .I2(n125_adj_4597), 
            .I3(GND_net), .O(n20440[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5185_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1936_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n52100), .O(n51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5185_2 (.CI(GND_net), .I0(n56_adj_4596), .I1(n125_adj_4597), 
            .CO(n51602));
    SB_CARRY counter_1936_add_4_10 (.CI(n52100), .I0(GND_net), .I1(counter[8]), 
            .CO(n52101));
    SB_LUT4 counter_1936_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n52099), .O(n51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_9 (.CI(n52099), .I0(GND_net), .I1(counter[7]), 
            .CO(n52100));
    SB_LUT4 counter_1936_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n52098), .O(n51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_8 (.CI(n52098), .I0(GND_net), .I1(counter[6]), 
            .CO(n52099));
    SB_LUT4 counter_1936_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n52097), .O(n51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51289_3_lut (.I0(n68304), .I1(n356[18]), .I2(n37_adj_4598), 
            .I3(GND_net), .O(n68305));   // verilog/motorControl.v(51[12:29])
    defparam i51289_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1936_add_4_7 (.CI(n52097), .I0(GND_net), .I1(counter[5]), 
            .CO(n52098));
    SB_LUT4 counter_1936_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n52096), .O(n51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_6 (.CI(n52096), .I0(GND_net), .I1(counter[4]), 
            .CO(n52097));
    SB_LUT4 counter_1936_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n52095), .O(n51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_5 (.CI(n52095), .I0(GND_net), .I1(counter[3]), 
            .CO(n52096));
    SB_LUT4 counter_1936_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n52094), .O(n51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_4590), 
            .I3(GND_net), .O(n10_adj_4566));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1936_add_4_4 (.CI(n52094), .I0(GND_net), .I1(counter[2]), 
            .CO(n52095));
    SB_LUT4 counter_1936_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n52093), .O(n51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1936_add_4_3 (.CI(n52093), .I0(GND_net), .I1(counter[1]), 
            .CO(n52094));
    SB_LUT4 counter_1936_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1936_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i138_2_lut (.I0(\Kp[2] ), .I1(n49[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204_adj_4600));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35273_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n49[22]), .I3(n49[21]), 
            .O(n20608[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35273_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i89_2_lut (.I0(\Kp[1] ), .I1(n49[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i42_2_lut (.I0(\Kp[0] ), .I1(n49[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1936_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52093));
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4588));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_4592), .I1(n363), .I2(n35_adj_4567), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_945 (.I0(\Kp[4] ), .I1(\Kp[5] ), .I2(n49[19]), 
            .I3(n49[18]), .O(n62070));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_3_lut (.I0(\Kp[3] ), .I1(n62070), .I2(n49[20]), .I3(GND_net), 
            .O(n62072));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i142_2_lut (.I0(\Kp[2] ), .I1(n49[21]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\Kp[1] ), .I1(n210), .I2(n49[22]), .I3(n62072), 
            .O(n62076));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h936c;
    SB_LUT4 i35275_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n49[22]), .I3(n49[21]), 
            .O(n50901));   // verilog/motorControl.v(50[18:24])
    defparam i35275_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_947 (.I0(n50901), .I1(\Kp[0] ), .I2(n62076), 
            .I3(n49[23]), .O(n62080));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h695a;
    SB_LUT4 i35233_4_lut (.I0(n20560[2]), .I1(\Kp[4] ), .I2(n6_adj_4571), 
            .I3(n49[18]), .O(n8_adj_4602));   // verilog/motorControl.v(50[18:24])
    defparam i35233_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n6_adj_4603), .I1(n8_adj_4602), .I2(n4_adj_4604), 
            .I3(n62080), .O(n60592));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i51261_3_lut (.I0(n68305), .I1(n356[19]), .I2(n39_adj_4605), 
            .I3(GND_net), .O(n68277));   // verilog/motorControl.v(51[12:29])
    defparam i51261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n207[12]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i13_3_lut (.I0(n207[12]), .I1(IntegralLimit[12]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [12]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4587));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4586));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50262_4_lut (.I0(n13_adj_4590), .I1(n11_adj_4591), .I2(n9_adj_4608), 
            .I3(n65598), .O(n67278));
    defparam i50262_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[19]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49420_4_lut (.I0(n43_adj_4609), .I1(n41_adj_4610), .I2(n39_adj_4605), 
            .I3(n68219), .O(n66436));
    defparam i49420_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50256_4_lut (.I0(n19_adj_4611), .I1(n17_adj_4612), .I2(n15_adj_4589), 
            .I3(n67278), .O(n67272));
    defparam i50256_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51108_4_lut (.I0(n25_adj_4613), .I1(n23_adj_4614), .I2(n21_adj_4615), 
            .I3(n67272), .O(n68124));
    defparam i51108_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50591_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n68124), 
            .O(n67607));
    defparam i50591_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51203_4_lut (.I0(n37_adj_4598), .I1(n35_adj_4567), .I2(n33), 
            .I3(n67607), .O(n68219));
    defparam i51203_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50839_3_lut (.I0(n6_adj_4616), .I1(n356[10]), .I2(n21_adj_4615), 
            .I3(GND_net), .O(n67855));   // verilog/motorControl.v(51[12:29])
    defparam i50839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_4609), 
            .I3(GND_net), .O(n16_adj_4617));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_4612), 
            .I3(GND_net), .O(n8_adj_4618));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_4617), .I1(n356[22]), .I2(n45_adj_4619), 
            .I3(GND_net), .O(n24_adj_4620));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49459_4_lut (.I0(n21_adj_4615), .I1(n19_adj_4611), .I2(n17_adj_4612), 
            .I3(n9_adj_4608), .O(n66475));
    defparam i49459_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50840_3_lut (.I0(n67855), .I1(n356[11]), .I2(n23_adj_4614), 
            .I3(GND_net), .O(n67856));   // verilog/motorControl.v(51[12:29])
    defparam i50840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49416_4_lut (.I0(n43_adj_4609), .I1(n25_adj_4613), .I2(n23_adj_4614), 
            .I3(n66475), .O(n66432));
    defparam i49416_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50646_4_lut (.I0(n24_adj_4620), .I1(n8_adj_4618), .I2(n45_adj_4619), 
            .I3(n66426), .O(n67662));   // verilog/motorControl.v(51[12:29])
    defparam i50646_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49620_3_lut (.I0(n67856), .I1(n356[12]), .I2(n25_adj_4613), 
            .I3(GND_net), .O(n66636));   // verilog/motorControl.v(51[12:29])
    defparam i49620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n382[7]), .I1(n382[16]), .I2(n356[16]), 
            .I3(GND_net), .O(n12_adj_4621));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i4_3_lut (.I0(n65413), .I1(n382[1]), .I2(n356[1]), 
            .I3(GND_net), .O(n4_adj_4622));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50831_3_lut (.I0(n4_adj_4622), .I1(n382[13]), .I2(n356[13]), 
            .I3(GND_net), .O(n67847));   // verilog/motorControl.v(51[33:53])
    defparam i50831_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50832_3_lut (.I0(n67847), .I1(n382[14]), .I2(n356[14]), .I3(GND_net), 
            .O(n67848));   // verilog/motorControl.v(51[33:53])
    defparam i50832_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49313_4_lut (.I0(n356[16]), .I1(n356[7]), .I2(n382[16]), 
            .I3(n382[7]), .O(n66329));
    defparam i49313_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i35_rep_96_2_lut (.I0(n363), .I1(n382[17]), .I2(GND_net), 
            .I3(GND_net), .O(n69113));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i35_rep_96_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n382[5]), .I1(n382[6]), .I2(n356[6]), 
            .I3(GND_net), .O(n10_adj_4623));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_4621), .I1(n382[17]), .I2(n363), 
            .I3(GND_net), .O(n30_adj_4624));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5094_12_lut (.I0(GND_net), .I1(n19736[9]), .I2(n840_adj_4625), 
            .I3(n51587), .O(n19472[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5094_11_lut (.I0(GND_net), .I1(n19736[8]), .I2(n767_adj_4626), 
            .I3(n51586), .O(n19472[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_11 (.CI(n51586), .I0(n19736[8]), .I1(n767_adj_4626), 
            .CO(n51587));
    SB_LUT4 add_5094_10_lut (.I0(GND_net), .I1(n19736[7]), .I2(n694_adj_4627), 
            .I3(n51585), .O(n19472[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49315_4_lut (.I0(n356[16]), .I1(n69086), .I2(n382[16]), .I3(n67176), 
            .O(n66331));
    defparam i49315_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_5094_10 (.CI(n51585), .I0(n19736[7]), .I1(n694_adj_4627), 
            .CO(n51586));
    SB_LUT4 add_5094_9_lut (.I0(GND_net), .I1(n19736[6]), .I2(n621_adj_4628), 
            .I3(n51584), .O(n19472[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_9 (.CI(n51584), .I0(n19736[6]), .I1(n621_adj_4628), 
            .CO(n51585));
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5094_8_lut (.I0(GND_net), .I1(n19736[5]), .I2(n548_adj_4630), 
            .I3(n51583), .O(n19472[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_8 (.CI(n51583), .I0(n19736[5]), .I1(n548_adj_4630), 
            .CO(n51584));
    SB_LUT4 add_5094_7_lut (.I0(GND_net), .I1(n19736[4]), .I2(n475_adj_4631), 
            .I3(n51582), .O(n19472[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_7 (.CI(n51582), .I0(n19736[4]), .I1(n475_adj_4631), 
            .CO(n51583));
    SB_LUT4 add_5094_6_lut (.I0(GND_net), .I1(n19736[3]), .I2(n402_adj_4632), 
            .I3(n51581), .O(n19472[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_6 (.CI(n51581), .I0(n19736[3]), .I1(n402_adj_4632), 
            .CO(n51582));
    SB_LUT4 i51122_4_lut (.I0(n66636), .I1(n67662), .I2(n45_adj_4619), 
            .I3(n66432), .O(n68138));   // verilog/motorControl.v(51[12:29])
    defparam i51122_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5094_5_lut (.I0(GND_net), .I1(n19736[2]), .I2(n329_adj_4633), 
            .I3(n51580), .O(n19472[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_5 (.CI(n51580), .I0(n19736[2]), .I1(n329_adj_4633), 
            .CO(n51581));
    SB_LUT4 add_5094_4_lut (.I0(GND_net), .I1(n19736[1]), .I2(n256_adj_4634), 
            .I3(n51579), .O(n19472[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51157_4_lut (.I0(n30_adj_4624), .I1(n10_adj_4623), .I2(n69113), 
            .I3(n66329), .O(n68173));   // verilog/motorControl.v(51[33:53])
    defparam i51157_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5094_4 (.CI(n51579), .I0(n19736[1]), .I1(n256_adj_4634), 
            .CO(n51580));
    SB_LUT4 add_5094_3_lut (.I0(GND_net), .I1(n19736[0]), .I2(n183_adj_4636), 
            .I3(n51578), .O(n19472[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_3 (.CI(n51578), .I0(n19736[0]), .I1(n183_adj_4636), 
            .CO(n51579));
    SB_LUT4 add_5094_2_lut (.I0(GND_net), .I1(n41_adj_4637), .I2(n110_adj_4638), 
            .I3(GND_net), .O(n19472[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5094_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n10755[0]), .I2(n10161[0]), 
            .I3(n51247), .O(n356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n306[22]), 
            .I3(n51246), .O(n356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5094_2 (.CI(GND_net), .I0(n41_adj_4637), .I1(n110_adj_4638), 
            .CO(n51578));
    SB_CARRY add_18_24 (.CI(n51246), .I0(n257[22]), .I1(n306[22]), .CO(n51247));
    SB_LUT4 i49632_3_lut (.I0(n67848), .I1(n382[15]), .I2(n356[15]), .I3(GND_net), 
            .O(n66648));   // verilog/motorControl.v(51[33:53])
    defparam i49632_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n306[21]), 
            .I3(n51245), .O(n356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4585));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49628_3_lut (.I0(n68277), .I1(n356[20]), .I2(n41_adj_4610), 
            .I3(GND_net), .O(n66644));   // verilog/motorControl.v(51[12:29])
    defparam i49628_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_18_23 (.CI(n51245), .I0(n257[21]), .I1(n306[21]), .CO(n51246));
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n306[20]), 
            .I3(n51244), .O(n356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4639));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4430));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4429));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[20]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4428));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4584));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_22 (.CI(n51244), .I0(n257[20]), .I1(n306[20]), .CO(n51245));
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n306[19]), 
            .I3(n51243), .O(n356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_21 (.CI(n51243), .I0(n257[19]), .I1(n306[19]), .CO(n51244));
    SB_LUT4 i51290_4_lut (.I0(n66648), .I1(n68173), .I2(n69113), .I3(n66331), 
            .O(n68306));   // verilog/motorControl.v(51[33:53])
    defparam i51290_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n306[18]), 
            .I3(n51242), .O(n356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51291_3_lut (.I0(n68306), .I1(n382[18]), .I2(n356[18]), .I3(GND_net), 
            .O(n68307));   // verilog/motorControl.v(51[33:53])
    defparam i51291_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_18_20 (.CI(n51242), .I0(n257[18]), .I1(n306[18]), .CO(n51243));
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51124_4_lut (.I0(n66644), .I1(n68138), .I2(n45_adj_4619), 
            .I3(n66436), .O(n68140));   // verilog/motorControl.v(51[12:29])
    defparam i51124_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n306[17]), 
            .I3(n51241), .O(n363)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n51241), .I0(n257[17]), .I1(n306[17]), .CO(n51242));
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4643));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48854_4_lut (.I0(n21_adj_4644), .I1(n19_adj_4645), .I2(n17_adj_4646), 
            .I3(n9_adj_4647), .O(n65870));
    defparam i48854_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48684_4_lut (.I0(n27_adj_4648), .I1(n15_adj_4649), .I2(n13_adj_4650), 
            .I3(n11_adj_4651), .O(n65700));
    defparam i48684_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_4652), 
            .I3(GND_net), .O(n12_adj_4653));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n382[2]), .I1(n382[3]), .I2(n356[3]), 
            .I3(GND_net), .O(n6_adj_4654));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n306[16]), 
            .I3(n51240), .O(n356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50833_3_lut (.I0(n6_adj_4654), .I1(n382[10]), .I2(n356[10]), 
            .I3(GND_net), .O(n67849));   // verilog/motorControl.v(51[33:53])
    defparam i50833_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_18_18 (.CI(n51240), .I0(n257[16]), .I1(n306[16]), .CO(n51241));
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_4650), 
            .I3(GND_net), .O(n10_adj_4656));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_4653), .I1(n182[17]), .I2(n35_adj_4643), 
            .I3(GND_net), .O(n30_adj_4658));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50834_3_lut (.I0(n67849), .I1(n382[11]), .I2(n356[11]), .I3(GND_net), 
            .O(n67850));   // verilog/motorControl.v(51[33:53])
    defparam i50834_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n306[15]), 
            .I3(n51239), .O(n356[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_17 (.CI(n51239), .I0(n257[15]), .I1(n306[15]), .CO(n51240));
    SB_LUT4 i49814_4_lut (.I0(n13_adj_4650), .I1(n11_adj_4651), .I2(n9_adj_4647), 
            .I3(n65914), .O(n66830));
    defparam i49814_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_5115_11_lut (.I0(GND_net), .I1(n19956[8]), .I2(n770), 
            .I3(n51565), .O(n19736[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_10_lut (.I0(GND_net), .I1(n19956[7]), .I2(n697), 
            .I3(n51564), .O(n19736[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [3]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n306[14]), 
            .I3(n51238), .O(n356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_10 (.CI(n51564), .I0(n19956[7]), .I1(n697), .CO(n51565));
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5115_9_lut (.I0(GND_net), .I1(n19956[6]), .I2(n624), .I3(n51563), 
            .O(n19736[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_9 (.CI(n51563), .I0(n19956[6]), .I1(n624), .CO(n51564));
    SB_CARRY add_18_16 (.CI(n51238), .I0(n257[14]), .I1(n306[14]), .CO(n51239));
    SB_LUT4 add_5115_8_lut (.I0(GND_net), .I1(n19956[5]), .I2(n551), .I3(n51562), 
            .O(n19736[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n306[13]), 
            .I3(n51237), .O(n356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_8 (.CI(n51562), .I0(n19956[5]), .I1(n551), .CO(n51563));
    SB_CARRY add_18_15 (.CI(n51237), .I0(n257[13]), .I1(n306[13]), .CO(n51238));
    SB_LUT4 i49790_4_lut (.I0(n19_adj_4645), .I1(n17_adj_4646), .I2(n15_adj_4649), 
            .I3(n66830), .O(n66806));
    defparam i49790_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50957_4_lut (.I0(n25_adj_4661), .I1(n23_adj_4662), .I2(n21_adj_4644), 
            .I3(n66806), .O(n67973));
    defparam i50957_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51128_4_lut (.I0(n66654), .I1(n68142), .I2(n69076), .I3(n66285), 
            .O(n68144));   // verilog/motorControl.v(51[33:53])
    defparam i51128_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50294_4_lut (.I0(n31_adj_4639), .I1(n29_adj_4663), .I2(n27_adj_4648), 
            .I3(n67973), .O(n67310));
    defparam i50294_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49266_4_lut (.I0(n356[21]), .I1(n69102), .I2(n382[21]), .I3(n67196), 
            .O(n66282));
    defparam i49266_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5115_7_lut (.I0(GND_net), .I1(n19956[4]), .I2(n478), .I3(n51561), 
            .O(n19736[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_7 (.CI(n51561), .I0(n19956[4]), .I1(n478), .CO(n51562));
    SB_LUT4 add_5115_6_lut (.I0(GND_net), .I1(n19956[3]), .I2(n405_adj_4665), 
            .I3(n51560), .O(n19736[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_6 (.CI(n51560), .I0(n19956[3]), .I1(n405_adj_4665), 
            .CO(n51561));
    SB_LUT4 i1_4_lut_adj_949 (.I0(n68140), .I1(control_update), .I2(deadband[23]), 
            .I3(n356[23]), .O(n62056));
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h4c04;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n62056), .I1(n68144), .I2(n356[23]), 
            .I3(n47), .O(n61055));
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h0a22;
    SB_LUT4 i51112_4_lut (.I0(n37), .I1(n35_adj_4643), .I2(n33_adj_4652), 
            .I3(n67310), .O(n68128));
    defparam i51112_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4666));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50819_3_lut (.I0(n6_adj_4667), .I1(n182[10]), .I2(n21_adj_4644), 
            .I3(GND_net), .O(n67835));   // verilog/motorControl.v(47[21:44])
    defparam i50819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50820_3_lut (.I0(n67835), .I1(n182[11]), .I2(n23_adj_4662), 
            .I3(GND_net), .O(n67836));   // verilog/motorControl.v(47[21:44])
    defparam i50820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_4646), 
            .I3(GND_net), .O(n8_adj_4668));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_4666), .I1(n182[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4669));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4583));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5115_5_lut (.I0(GND_net), .I1(n19956[2]), .I2(n332_adj_4670), 
            .I3(n51559), .O(n19736[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_5 (.CI(n51559), .I0(n19956[2]), .I1(n332_adj_4670), 
            .CO(n51560));
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n306[12]), 
            .I3(n51236), .O(n356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_14 (.CI(n51236), .I0(n257[12]), .I1(n306[12]), .CO(n51237));
    SB_LUT4 add_5115_4_lut (.I0(GND_net), .I1(n19956[1]), .I2(n259), .I3(n51558), 
            .O(n19736[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5115_4 (.CI(n51558), .I0(n19956[1]), .I1(n259), .CO(n51559));
    SB_LUT4 i48593_4_lut (.I0(n43), .I1(n25_adj_4661), .I2(n23_adj_4662), 
            .I3(n65870), .O(n65609));
    defparam i48593_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50644_4_lut (.I0(n24_adj_4669), .I1(n8_adj_4668), .I2(n45), 
            .I3(n65600), .O(n67660));   // verilog/motorControl.v(47[21:44])
    defparam i50644_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50639_3_lut (.I0(n67836), .I1(n182[12]), .I2(n25_adj_4661), 
            .I3(GND_net), .O(n67655));   // verilog/motorControl.v(47[21:44])
    defparam i50639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_4672));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50817_3_lut (.I0(n4_adj_4672), .I1(n182[13]), .I2(n27_adj_4648), 
            .I3(GND_net), .O(n67833));   // verilog/motorControl.v(47[21:44])
    defparam i50817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n306[11]), 
            .I3(n51235), .O(n356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_13 (.CI(n51235), .I0(n257[11]), .I1(n306[11]), .CO(n51236));
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n306[10]), 
            .I3(n51234), .O(n356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5115_3_lut (.I0(GND_net), .I1(n19956[0]), .I2(n186_adj_4674), 
            .I3(n51557), .O(n19736[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50818_3_lut (.I0(n67833), .I1(n182[14]), .I2(n29_adj_4663), 
            .I3(GND_net), .O(n67834));   // verilog/motorControl.v(47[21:44])
    defparam i50818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48645_4_lut (.I0(n33_adj_4652), .I1(n31_adj_4639), .I2(n29_adj_4663), 
            .I3(n65700), .O(n65661));
    defparam i48645_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51151_4_lut (.I0(n30_adj_4658), .I1(n10_adj_4656), .I2(n35_adj_4643), 
            .I3(n65647), .O(n68167));   // verilog/motorControl.v(47[21:44])
    defparam i51151_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50641_3_lut (.I0(n67834), .I1(n182[15]), .I2(n31_adj_4639), 
            .I3(GND_net), .O(n67657));   // verilog/motorControl.v(47[21:44])
    defparam i50641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51308_4_lut (.I0(n67657), .I1(n68167), .I2(n35_adj_4643), 
            .I3(n65661), .O(n68324));   // verilog/motorControl.v(47[21:44])
    defparam i51308_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5115_3 (.CI(n51557), .I0(n19956[0]), .I1(n186_adj_4674), 
            .CO(n51558));
    SB_LUT4 add_5115_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19736[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5115_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_12 (.CI(n51234), .I0(n257[10]), .I1(n306[10]), .CO(n51235));
    SB_CARRY add_5115_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n51557));
    SB_LUT4 i51309_3_lut (.I0(n68324), .I1(n182[18]), .I2(n37), .I3(GND_net), 
            .O(n68325));   // verilog/motorControl.v(47[21:44])
    defparam i51309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51234_3_lut (.I0(n68325), .I1(n182[19]), .I2(n39), .I3(GND_net), 
            .O(n68250));   // verilog/motorControl.v(47[21:44])
    defparam i51234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48595_4_lut (.I0(n43), .I1(n41_adj_4568), .I2(n39), .I3(n68128), 
            .O(n65611));
    defparam i48595_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50945_4_lut (.I0(n67655), .I1(n67660), .I2(n45), .I3(n65609), 
            .O(n67961));   // verilog/motorControl.v(47[21:44])
    defparam i50945_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51222_3_lut (.I0(n68250), .I1(n182[20]), .I2(n41_adj_4568), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(47[21:44])
    defparam i51222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50947_4_lut (.I0(n40), .I1(n67961), .I2(n45), .I3(n65611), 
            .O(n67963));   // verilog/motorControl.v(47[21:44])
    defparam i50947_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50948_3_lut (.I0(n67963), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(47[21:44])
    defparam i50948_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35406_3_lut_4_lut (.I0(\Kp[2] ), .I1(n49[20]), .I2(n51029), 
            .I3(n20608[0]), .O(n4_adj_4604));   // verilog/motorControl.v(50[18:24])
    defparam i35406_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i50648_4_lut (.I0(n24_adj_4565), .I1(n8_adj_4549), .I2(n69076), 
            .I3(n66262), .O(n67664));   // verilog/motorControl.v(51[33:53])
    defparam i50648_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[2] ), .I1(n49[20]), .I2(n20608[0]), 
            .I3(n51029), .O(n20591[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i35393_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n49[21]), .I2(n49[20]), 
            .I3(\Kp[1] ), .O(n20591[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35393_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i49630_3_lut (.I0(n67850), .I1(n382[12]), .I2(n356[12]), .I3(GND_net), 
            .O(n66646));   // verilog/motorControl.v(51[33:53])
    defparam i49630_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n306[9]), .I3(n51233), 
            .O(n356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_11 (.CI(n51233), .I0(n257[9]), .I1(n306[9]), .CO(n51234));
    SB_LUT4 i35395_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n49[21]), .I2(n49[20]), 
            .I3(\Kp[1] ), .O(n51029));   // verilog/motorControl.v(50[18:24])
    defparam i35395_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n306[8]), .I3(n51232), 
            .O(n356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_10 (.CI(n51232), .I0(n257[8]), .I1(n306[8]), .CO(n51233));
    SB_LUT4 i51259_3_lut (.I0(n68307), .I1(n382[19]), .I2(n356[19]), .I3(GND_net), 
            .O(n68275));   // verilog/motorControl.v(51[33:53])
    defparam i51259_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49269_4_lut (.I0(n356[21]), .I1(n69078), .I2(n382[21]), .I3(n68292), 
            .O(n66285));
    defparam i49269_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i45_rep_59_2_lut (.I0(n356[22]), .I1(n382[22]), 
            .I2(GND_net), .I3(GND_net), .O(n69076));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i45_rep_59_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n306[7]), .I3(n51231), 
            .O(n356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51126_4_lut (.I0(n66646), .I1(n67664), .I2(n69076), .I3(n66282), 
            .O(n68142));   // verilog/motorControl.v(51[33:53])
    defparam i51126_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_18_9 (.CI(n51231), .I0(n257[7]), .I1(n306[7]), .CO(n51232));
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n306[6]), .I3(n51230), 
            .O(n356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4581));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49638_3_lut (.I0(n68275), .I1(n382[20]), .I2(n356[20]), .I3(GND_net), 
            .O(n66654));   // verilog/motorControl.v(51[33:53])
    defparam i49638_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(deadband[0]), .I1(n356[1]), .I2(deadband[1]), 
            .I3(n356[0]), .O(n4_adj_4678));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4580));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35225_3_lut_4_lut (.I0(\Kp[3] ), .I1(n49[18]), .I2(n4_adj_4679), 
            .I3(n20560[1]), .O(n6_adj_4571));   // verilog/motorControl.v(50[18:24])
    defparam i35225_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_951 (.I0(\Kp[3] ), .I1(n49[18]), .I2(n20560[1]), 
            .I3(n4_adj_4679), .O(n20511[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_951.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_952 (.I0(\Kp[2] ), .I1(n49[18]), .I2(n20560[0]), 
            .I3(n50826), .O(n20511[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_952.LUT_INIT = 16'h8778;
    SB_LUT4 i35217_3_lut_4_lut (.I0(\Kp[2] ), .I1(n49[18]), .I2(n50826), 
            .I3(n20560[0]), .O(n4_adj_4679));   // verilog/motorControl.v(50[18:24])
    defparam i35217_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i35204_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n49[19]), .I2(n49[18]), 
            .I3(\Kp[1] ), .O(n20511[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35204_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_18_8 (.CI(n51230), .I0(n257[6]), .I1(n306[6]), .CO(n51231));
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n306[5]), .I3(n51229), 
            .O(n356[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_7 (.CI(n51229), .I0(n257[5]), .I1(n306[5]), .CO(n51230));
    SB_LUT4 i48900_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n65916));
    defparam i48900_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n306[4]), .I3(n51228), 
            .O(n356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35206_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n49[19]), .I2(n49[18]), 
            .I3(\Kp[1] ), .O(n50826));   // verilog/motorControl.v(50[18:24])
    defparam i35206_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4579));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4578));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n29183), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n29182), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n29181), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n29180), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n29179), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n29178), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n29177), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n29176), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n29175), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n29174), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n29173), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n29172), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n29171), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n29170), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n29169), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n29168), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n29164), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n29160), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n29159), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n29158), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n29157), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n29156), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n29155), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4577));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4576));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4575));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4574));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_6 (.CI(n51228), .I0(n257[4]), .I1(n306[4]), .CO(n51229));
    SB_LUT4 i1_3_lut_4_lut_adj_953 (.I0(\Kp[3] ), .I1(n49[19]), .I2(n20591[1]), 
            .I3(n4_adj_4681), .O(n20560[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_953.LUT_INIT = 16'h8778;
    SB_LUT4 i35444_3_lut_4_lut (.I0(\Kp[3] ), .I1(n49[19]), .I2(n4_adj_4681), 
            .I3(n20591[1]), .O(n6_adj_4603));   // verilog/motorControl.v(50[18:24])
    defparam i35444_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12_adj_4682));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n306[3]), .I3(n51227), 
            .O(n356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1936__i0 (.Q(counter[0]), .C(clk16MHz), .D(n51[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_CARRY add_18_5 (.CI(n51227), .I0(n257[3]), .I1(n306[3]), .CO(n51228));
    SB_LUT4 i4_3_lut (.I0(counter[5]), .I1(counter[2]), .I2(counter[0]), 
            .I3(GND_net), .O(n11_adj_4683));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut (.I0(counter[19]), .I1(counter[29]), .I2(counter[28]), 
            .I3(GND_net), .O(n8_adj_4684));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2609_4_lut (.I0(n11_adj_4683), .I1(counter[8]), .I2(counter[7]), 
            .I3(n12_adj_4682), .O(n18_adj_4685));
    defparam i2609_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_4686));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_4_lut (.I0(counter[24]), .I1(counter[30]), .I2(n8_adj_4684), 
            .I3(counter[27]), .O(n16_adj_4687));
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_954 (.I0(counter[23]), .I1(counter[12]), .I2(n10_adj_4686), 
            .I3(n18_adj_4685), .O(n15_adj_4688));
    defparam i1_4_lut_adj_954.LUT_INIT = 16'heaaa;
    SB_LUT4 i10_4_lut (.I0(counter[21]), .I1(counter[18]), .I2(counter[22]), 
            .I3(counter[26]), .O(n24_adj_4689));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(counter[17]), .I1(counter[20]), .I2(counter[16]), 
            .I3(counter[14]), .O(n23_adj_4690));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(counter[15]), .I1(n15_adj_4688), .I2(counter[25]), 
            .I3(n16_adj_4687), .O(n25_adj_4691));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23343_4_lut (.I0(n25_adj_4691), .I1(counter[31]), .I2(n23_adj_4690), 
            .I3(n24_adj_4689), .O(counter_31__N_3714));   // verilog/motorControl.v(26[8:41])
    defparam i23343_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i35436_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204_adj_4600), 
            .I3(n20591[0]), .O(n4_adj_4681));   // verilog/motorControl.v(50[18:24])
    defparam i35436_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_955 (.I0(n62), .I1(n131), .I2(n204_adj_4600), 
            .I3(n20591[0]), .O(n20560[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_955.LUT_INIT = 16'h8778;
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n306[2]), .I3(n51226), 
            .O(n356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_4 (.CI(n51226), .I0(n257[2]), .I1(n306[2]), .CO(n51227));
    SB_LUT4 i48934_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n65950));
    defparam i48934_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n306[1]), .I3(n51225), 
            .O(n356[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_3 (.CI(n51225), .I0(n257[1]), .I1(n306[1]), .CO(n51226));
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n306[0]), .I3(GND_net), 
            .O(n356[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n306[0]), .CO(n51225));
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n49[23]), .I3(n51224), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29023), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n49[22]), .I3(n51223), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[21]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[22]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[23]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .I1(n10731[21]), .I2(GND_net), .I3(n51983), .O(n10161[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4324_2_lut_4_lut (.I0(control_update), .I1(n68148), .I2(PWMLimit[23]), 
            .I3(n356[23]), .O(n9647));
    defparam i4324_2_lut_4_lut.LUT_INIT = 16'h2a02;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n356[7]), .I1(n436[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4693));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4694));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4695));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i45_2_lut (.I0(PWMLimit[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4696));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n10731[20]), .I2(GND_net), 
            .I3(n51982), .O(n306[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4697));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4698));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35288_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .O(n20536[0]));   // verilog/motorControl.v(50[27:38])
    defparam i35288_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4699));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4700));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4701));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4702));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n356[4]), .I1(n436[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4703));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n356[5]), .I1(n436[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4704));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n356[6]), .I1(n436[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4705));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4591));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4590));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4589));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4608));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4612));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4611));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4615));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4614));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4613));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4706));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4707));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4708));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4709));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4711));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4712));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4714));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4716));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4717));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4719));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4647));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4651));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4650));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4649));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4644));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4645));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4646));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4662));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4661));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4648));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4663));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_17_add_1225_23 (.CI(n51982), .I0(n10731[20]), .I1(GND_net), 
            .CO(n51983));
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4652));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n10731[19]), .I2(GND_net), 
            .I3(n51981), .O(n306[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_24 (.CI(n51223), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n49[22]), .CO(n51224));
    SB_CARRY mult_17_add_1225_22 (.CI(n51981), .I0(n10731[19]), .I1(GND_net), 
            .CO(n51982));
    SB_DFFER result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n1[23]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n49[21]), .I3(n51222), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n10731[18]), .I2(GND_net), 
            .I3(n51980), .O(n306[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_21 (.CI(n51980), .I0(n10731[18]), .I1(GND_net), 
            .CO(n51981));
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n10731[17]), .I2(GND_net), 
            .I3(n51979), .O(n306[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_20 (.CI(n51979), .I0(n10731[17]), .I1(GND_net), 
            .CO(n51980));
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n10731[16]), .I2(GND_net), 
            .I3(n51978), .O(n306[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n51978), .I0(n10731[16]), .I1(GND_net), 
            .CO(n51979));
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n10731[15]), .I2(GND_net), 
            .I3(n51977), .O(n306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n51977), .I0(n10731[15]), .I1(GND_net), 
            .CO(n51978));
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n10731[14]), .I2(GND_net), 
            .I3(n51976), .O(n306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n51222), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n49[21]), .CO(n51223));
    SB_CARRY mult_17_add_1225_17 (.CI(n51976), .I0(n10731[14]), .I1(GND_net), 
            .CO(n51977));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n10731[13]), .I2(n1096), 
            .I3(n51975), .O(n306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n51975), .I0(n10731[13]), .I1(n1096), 
            .CO(n51976));
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n10731[12]), .I2(n1023), 
            .I3(n51974), .O(n306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_15 (.CI(n51974), .I0(n10731[12]), .I1(n1023), 
            .CO(n51975));
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n49[20]), .I3(n51221), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_22 (.CI(n51221), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n49[20]), .CO(n51222));
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n49[19]), .I3(n51220), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n10731[11]), .I2(n950), 
            .I3(n51973), .O(n306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_14 (.CI(n51973), .I0(n10731[11]), .I1(n950), 
            .CO(n51974));
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n10731[10]), .I2(n877), 
            .I3(n51972), .O(n306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_13 (.CI(n51972), .I0(n10731[10]), .I1(n877), 
            .CO(n51973));
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n10731[9]), .I2(n804), 
            .I3(n51971), .O(n306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_21 (.CI(n51220), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n49[19]), .CO(n51221));
    SB_CARRY mult_17_add_1225_12 (.CI(n51971), .I0(n10731[9]), .I1(n804), 
            .CO(n51972));
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n10731[8]), .I2(n731), 
            .I3(n51970), .O(n306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_11 (.CI(n51970), .I0(n10731[8]), .I1(n731), 
            .CO(n51971));
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n10731[7]), .I2(n658), 
            .I3(n51969), .O(n306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n49[18]), .I3(n51219), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_10 (.CI(n51969), .I0(n10731[7]), .I1(n658), 
            .CO(n51970));
    SB_CARRY add_9_20 (.CI(n51219), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n49[18]), .CO(n51220));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n10731[6]), .I2(n585), 
            .I3(n51968), .O(n306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n49[17]), .I3(n51218), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_9 (.CI(n51968), .I0(n10731[6]), .I1(n585), 
            .CO(n51969));
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n10731[5]), .I2(n512), 
            .I3(n51967), .O(n306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n1[22]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY mult_17_add_1225_8 (.CI(n51967), .I0(n10731[5]), .I1(n512), 
            .CO(n51968));
    SB_DFFER result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n1[21]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n1[20]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n1[19]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n1[18]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n1[17]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n1[16]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n1[15]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n1[14]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n1[13]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n1[12]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n1[11]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n1[10]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n1[9]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n1[8]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n1[7]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n1[6]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n1[5]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n1[4]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n1[3]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n1[2]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n1[1]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_5134_10_lut (.I0(GND_net), .I1(n20136[7]), .I2(n700), 
            .I3(n51515), .O(n19956[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n51218), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n49[17]), .CO(n51219));
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n49[16]), .I3(n51217), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n10731[4]), .I2(n439_adj_4730), 
            .I3(n51966), .O(n306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i33_2_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4731));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5134_9_lut (.I0(GND_net), .I1(n20136[6]), .I2(n627), .I3(n51514), 
            .O(n19956[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5134_9 (.CI(n51514), .I0(n20136[6]), .I1(n627), .CO(n51515));
    SB_CARRY add_9_18 (.CI(n51217), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n49[16]), .CO(n51218));
    SB_CARRY mult_17_add_1225_7 (.CI(n51966), .I0(n10731[4]), .I1(n439_adj_4730), 
            .CO(n51967));
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n49[15]), .I3(n51216), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5134_8_lut (.I0(GND_net), .I1(n20136[5]), .I2(n554), .I3(n51513), 
            .O(n19956[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_17 (.CI(n51216), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n49[15]), .CO(n51217));
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n10731[3]), .I2(n366_adj_4733), 
            .I3(n51965), .O(n306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5134_8 (.CI(n51513), .I0(n20136[5]), .I1(n554), .CO(n51514));
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n49[14]), .I3(n51215), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_6 (.CI(n51965), .I0(n10731[3]), .I1(n366_adj_4733), 
            .CO(n51966));
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n10731[2]), .I2(n293_adj_4734), 
            .I3(n51964), .O(n306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5134_7_lut (.I0(GND_net), .I1(n20136[4]), .I2(n481), .I3(n51512), 
            .O(n19956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4735));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4736));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4737));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4738));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4739));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4740));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4741));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4742));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4743));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4744));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4745));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4746));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4747));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4748));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_5 (.CI(n51964), .I0(n10731[2]), .I1(n293_adj_4734), 
            .CO(n51965));
    SB_CARRY add_9_16 (.CI(n51215), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n49[14]), .CO(n51216));
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n49[13]), .I3(n51214), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5134_7 (.CI(n51512), .I0(n20136[4]), .I1(n481), .CO(n51513));
    SB_LUT4 add_5134_6_lut (.I0(GND_net), .I1(n20136[3]), .I2(n408), .I3(n51511), 
            .O(n19956[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5134_6 (.CI(n51511), .I0(n20136[3]), .I1(n408), .CO(n51512));
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n10731[1]), .I2(n220), 
            .I3(n51963), .O(n306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5134_5_lut (.I0(GND_net), .I1(n20136[2]), .I2(n335_adj_4749), 
            .I3(n51510), .O(n19956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5134_5 (.CI(n51510), .I0(n20136[2]), .I1(n335_adj_4749), 
            .CO(n51511));
    SB_LUT4 add_5134_4_lut (.I0(GND_net), .I1(n20136[1]), .I2(n262), .I3(n51509), 
            .O(n19956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5134_4 (.CI(n51509), .I0(n20136[1]), .I1(n262), .CO(n51510));
    SB_CARRY mult_17_add_1225_4 (.CI(n51963), .I0(n10731[1]), .I1(n220), 
            .CO(n51964));
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n10731[0]), .I2(n147_adj_4750), 
            .I3(n51962), .O(n306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5134_3_lut (.I0(GND_net), .I1(n20136[0]), .I2(n189_adj_4751), 
            .I3(n51508), .O(n19956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_3 (.CI(n51962), .I0(n10731[0]), .I1(n147_adj_4750), 
            .CO(n51963));
    SB_CARRY add_5134_3 (.CI(n51508), .I0(n20136[0]), .I1(n189_adj_4751), 
            .CO(n51509));
    SB_LUT4 add_5134_2_lut (.I0(GND_net), .I1(n47_adj_4752), .I2(n116), 
            .I3(GND_net), .O(n19956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5134_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5134_2 (.CI(GND_net), .I0(n47_adj_4752), .I1(n116), .CO(n51508));
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n49[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4753));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_15 (.CI(n51214), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n49[13]), .CO(n51215));
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n49[12]), .I3(n51213), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4755));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_14 (.CI(n51213), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n49[12]), .CO(n51214));
    SB_LUT4 LessThan_23_i27_2_lut (.I0(PWMLimit[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4756));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4757), .I2(n74), 
            .I3(GND_net), .O(n306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n49[11]), .I3(n51212), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_13 (.CI(n51212), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n49[11]), .CO(n51213));
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4758));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n49[10]), .I3(n51211), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5_adj_4757), .I1(n74), 
            .CO(n51962));
    SB_LUT4 LessThan_23_i29_2_lut (.I0(PWMLimit[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4759));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_23_lut (.I0(GND_net), .I1(n12441[20]), .I2(GND_net), 
            .I3(n51961), .O(n10731[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_22_lut (.I0(GND_net), .I1(n12441[19]), .I2(GND_net), 
            .I3(n51960), .O(n10731[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_12 (.CI(n51211), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n49[10]), .CO(n51212));
    SB_LUT4 LessThan_23_i31_2_lut (.I0(PWMLimit[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4760));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49214_4_lut (.I0(n21_adj_4736), .I1(n19_adj_4697), .I2(n17_adj_4698), 
            .I3(n9_adj_4699), .O(n66230));
    defparam i49214_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49197_4_lut (.I0(n27_adj_4756), .I1(n15_adj_4702), .I2(n13_adj_4701), 
            .I3(n11_adj_4700), .O(n66213));
    defparam i49197_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n49[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4762));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n49[9]), .I3(n51210), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33_adj_4731), 
            .I3(GND_net), .O(n12_adj_4764));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4765));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4766));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_11 (.CI(n51210), .I0(\PID_CONTROLLER.integral [9]), .I1(n49[9]), 
            .CO(n51211));
    SB_CARRY add_4426_22 (.CI(n51960), .I0(n12441[19]), .I1(GND_net), 
            .CO(n51961));
    SB_LUT4 add_4426_21_lut (.I0(GND_net), .I1(n12441[18]), .I2(GND_net), 
            .I3(n51959), .O(n10731[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_21 (.CI(n51959), .I0(n12441[18]), .I1(GND_net), 
            .CO(n51960));
    SB_LUT4 add_4426_20_lut (.I0(GND_net), .I1(n12441[17]), .I2(GND_net), 
            .I3(n51958), .O(n10731[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4767));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_20 (.CI(n51958), .I0(n12441[17]), .I1(GND_net), 
            .CO(n51959));
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_19_lut (.I0(GND_net), .I1(n12441[16]), .I2(GND_net), 
            .I3(n51957), .O(n10731[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n49[8]), .I3(n51209), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_4701), 
            .I3(GND_net), .O(n10_adj_4768));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_9_10 (.CI(n51209), .I0(\PID_CONTROLLER.integral [8]), .I1(n49[8]), 
            .CO(n51210));
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n49[7]), .I3(n51208), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_19 (.CI(n51957), .I0(n12441[16]), .I1(GND_net), 
            .CO(n51958));
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_18_lut (.I0(GND_net), .I1(n12441[15]), .I2(GND_net), 
            .I3(n51956), .O(n10731[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_9 (.CI(n51208), .I0(\PID_CONTROLLER.integral [7]), .I1(n49[7]), 
            .CO(n51209));
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n49[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4770));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n49[6]), .I3(n51207), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_8 (.CI(n51207), .I0(\PID_CONTROLLER.integral [6]), .I1(n49[6]), 
            .CO(n51208));
    SB_CARRY add_4426_18 (.CI(n51956), .I0(n12441[15]), .I1(GND_net), 
            .CO(n51957));
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4771));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4772));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4773));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i30_3_lut (.I0(n12_adj_4764), .I1(n363), .I2(n35), 
            .I3(GND_net), .O(n30_adj_4775));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4776));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4777));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_17_lut (.I0(GND_net), .I1(n12441[14]), .I2(GND_net), 
            .I3(n51955), .O(n10731[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50098_4_lut (.I0(n13_adj_4701), .I1(n11_adj_4700), .I2(n9_adj_4699), 
            .I3(n66259), .O(n67114));
    defparam i50098_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_17 (.CI(n51955), .I0(n12441[14]), .I1(GND_net), 
            .CO(n51956));
    SB_LUT4 add_4426_16_lut (.I0(GND_net), .I1(n12441[13]), .I2(n1099), 
            .I3(n51954), .O(n10731[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_1936__i1 (.Q(counter[1]), .C(clk16MHz), .D(n51[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i2 (.Q(counter[2]), .C(clk16MHz), .D(n51[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 i50084_4_lut (.I0(n19_adj_4697), .I1(n17_adj_4698), .I2(n15_adj_4702), 
            .I3(n67114), .O(n67100));
    defparam i50084_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_16 (.CI(n51954), .I0(n12441[13]), .I1(n1099), .CO(n51955));
    SB_LUT4 add_4426_15_lut (.I0(GND_net), .I1(n12441[12]), .I2(n1026), 
            .I3(n51953), .O(n10731[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_1936__i3 (.Q(counter[3]), .C(clk16MHz), .D(n51[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i4 (.Q(counter[4]), .C(clk16MHz), .D(n51[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i5 (.Q(counter[5]), .C(clk16MHz), .D(n51[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i6 (.Q(counter[6]), .C(clk16MHz), .D(n51[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i7 (.Q(counter[7]), .C(clk16MHz), .D(n51[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i8 (.Q(counter[8]), .C(clk16MHz), .D(n51[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i9 (.Q(counter[9]), .C(clk16MHz), .D(n51[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i10 (.Q(counter[10]), .C(clk16MHz), .D(n51[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i11 (.Q(counter[11]), .C(clk16MHz), .D(n51[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i12 (.Q(counter[12]), .C(clk16MHz), .D(n51[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i13 (.Q(counter[13]), .C(clk16MHz), .D(n51[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i14 (.Q(counter[14]), .C(clk16MHz), .D(n51[14]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i15 (.Q(counter[15]), .C(clk16MHz), .D(n51[15]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i16 (.Q(counter[16]), .C(clk16MHz), .D(n51[16]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i17 (.Q(counter[17]), .C(clk16MHz), .D(n51[17]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i18 (.Q(counter[18]), .C(clk16MHz), .D(n51[18]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i19 (.Q(counter[19]), .C(clk16MHz), .D(n51[19]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i20 (.Q(counter[20]), .C(clk16MHz), .D(n51[20]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i21 (.Q(counter[21]), .C(clk16MHz), .D(n51[21]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i22 (.Q(counter[22]), .C(clk16MHz), .D(n51[22]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i23 (.Q(counter[23]), .C(clk16MHz), .D(n51[23]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i24 (.Q(counter[24]), .C(clk16MHz), .D(n51[24]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i25 (.Q(counter[25]), .C(clk16MHz), .D(n51[25]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i26 (.Q(counter[26]), .C(clk16MHz), .D(n51[26]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i27 (.Q(counter[27]), .C(clk16MHz), .D(n51[27]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i28 (.Q(counter[28]), .C(clk16MHz), .D(n51[28]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i29 (.Q(counter[29]), .C(clk16MHz), .D(n51[29]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i30 (.Q(counter[30]), .C(clk16MHz), .D(n51[30]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1936__i31 (.Q(counter[31]), .C(clk16MHz), .D(n51[31]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_15 (.CI(n51953), .I0(n12441[12]), .I1(n1026), .CO(n51954));
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n49[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4778));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4779));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_14_lut (.I0(GND_net), .I1(n12441[11]), .I2(n953), 
            .I3(n51952), .O(n10731[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_14 (.CI(n51952), .I0(n12441[11]), .I1(n953), .CO(n51953));
    SB_LUT4 i51072_4_lut (.I0(n25_adj_4739), .I1(n23_adj_4737), .I2(n21_adj_4736), 
            .I3(n67100), .O(n68088));
    defparam i51072_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4780));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_13_lut (.I0(GND_net), .I1(n12441[10]), .I2(n880), 
            .I3(n51951), .O(n10731[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4781));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4782));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50503_4_lut (.I0(n31_adj_4760), .I1(n29_adj_4759), .I2(n27_adj_4756), 
            .I3(n68088), .O(n67519));
    defparam i50503_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4783));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_13 (.CI(n51951), .I0(n12441[10]), .I1(n880), .CO(n51952));
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51195_4_lut (.I0(n37_adj_4735), .I1(n35), .I2(n33_adj_4731), 
            .I3(n67519), .O(n68211));
    defparam i51195_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_12_lut (.I0(GND_net), .I1(n12441[9]), .I2(n807), 
            .I3(n51950), .O(n10731[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_12 (.CI(n51950), .I0(n12441[9]), .I1(n807), .CO(n51951));
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_11_lut (.I0(GND_net), .I1(n12441[8]), .I2(n734), 
            .I3(n51949), .O(n10731[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_11 (.CI(n51949), .I0(n12441[8]), .I1(n734), .CO(n51950));
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n49[5]), .I3(n51206), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4426_10_lut (.I0(GND_net), .I1(n12441[7]), .I2(n661), 
            .I3(n51948), .O(n10731[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_10 (.CI(n51948), .I0(n12441[7]), .I1(n661), .CO(n51949));
    SB_LUT4 add_4426_9_lut (.I0(GND_net), .I1(n12441[6]), .I2(n588), .I3(n51947), 
            .O(n10731[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_9 (.CI(n51947), .I0(n12441[6]), .I1(n588), .CO(n51948));
    SB_LUT4 add_4426_8_lut (.I0(GND_net), .I1(n12441[5]), .I2(n515), .I3(n51946), 
            .O(n10731[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_8 (.CI(n51946), .I0(n12441[5]), .I1(n515), .CO(n51947));
    SB_LUT4 add_4426_7_lut (.I0(GND_net), .I1(n12441[4]), .I2(n442_adj_4784), 
            .I3(n51945), .O(n10731[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_7 (.CI(n51945), .I0(n12441[4]), .I1(n442_adj_4784), 
            .CO(n51946));
    SB_LUT4 add_4426_6_lut (.I0(GND_net), .I1(n12441[3]), .I2(n369_adj_4785), 
            .I3(n51944), .O(n10731[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_6 (.CI(n51944), .I0(n12441[3]), .I1(n369_adj_4785), 
            .CO(n51945));
    SB_LUT4 add_4426_5_lut (.I0(GND_net), .I1(n12441[2]), .I2(n296_adj_4786), 
            .I3(n51943), .O(n10731[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4426_5 (.CI(n51943), .I0(n12441[2]), .I1(n296_adj_4786), 
            .CO(n51944));
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n49[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4787));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4788));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_4_lut (.I0(GND_net), .I1(n12441[1]), .I2(n223), .I3(n51942), 
            .O(n10731[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4789));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_4 (.CI(n51942), .I0(n12441[1]), .I1(n223), .CO(n51943));
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4790));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4426_3_lut (.I0(GND_net), .I1(n12441[0]), .I2(n150_adj_4791), 
            .I3(n51941), .O(n10731[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4792));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4793));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_3 (.CI(n51941), .I0(n12441[0]), .I1(n150_adj_4791), 
            .CO(n51942));
    SB_LUT4 add_4426_2_lut (.I0(GND_net), .I1(n8_adj_4794), .I2(n77_adj_4795), 
            .I3(GND_net), .O(n10731[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4426_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4796));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4426_2 (.CI(GND_net), .I0(n8_adj_4794), .I1(n77_adj_4795), 
            .CO(n51941));
    SB_LUT4 add_4721_22_lut (.I0(GND_net), .I1(n13743[19]), .I2(GND_net), 
            .I3(n51940), .O(n12441[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4797));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4798));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_21_lut (.I0(GND_net), .I1(n13743[18]), .I2(GND_net), 
            .I3(n51939), .O(n12441[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_21 (.CI(n51939), .I0(n13743[18]), .I1(GND_net), 
            .CO(n51940));
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4799));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4800));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4801));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4802));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_20_lut (.I0(GND_net), .I1(n13743[17]), .I2(GND_net), 
            .I3(n51938), .O(n12441[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_20 (.CI(n51938), .I0(n13743[17]), .I1(GND_net), 
            .CO(n51939));
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4803));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4804));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4805));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n49[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4806));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4807));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_19_lut (.I0(GND_net), .I1(n13743[16]), .I2(GND_net), 
            .I3(n51937), .O(n12441[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_19 (.CI(n51937), .I0(n13743[16]), .I1(GND_net), 
            .CO(n51938));
    SB_LUT4 add_4721_18_lut (.I0(GND_net), .I1(n13743[15]), .I2(GND_net), 
            .I3(n51936), .O(n12441[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_18 (.CI(n51936), .I0(n13743[15]), .I1(GND_net), 
            .CO(n51937));
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4808));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_17_lut (.I0(GND_net), .I1(n13743[14]), .I2(GND_net), 
            .I3(n51935), .O(n12441[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_17 (.CI(n51935), .I0(n13743[14]), .I1(GND_net), 
            .CO(n51936));
    SB_CARRY add_9_7 (.CI(n51206), .I0(\PID_CONTROLLER.integral [5]), .I1(n49[5]), 
            .CO(n51207));
    SB_LUT4 add_4721_16_lut (.I0(GND_net), .I1(n13743[13]), .I2(n1102_adj_4809), 
            .I3(n51934), .O(n12441[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4810));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4721_16 (.CI(n51934), .I0(n13743[13]), .I1(n1102_adj_4809), 
            .CO(n51935));
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4752));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_15_lut (.I0(GND_net), .I1(n13743[12]), .I2(n1029_adj_4811), 
            .I3(n51933), .O(n12441[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4812));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4721_15 (.CI(n51933), .I0(n13743[12]), .I1(n1029_adj_4811), 
            .CO(n51934));
    SB_LUT4 add_4721_14_lut (.I0(GND_net), .I1(n13743[11]), .I2(n956_adj_4813), 
            .I3(n51932), .O(n12441[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_14 (.CI(n51932), .I0(n13743[11]), .I1(n956_adj_4813), 
            .CO(n51933));
    SB_LUT4 add_4721_13_lut (.I0(GND_net), .I1(n13743[10]), .I2(n883_adj_4814), 
            .I3(n51931), .O(n12441[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_13 (.CI(n51931), .I0(n13743[10]), .I1(n883_adj_4814), 
            .CO(n51932));
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4815));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_12_lut (.I0(GND_net), .I1(n13743[9]), .I2(n810_adj_4816), 
            .I3(n51930), .O(n12441[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_12 (.CI(n51930), .I0(n13743[9]), .I1(n810_adj_4816), 
            .CO(n51931));
    SB_LUT4 add_4721_11_lut (.I0(GND_net), .I1(n13743[8]), .I2(n737_adj_4817), 
            .I3(n51929), .O(n12441[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4818));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4819));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n49[4]), .I3(n51205), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_4742), 
            .I3(GND_net), .O(n16_adj_4820));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4721_11 (.CI(n51929), .I0(n13743[8]), .I1(n737_adj_4817), 
            .CO(n51930));
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4821));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4822));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_10_lut (.I0(GND_net), .I1(n13743[7]), .I2(n664_adj_4823), 
            .I3(n51928), .O(n12441[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_10 (.CI(n51928), .I0(n13743[7]), .I1(n664_adj_4823), 
            .CO(n51929));
    SB_LUT4 add_4721_9_lut (.I0(GND_net), .I1(n13743[6]), .I2(n591_adj_4824), 
            .I3(n51927), .O(n12441[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_9 (.CI(n51927), .I0(n13743[6]), .I1(n591_adj_4824), 
            .CO(n51928));
    SB_LUT4 add_4721_8_lut (.I0(GND_net), .I1(n13743[5]), .I2(n518_adj_4825), 
            .I3(n51926), .O(n12441[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4826));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4827));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4828));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4829));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4830));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4831));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4832));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4833));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4834));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4721_8 (.CI(n51926), .I0(n13743[5]), .I1(n518_adj_4825), 
            .CO(n51927));
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4835));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4836));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4837));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4838));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4839));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4721_7_lut (.I0(GND_net), .I1(n13743[4]), .I2(n445_adj_4840), 
            .I3(n51925), .O(n12441[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4841));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4842));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4843));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50825_3_lut (.I0(n6_adj_4844), .I1(n356[10]), .I2(n21_adj_4736), 
            .I3(GND_net), .O(n67841));   // verilog/motorControl.v(52[14:29])
    defparam i50825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4845));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4721_7 (.CI(n51925), .I0(n13743[4]), .I1(n445_adj_4840), 
            .CO(n51926));
    SB_LUT4 add_4721_6_lut (.I0(GND_net), .I1(n13743[3]), .I2(n372_adj_4846), 
            .I3(n51924), .O(n12441[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_6 (.CI(n51924), .I0(n13743[3]), .I1(n372_adj_4846), 
            .CO(n51925));
    SB_LUT4 add_4721_5_lut (.I0(GND_net), .I1(n13743[2]), .I2(n299_adj_4847), 
            .I3(n51923), .O(n12441[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_6 (.CI(n51205), .I0(\PID_CONTROLLER.integral [4]), .I1(n49[4]), 
            .CO(n51206));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n49[3]), .I3(n51204), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_5 (.CI(n51923), .I0(n13743[2]), .I1(n299_adj_4847), 
            .CO(n51924));
    SB_LUT4 add_4721_4_lut (.I0(GND_net), .I1(n13743[1]), .I2(n226_adj_4848), 
            .I3(n51922), .O(n12441[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_4 (.CI(n51922), .I0(n13743[1]), .I1(n226_adj_4848), 
            .CO(n51923));
    SB_LUT4 add_4721_3_lut (.I0(GND_net), .I1(n13743[0]), .I2(n153_adj_4849), 
            .I3(n51921), .O(n12441[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_3 (.CI(n51921), .I0(n13743[0]), .I1(n153_adj_4849), 
            .CO(n51922));
    SB_LUT4 add_4721_2_lut (.I0(GND_net), .I1(n11_adj_4850), .I2(n80_adj_4851), 
            .I3(GND_net), .O(n12441[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4721_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4721_2 (.CI(GND_net), .I0(n11_adj_4850), .I1(n80_adj_4851), 
            .CO(n51921));
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4852));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4853));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4854));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4779_21_lut (.I0(GND_net), .I1(n14896[18]), .I2(GND_net), 
            .I3(n51920), .O(n13743[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_20_lut (.I0(GND_net), .I1(n14896[17]), .I2(GND_net), 
            .I3(n51919), .O(n13743[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_5 (.CI(n51204), .I0(\PID_CONTROLLER.integral [3]), .I1(n49[3]), 
            .CO(n51205));
    SB_CARRY add_4779_20 (.CI(n51919), .I0(n14896[17]), .I1(GND_net), 
            .CO(n51920));
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4855));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4856));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4857));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50826_3_lut (.I0(n67841), .I1(n356[11]), .I2(n23_adj_4737), 
            .I3(GND_net), .O(n67842));   // verilog/motorControl.v(52[14:29])
    defparam i50826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4858));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4859));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4860));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n49[2]), .I3(n51203), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_4 (.CI(n51203), .I0(\PID_CONTROLLER.integral [2]), .I1(n49[2]), 
            .CO(n51204));
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4861));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n49[1]), .I3(n51202), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4779_19_lut (.I0(GND_net), .I1(n14896[16]), .I2(GND_net), 
            .I3(n51918), .O(n13743[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4862));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4779_19 (.CI(n51918), .I0(n14896[16]), .I1(GND_net), 
            .CO(n51919));
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4863));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4864));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4779_18_lut (.I0(GND_net), .I1(n14896[15]), .I2(GND_net), 
            .I3(n51917), .O(n13743[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_18 (.CI(n51917), .I0(n14896[15]), .I1(GND_net), 
            .CO(n51918));
    SB_LUT4 add_4779_17_lut (.I0(GND_net), .I1(n14896[14]), .I2(GND_net), 
            .I3(n51916), .O(n13743[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_17 (.CI(n51916), .I0(n14896[14]), .I1(GND_net), 
            .CO(n51917));
    SB_LUT4 add_4779_16_lut (.I0(GND_net), .I1(n14896[13]), .I2(n1105_adj_4865), 
            .I3(n51915), .O(n13743[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_3 (.CI(n51202), .I0(\PID_CONTROLLER.integral [1]), .I1(n49[1]), 
            .CO(n51203));
    SB_CARRY add_4779_16 (.CI(n51915), .I0(n14896[13]), .I1(n1105_adj_4865), 
            .CO(n51916));
    SB_LUT4 add_4779_15_lut (.I0(GND_net), .I1(n14896[12]), .I2(n1032_adj_4866), 
            .I3(n51914), .O(n13743[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4867));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4868));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n49[0]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n49[0]), 
            .CO(n51202));
    SB_CARRY add_4779_15 (.CI(n51914), .I0(n14896[12]), .I1(n1032_adj_4866), 
            .CO(n51915));
    SB_LUT4 add_4779_14_lut (.I0(GND_net), .I1(n14896[11]), .I2(n959_adj_4869), 
            .I3(n51913), .O(n13743[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_14 (.CI(n51913), .I0(n14896[11]), .I1(n959_adj_4869), 
            .CO(n51914));
    SB_LUT4 add_4779_13_lut (.I0(GND_net), .I1(n14896[10]), .I2(n886_adj_4870), 
            .I3(n51912), .O(n13743[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_13 (.CI(n51912), .I0(n14896[10]), .I1(n886_adj_4870), 
            .CO(n51913));
    SB_LUT4 add_4779_12_lut (.I0(GND_net), .I1(n14896[9]), .I2(n813_adj_4871), 
            .I3(n51911), .O(n13743[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4872));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4873));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4874));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n51201), .O(n49[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_4698), 
            .I3(GND_net), .O(n8_adj_4875));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4876));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n51200), .O(n49[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_24 (.CI(n51200), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n51201));
    SB_CARRY add_4779_12 (.CI(n51911), .I0(n14896[9]), .I1(n813_adj_4871), 
            .CO(n51912));
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4779_11_lut (.I0(GND_net), .I1(n14896[8]), .I2(n740_adj_4878), 
            .I3(n51910), .O(n13743[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_11 (.CI(n51910), .I0(n14896[8]), .I1(n740_adj_4878), 
            .CO(n51911));
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4879));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4779_10_lut (.I0(GND_net), .I1(n14896[7]), .I2(n667_adj_4880), 
            .I3(n51909), .O(n13743[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4881));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4779_10 (.CI(n51909), .I0(n14896[7]), .I1(n667_adj_4880), 
            .CO(n51910));
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4882));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4883));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4884));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4885));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4779_9_lut (.I0(GND_net), .I1(n14896[6]), .I2(n594_adj_4886), 
            .I3(n51908), .O(n13743[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_9 (.CI(n51908), .I0(n14896[6]), .I1(n594_adj_4886), 
            .CO(n51909));
    SB_LUT4 add_4779_8_lut (.I0(GND_net), .I1(n14896[5]), .I2(n521_adj_4887), 
            .I3(n51907), .O(n13743[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_8 (.CI(n51907), .I0(n14896[5]), .I1(n521_adj_4887), 
            .CO(n51908));
    SB_LUT4 add_4779_7_lut (.I0(GND_net), .I1(n14896[4]), .I2(n448_adj_4888), 
            .I3(n51906), .O(n13743[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_7 (.CI(n51906), .I0(n14896[4]), .I1(n448_adj_4888), 
            .CO(n51907));
    SB_LUT4 add_4779_6_lut (.I0(GND_net), .I1(n14896[3]), .I2(n375_adj_4889), 
            .I3(n51905), .O(n13743[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_6 (.CI(n51905), .I0(n14896[3]), .I1(n375_adj_4889), 
            .CO(n51906));
    SB_LUT4 add_4779_5_lut (.I0(GND_net), .I1(n14896[2]), .I2(n302_adj_4890), 
            .I3(n51904), .O(n13743[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_5 (.CI(n51904), .I0(n14896[2]), .I1(n302_adj_4890), 
            .CO(n51905));
    SB_LUT4 add_4779_4_lut (.I0(GND_net), .I1(n14896[1]), .I2(n229_adj_4891), 
            .I3(n51903), .O(n13743[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_4 (.CI(n51903), .I0(n14896[1]), .I1(n229_adj_4891), 
            .CO(n51904));
    SB_LUT4 add_4779_3_lut (.I0(GND_net), .I1(n14896[0]), .I2(n156_adj_4892), 
            .I3(n51902), .O(n13743[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_3 (.CI(n51902), .I0(n14896[0]), .I1(n156_adj_4892), 
            .CO(n51903));
    SB_LUT4 add_4779_2_lut (.I0(GND_net), .I1(n14_adj_4893), .I2(n83_adj_4894), 
            .I3(GND_net), .O(n13743[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4779_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4779_2 (.CI(GND_net), .I0(n14_adj_4893), .I1(n83_adj_4894), 
            .CO(n51902));
    SB_LUT4 add_5125_11_lut (.I0(GND_net), .I1(n20055[8]), .I2(n770_adj_4895), 
            .I3(n51901), .O(n19856[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5125_10_lut (.I0(GND_net), .I1(n20055[7]), .I2(n697_adj_4896), 
            .I3(n51900), .O(n19856[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_10 (.CI(n51900), .I0(n20055[7]), .I1(n697_adj_4896), 
            .CO(n51901));
    SB_LUT4 add_5125_9_lut (.I0(GND_net), .I1(n20055[6]), .I2(n624_adj_4897), 
            .I3(n51899), .O(n19856[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_9 (.CI(n51899), .I0(n20055[6]), .I1(n624_adj_4897), 
            .CO(n51900));
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n51199), .O(n49[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_23 (.CI(n51199), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n51200));
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n51198), .O(n49[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_22 (.CI(n51198), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n51199));
    SB_LUT4 add_5125_8_lut (.I0(GND_net), .I1(n20055[5]), .I2(n551_adj_4898), 
            .I3(n51898), .O(n19856[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_8 (.CI(n51898), .I0(n20055[5]), .I1(n551_adj_4898), 
            .CO(n51899));
    SB_LUT4 add_5125_7_lut (.I0(GND_net), .I1(n20055[4]), .I2(n478_adj_4899), 
            .I3(n51897), .O(n19856[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_7 (.CI(n51897), .I0(n20055[4]), .I1(n478_adj_4899), 
            .CO(n51898));
    SB_LUT4 add_5125_6_lut (.I0(GND_net), .I1(n20055[3]), .I2(n405_adj_4900), 
            .I3(n51896), .O(n19856[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_6 (.CI(n51896), .I0(n20055[3]), .I1(n405_adj_4900), 
            .CO(n51897));
    SB_LUT4 add_5125_5_lut (.I0(GND_net), .I1(n20055[2]), .I2(n332_adj_4901), 
            .I3(n51895), .O(n19856[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_5 (.CI(n51895), .I0(n20055[2]), .I1(n332_adj_4901), 
            .CO(n51896));
    SB_LUT4 add_5125_4_lut (.I0(GND_net), .I1(n20055[1]), .I2(n259_adj_4902), 
            .I3(n51894), .O(n19856[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_4 (.CI(n51894), .I0(n20055[1]), .I1(n259_adj_4902), 
            .CO(n51895));
    SB_LUT4 add_5125_3_lut (.I0(GND_net), .I1(n20055[0]), .I2(n186_adj_4903), 
            .I3(n51893), .O(n19856[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_3 (.CI(n51893), .I0(n20055[0]), .I1(n186_adj_4903), 
            .CO(n51894));
    SB_LUT4 add_5125_2_lut (.I0(GND_net), .I1(n44_adj_4904), .I2(n113_adj_4905), 
            .I3(GND_net), .O(n19856[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5125_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5125_2 (.CI(GND_net), .I0(n44_adj_4904), .I1(n113_adj_4905), 
            .CO(n51893));
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n51197), .O(n49[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_21 (.CI(n51197), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n51198));
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(n14), 
            .I3(n51196), .O(n49[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_20 (.CI(n51196), .I0(setpoint[18]), .I1(n14), 
            .CO(n51197));
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n51195), .O(n49[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_19 (.CI(n51195), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n51196));
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n51194), .O(n49[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51380_4_lut (.I0(\encoder1_position_scaled[0] ), .I1(n15), 
            .I2(n65364), .I3(n15_adj_1), .O(motor_state[0]));   // verilog/motorControl.v(43[15:31])
    defparam i51380_4_lut.LUT_INIT = 16'h3f77;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4909));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_18 (.CI(n51194), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n51195));
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4910));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4911));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n51193), .O(n49[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_17 (.CI(n51193), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n51194));
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n51192), .O(n49[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_16 (.CI(n51192), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n51193));
    SB_LUT4 i51498_4_lut (.I0(\encoder1_position_scaled[1] ), .I1(n15), 
            .I2(n65475), .I3(n15_adj_1), .O(motor_state[1]));   // verilog/motorControl.v(43[15:31])
    defparam i51498_4_lut.LUT_INIT = 16'h3f77;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4912));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4913));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n51191), .O(n49[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51495_4_lut (.I0(\encoder1_position_scaled[2] ), .I1(n15), 
            .I2(n65474), .I3(n15_adj_1), .O(motor_state[2]));   // verilog/motorControl.v(43[15:31])
    defparam i51495_4_lut.LUT_INIT = 16'h3f77;
    SB_CARRY sub_8_add_2_15 (.CI(n51191), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n51192));
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4914));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n51190), .O(n49[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_14 (.CI(n51190), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n51191));
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n51189), .O(n49[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4915));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4916));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4917));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i24_3_lut (.I0(n16_adj_4820), .I1(n356[22]), .I2(n45_adj_4696), 
            .I3(GND_net), .O(n24_adj_4918));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4919));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4920));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49167_4_lut (.I0(n43_adj_4742), .I1(n25_adj_4739), .I2(n23_adj_4737), 
            .I3(n66230), .O(n66183));
    defparam i49167_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50650_4_lut (.I0(n24_adj_4918), .I1(n8_adj_4875), .I2(n45_adj_4696), 
            .I3(n66177), .O(n67666));   // verilog/motorControl.v(52[14:29])
    defparam i50650_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4921));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4922));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4923));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49640_3_lut (.I0(n67842), .I1(n356[12]), .I2(n25_adj_4739), 
            .I3(GND_net), .O(n66656));   // verilog/motorControl.v(52[14:29])
    defparam i49640_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_8_add_2_13 (.CI(n51189), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n51190));
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n51188), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_12 (.CI(n51188), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n51189));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(n38106), 
            .I3(n51187), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_11 (.CI(n51187), .I0(setpoint[9]), .I1(n38106), 
            .CO(n51188));
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4924));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4925));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n51186), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i4_4_lut (.I0(PWMLimit[0]), .I1(n356[1]), .I2(PWMLimit[1]), 
            .I3(n356[0]), .O(n4_adj_4926));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY sub_8_add_2_10 (.CI(n51186), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n51187));
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n51185), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50823_3_lut (.I0(n4_adj_4926), .I1(n356[13]), .I2(n27_adj_4756), 
            .I3(GND_net), .O(n67839));   // verilog/motorControl.v(52[14:29])
    defparam i50823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50824_3_lut (.I0(n67839), .I1(n356[14]), .I2(n29_adj_4759), 
            .I3(GND_net), .O(n67840));   // verilog/motorControl.v(52[14:29])
    defparam i50824_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_8_add_2_9 (.CI(n51185), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n51186));
    SB_LUT4 add_4831_20_lut (.I0(GND_net), .I1(n15911[17]), .I2(GND_net), 
            .I3(n51869), .O(n14896[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4831_19_lut (.I0(GND_net), .I1(n15911[16]), .I2(GND_net), 
            .I3(n51868), .O(n14896[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_19 (.CI(n51868), .I0(n15911[16]), .I1(GND_net), 
            .CO(n51869));
    SB_LUT4 add_4831_18_lut (.I0(GND_net), .I1(n15911[15]), .I2(GND_net), 
            .I3(n51867), .O(n14896[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n51184), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_18 (.CI(n51867), .I0(n15911[15]), .I1(GND_net), 
            .CO(n51868));
    SB_CARRY sub_8_add_2_8 (.CI(n51184), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n51185));
    SB_LUT4 add_4831_17_lut (.I0(GND_net), .I1(n15911[14]), .I2(GND_net), 
            .I3(n51866), .O(n14896[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_17 (.CI(n51866), .I0(n15911[14]), .I1(GND_net), 
            .CO(n51867));
    SB_LUT4 add_4831_16_lut (.I0(GND_net), .I1(n15911[13]), .I2(n1108_adj_4925), 
            .I3(n51865), .O(n14896[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n51183), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n51183), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n51184));
    SB_CARRY add_4831_16 (.CI(n51865), .I0(n15911[13]), .I1(n1108_adj_4925), 
            .CO(n51866));
    SB_LUT4 add_4831_15_lut (.I0(GND_net), .I1(n15911[12]), .I2(n1035_adj_4924), 
            .I3(n51864), .O(n14896[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n51182), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49191_4_lut (.I0(n33_adj_4731), .I1(n31_adj_4760), .I2(n29_adj_4759), 
            .I3(n66213), .O(n66207));
    defparam i49191_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4831_15 (.CI(n51864), .I0(n15911[12]), .I1(n1035_adj_4924), 
            .CO(n51865));
    SB_LUT4 add_4831_14_lut (.I0(GND_net), .I1(n15911[11]), .I2(n962_adj_4923), 
            .I3(n51863), .O(n14896[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_14 (.CI(n51863), .I0(n15911[11]), .I1(n962_adj_4923), 
            .CO(n51864));
    SB_LUT4 add_4831_13_lut (.I0(GND_net), .I1(n15911[10]), .I2(n889_adj_4922), 
            .I3(n51862), .O(n14896[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_13 (.CI(n51862), .I0(n15911[10]), .I1(n889_adj_4922), 
            .CO(n51863));
    SB_LUT4 add_4831_12_lut (.I0(GND_net), .I1(n15911[9]), .I2(n816_adj_4921), 
            .I3(n51861), .O(n14896[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_6 (.CI(n51182), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n51183));
    SB_LUT4 sub_8_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(\motor_state[3] ), 
            .I3(n51181), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_12 (.CI(n51861), .I0(n15911[9]), .I1(n816_adj_4921), 
            .CO(n51862));
    SB_LUT4 add_4831_11_lut (.I0(GND_net), .I1(n15911[8]), .I2(n743_adj_4920), 
            .I3(n51860), .O(n14896[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_11 (.CI(n51860), .I0(n15911[8]), .I1(n743_adj_4920), 
            .CO(n51861));
    SB_LUT4 add_4831_10_lut (.I0(GND_net), .I1(n15911[7]), .I2(n670_adj_4919), 
            .I3(n51859), .O(n14896[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_10 (.CI(n51859), .I0(n15911[7]), .I1(n670_adj_4919), 
            .CO(n51860));
    SB_LUT4 add_4831_9_lut (.I0(GND_net), .I1(n15911[6]), .I2(n597_adj_4917), 
            .I3(n51858), .O(n14896[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_9 (.CI(n51858), .I0(n15911[6]), .I1(n597_adj_4917), 
            .CO(n51859));
    SB_LUT4 add_4831_8_lut (.I0(GND_net), .I1(n15911[5]), .I2(n524_adj_4916), 
            .I3(n51857), .O(n14896[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_5 (.CI(n51181), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n51182));
    SB_CARRY add_4831_8 (.CI(n51857), .I0(n15911[5]), .I1(n524_adj_4916), 
            .CO(n51858));
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4905));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n49[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4904));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4903));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4831_7_lut (.I0(GND_net), .I1(n15911[4]), .I2(n451_adj_4915), 
            .I3(n51856), .O(n14896[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4902));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4831_7 (.CI(n51856), .I0(n15911[4]), .I1(n451_adj_4915), 
            .CO(n51857));
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4901));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4831_6_lut (.I0(GND_net), .I1(n15911[3]), .I2(n378_adj_4914), 
            .I3(n51855), .O(n14896[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4900));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4899));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4898));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4831_6 (.CI(n51855), .I0(n15911[3]), .I1(n378_adj_4914), 
            .CO(n51856));
    SB_LUT4 sub_8_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n51180), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4831_5_lut (.I0(GND_net), .I1(n15911[2]), .I2(n305_adj_4913), 
            .I3(n51854), .O(n14896[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_4 (.CI(n51180), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n51181));
    SB_CARRY add_4831_5 (.CI(n51854), .I0(n15911[2]), .I1(n305_adj_4913), 
            .CO(n51855));
    SB_LUT4 add_4831_4_lut (.I0(GND_net), .I1(n15911[1]), .I2(n232_adj_4912), 
            .I3(n51853), .O(n14896[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n51179), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_4 (.CI(n51853), .I0(n15911[1]), .I1(n232_adj_4912), 
            .CO(n51854));
    SB_LUT4 add_4831_3_lut (.I0(GND_net), .I1(n15911[0]), .I2(n159_adj_4911), 
            .I3(n51852), .O(n14896[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_3 (.CI(n51852), .I0(n15911[0]), .I1(n159_adj_4911), 
            .CO(n51853));
    SB_LUT4 add_4831_2_lut (.I0(GND_net), .I1(n17_adj_4910), .I2(n86_adj_4909), 
            .I3(GND_net), .O(n14896[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4831_2 (.CI(GND_net), .I0(n17_adj_4910), .I1(n86_adj_4909), 
            .CO(n51852));
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4897));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4896));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_3 (.CI(n51179), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n51180));
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4895));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4894));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4893));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51159_4_lut (.I0(n30_adj_4775), .I1(n10_adj_4768), .I2(n35), 
            .I3(n66205), .O(n68175));   // verilog/motorControl.v(52[14:29])
    defparam i51159_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4892));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4891));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49642_3_lut (.I0(n67840), .I1(n356[15]), .I2(n31_adj_4760), 
            .I3(GND_net), .O(n66658));   // verilog/motorControl.v(52[14:29])
    defparam i49642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4890));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4889));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4888));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4887));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n51179));
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4886));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4880));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4878));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51294_4_lut (.I0(n66658), .I1(n68175), .I2(n35), .I3(n66207), 
            .O(n68310));   // verilog/motorControl.v(52[14:29])
    defparam i51294_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4879_19_lut (.I0(GND_net), .I1(n16722[16]), .I2(GND_net), 
            .I3(n51810), .O(n15911[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4879_18_lut (.I0(GND_net), .I1(n16722[15]), .I2(GND_net), 
            .I3(n51809), .O(n15911[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_18 (.CI(n51809), .I0(n16722[15]), .I1(GND_net), 
            .CO(n51810));
    SB_LUT4 add_4879_17_lut (.I0(GND_net), .I1(n16722[14]), .I2(GND_net), 
            .I3(n51808), .O(n15911[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_17 (.CI(n51808), .I0(n16722[14]), .I1(GND_net), 
            .CO(n51809));
    SB_LUT4 add_4879_16_lut (.I0(GND_net), .I1(n16722[13]), .I2(n1111_adj_4885), 
            .I3(n51807), .O(n15911[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_16 (.CI(n51807), .I0(n16722[13]), .I1(n1111_adj_4885), 
            .CO(n51808));
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4871));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4870));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4869));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4879_15_lut (.I0(GND_net), .I1(n16722[12]), .I2(n1038_adj_4884), 
            .I3(n51806), .O(n15911[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_15 (.CI(n51806), .I0(n16722[12]), .I1(n1038_adj_4884), 
            .CO(n51807));
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4866));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4879_14_lut (.I0(GND_net), .I1(n16722[11]), .I2(n965_adj_4883), 
            .I3(n51805), .O(n15911[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_14 (.CI(n51805), .I0(n16722[11]), .I1(n965_adj_4883), 
            .CO(n51806));
    SB_LUT4 add_4879_13_lut (.I0(GND_net), .I1(n16722[10]), .I2(n892_adj_4882), 
            .I3(n51804), .O(n15911[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_13 (.CI(n51804), .I0(n16722[10]), .I1(n892_adj_4882), 
            .CO(n51805));
    SB_LUT4 add_4879_12_lut (.I0(GND_net), .I1(n16722[9]), .I2(n819_adj_4881), 
            .I3(n51803), .O(n15911[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_12 (.CI(n51803), .I0(n16722[9]), .I1(n819_adj_4881), 
            .CO(n51804));
    SB_LUT4 add_4879_11_lut (.I0(GND_net), .I1(n16722[8]), .I2(n746_adj_4879), 
            .I3(n51802), .O(n15911[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_11 (.CI(n51802), .I0(n16722[8]), .I1(n746_adj_4879), 
            .CO(n51803));
    SB_LUT4 add_4879_10_lut (.I0(GND_net), .I1(n16722[7]), .I2(n673_adj_4877), 
            .I3(n51801), .O(n15911[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_10 (.CI(n51801), .I0(n16722[7]), .I1(n673_adj_4877), 
            .CO(n51802));
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4865));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4879_9_lut (.I0(GND_net), .I1(n16722[6]), .I2(n600_adj_4876), 
            .I3(n51800), .O(n15911[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_9 (.CI(n51800), .I0(n16722[6]), .I1(n600_adj_4876), 
            .CO(n51801));
    SB_LUT4 add_4879_8_lut (.I0(GND_net), .I1(n16722[5]), .I2(n527_adj_4874), 
            .I3(n51799), .O(n15911[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_8 (.CI(n51799), .I0(n16722[5]), .I1(n527_adj_4874), 
            .CO(n51800));
    SB_LUT4 add_4879_7_lut (.I0(GND_net), .I1(n16722[4]), .I2(n454_adj_4873), 
            .I3(n51798), .O(n15911[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_7 (.CI(n51798), .I0(n16722[4]), .I1(n454_adj_4873), 
            .CO(n51799));
    SB_LUT4 add_4879_6_lut (.I0(GND_net), .I1(n16722[3]), .I2(n381_adj_4872), 
            .I3(n51797), .O(n15911[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_6 (.CI(n51797), .I0(n16722[3]), .I1(n381_adj_4872), 
            .CO(n51798));
    SB_LUT4 add_4879_5_lut (.I0(GND_net), .I1(n16722[2]), .I2(n308_adj_4868), 
            .I3(n51796), .O(n15911[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_5 (.CI(n51796), .I0(n16722[2]), .I1(n308_adj_4868), 
            .CO(n51797));
    SB_LUT4 add_4879_4_lut (.I0(GND_net), .I1(n16722[1]), .I2(n235_adj_4867), 
            .I3(n51795), .O(n15911[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_4 (.CI(n51795), .I0(n16722[1]), .I1(n235_adj_4867), 
            .CO(n51796));
    SB_LUT4 add_4879_3_lut (.I0(GND_net), .I1(n16722[0]), .I2(n162_adj_4864), 
            .I3(n51794), .O(n15911[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_3 (.CI(n51794), .I0(n16722[0]), .I1(n162_adj_4864), 
            .CO(n51795));
    SB_LUT4 add_4879_2_lut (.I0(GND_net), .I1(n20_adj_4863), .I2(n89_adj_4862), 
            .I3(GND_net), .O(n15911[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4879_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4879_2 (.CI(GND_net), .I0(n20_adj_4863), .I1(n89_adj_4862), 
            .CO(n51794));
    SB_LUT4 add_5143_10_lut (.I0(GND_net), .I1(n20216[7]), .I2(n700_adj_4861), 
            .I3(n51793), .O(n20055[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5143_9_lut (.I0(GND_net), .I1(n20216[6]), .I2(n627_adj_4860), 
            .I3(n51792), .O(n20055[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5143_9 (.CI(n51792), .I0(n20216[6]), .I1(n627_adj_4860), 
            .CO(n51793));
    SB_LUT4 add_5143_8_lut (.I0(GND_net), .I1(n20216[5]), .I2(n554_adj_4859), 
            .I3(n51791), .O(n20055[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4851));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4850));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5143_8 (.CI(n51791), .I0(n20216[5]), .I1(n554_adj_4859), 
            .CO(n51792));
    SB_LUT4 add_5143_7_lut (.I0(GND_net), .I1(n20216[4]), .I2(n481_adj_4858), 
            .I3(n51790), .O(n20055[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4849));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5143_7 (.CI(n51790), .I0(n20216[4]), .I1(n481_adj_4858), 
            .CO(n51791));
    SB_LUT4 add_5143_6_lut (.I0(GND_net), .I1(n20216[3]), .I2(n408_adj_4857), 
            .I3(n51789), .O(n20055[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5143_6 (.CI(n51789), .I0(n20216[3]), .I1(n408_adj_4857), 
            .CO(n51790));
    SB_LUT4 add_5143_5_lut (.I0(GND_net), .I1(n20216[2]), .I2(n335_adj_4856), 
            .I3(n51788), .O(n20055[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5143_5 (.CI(n51788), .I0(n20216[2]), .I1(n335_adj_4856), 
            .CO(n51789));
    SB_LUT4 add_5143_4_lut (.I0(GND_net), .I1(n20216[1]), .I2(n262_adj_4855), 
            .I3(n51787), .O(n20055[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5143_4 (.CI(n51787), .I0(n20216[1]), .I1(n262_adj_4855), 
            .CO(n51788));
    SB_LUT4 add_5143_3_lut (.I0(GND_net), .I1(n20216[0]), .I2(n189_adj_4854), 
            .I3(n51786), .O(n20055[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5143_3 (.CI(n51786), .I0(n20216[0]), .I1(n189_adj_4854), 
            .CO(n51787));
    SB_LUT4 add_5143_2_lut (.I0(GND_net), .I1(n47_adj_4853), .I2(n116_adj_4852), 
            .I3(GND_net), .O(n20055[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5143_2 (.CI(GND_net), .I0(n47_adj_4853), .I1(n116_adj_4852), 
            .CO(n51786));
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4848));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51295_3_lut (.I0(n68310), .I1(n356[18]), .I2(n37_adj_4735), 
            .I3(GND_net), .O(n68311));   // verilog/motorControl.v(52[14:29])
    defparam i51295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4847));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4846));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4840));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4825));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4924_18_lut (.I0(GND_net), .I1(n17338[15]), .I2(GND_net), 
            .I3(n51766), .O(n16722[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4924_17_lut (.I0(GND_net), .I1(n17338[14]), .I2(GND_net), 
            .I3(n51765), .O(n16722[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_17 (.CI(n51765), .I0(n17338[14]), .I1(GND_net), 
            .CO(n51766));
    SB_LUT4 add_4924_16_lut (.I0(GND_net), .I1(n17338[13]), .I2(n1114_adj_4845), 
            .I3(n51764), .O(n16722[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4824));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4924_16 (.CI(n51764), .I0(n17338[13]), .I1(n1114_adj_4845), 
            .CO(n51765));
    SB_LUT4 add_4924_15_lut (.I0(GND_net), .I1(n17338[12]), .I2(n1041_adj_4843), 
            .I3(n51763), .O(n16722[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_15 (.CI(n51763), .I0(n17338[12]), .I1(n1041_adj_4843), 
            .CO(n51764));
    SB_LUT4 add_4924_14_lut (.I0(GND_net), .I1(n17338[11]), .I2(n968_adj_4842), 
            .I3(n51762), .O(n16722[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_14 (.CI(n51762), .I0(n17338[11]), .I1(n968_adj_4842), 
            .CO(n51763));
    SB_LUT4 add_4924_13_lut (.I0(GND_net), .I1(n17338[10]), .I2(n895_adj_4841), 
            .I3(n51761), .O(n16722[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4924_13 (.CI(n51761), .I0(n17338[10]), .I1(n895_adj_4841), 
            .CO(n51762));
    SB_LUT4 add_4924_12_lut (.I0(GND_net), .I1(n17338[9]), .I2(n822), 
            .I3(n51760), .O(n16722[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4924_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4823));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4817));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4816));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4814));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4813));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4811));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4809));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4795));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4794));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4791));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4786));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4785));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4784));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51253_3_lut (.I0(n68311), .I1(n356[19]), .I2(n39_adj_4695), 
            .I3(GND_net), .O(n68269));   // verilog/motorControl.v(52[14:29])
    defparam i51253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49171_4_lut (.I0(n43_adj_4742), .I1(n41_adj_4694), .I2(n39_adj_4695), 
            .I3(n68211), .O(n66187));
    defparam i49171_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51130_4_lut (.I0(n66656), .I1(n67666), .I2(n45_adj_4696), 
            .I3(n66183), .O(n68146));   // verilog/motorControl.v(52[14:29])
    defparam i51130_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49648_3_lut (.I0(n68269), .I1(n356[20]), .I2(n41_adj_4694), 
            .I3(GND_net), .O(n66664));   // verilog/motorControl.v(52[14:29])
    defparam i49648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51132_4_lut (.I0(n66664), .I1(n68146), .I2(n45_adj_4696), 
            .I3(n66187), .O(n68148));   // verilog/motorControl.v(52[14:29])
    defparam i51132_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49066_2_lut_4_lut (.I0(n356[21]), .I1(n436[21]), .I2(n356[9]), 
            .I3(n436[9]), .O(n66082));
    defparam i49066_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51133_3_lut (.I0(n68148), .I1(PWMLimit[23]), .I2(n356[23]), 
            .I3(GND_net), .O(n409));   // verilog/motorControl.v(52[14:29])
    defparam i51133_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n356[20]), .I1(n436[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4927));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4757));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49103_2_lut_4_lut (.I0(n356[16]), .I1(n436[16]), .I2(n356[7]), 
            .I3(n436[7]), .O(n66119));
    defparam i49103_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5151_9_lut (.I0(GND_net), .I1(n20280[6]), .I2(n630_adj_4839), 
            .I3(n52413), .O(n20136[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5151_8_lut (.I0(GND_net), .I1(n20280[5]), .I2(n557_adj_4838), 
            .I3(n52412), .O(n20136[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_8 (.CI(n52412), .I0(n20280[5]), .I1(n557_adj_4838), 
            .CO(n52413));
    SB_LUT4 add_5151_7_lut (.I0(GND_net), .I1(n20280[4]), .I2(n484_adj_4837), 
            .I3(n52411), .O(n20136[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_7 (.CI(n52411), .I0(n20280[4]), .I1(n484_adj_4837), 
            .CO(n52412));
    SB_LUT4 add_5151_6_lut (.I0(GND_net), .I1(n20280[3]), .I2(n411_adj_4836), 
            .I3(n52410), .O(n20136[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_6 (.CI(n52410), .I0(n20280[3]), .I1(n411_adj_4836), 
            .CO(n52411));
    SB_LUT4 add_5151_5_lut (.I0(GND_net), .I1(n20280[2]), .I2(n338_adj_4835), 
            .I3(n52409), .O(n20136[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_5 (.CI(n52409), .I0(n20280[2]), .I1(n338_adj_4835), 
            .CO(n52410));
    SB_LUT4 add_5151_4_lut (.I0(GND_net), .I1(n20280[1]), .I2(n265_adj_4834), 
            .I3(n52408), .O(n20136[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_4 (.CI(n52408), .I0(n20280[1]), .I1(n265_adj_4834), 
            .CO(n52409));
    SB_LUT4 add_5151_3_lut (.I0(GND_net), .I1(n20280[0]), .I2(n192_adj_4833), 
            .I3(n52407), .O(n20136[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_3 (.CI(n52407), .I0(n20280[0]), .I1(n192_adj_4833), 
            .CO(n52408));
    SB_LUT4 add_5151_2_lut (.I0(GND_net), .I1(n50_adj_4832), .I2(n119_adj_4831), 
            .I3(GND_net), .O(n20136[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_2 (.CI(GND_net), .I0(n50_adj_4832), .I1(n119_adj_4831), 
            .CO(n52407));
    SB_LUT4 mult_16_add_1225_24_lut (.I0(n49[23]), .I1(n11262[21]), .I2(GND_net), 
            .I3(n52406), .O(n10755[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_16_add_1225_23_lut (.I0(GND_net), .I1(n11262[20]), .I2(GND_net), 
            .I3(n52405), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_23 (.CI(n52405), .I0(n11262[20]), .I1(GND_net), 
            .CO(n52406));
    SB_LUT4 mult_16_add_1225_22_lut (.I0(GND_net), .I1(n11262[19]), .I2(GND_net), 
            .I3(n52404), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n356[19]), .I1(n436[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4928));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_16_add_1225_22 (.CI(n52404), .I0(n11262[19]), .I1(GND_net), 
            .CO(n52405));
    SB_LUT4 mult_16_add_1225_21_lut (.I0(GND_net), .I1(n11262[18]), .I2(GND_net), 
            .I3(n52403), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_21 (.CI(n52403), .I0(n11262[18]), .I1(GND_net), 
            .CO(n52404));
    SB_LUT4 mult_16_add_1225_20_lut (.I0(GND_net), .I1(n11262[17]), .I2(GND_net), 
            .I3(n52402), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_20 (.CI(n52402), .I0(n11262[17]), .I1(GND_net), 
            .CO(n52403));
    SB_LUT4 mult_16_add_1225_19_lut (.I0(GND_net), .I1(n11262[16]), .I2(GND_net), 
            .I3(n52401), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_19 (.CI(n52401), .I0(n11262[16]), .I1(GND_net), 
            .CO(n52402));
    SB_LUT4 mult_16_add_1225_18_lut (.I0(GND_net), .I1(n11262[15]), .I2(GND_net), 
            .I3(n52400), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_18 (.CI(n52400), .I0(n11262[15]), .I1(GND_net), 
            .CO(n52401));
    SB_LUT4 mult_16_add_1225_17_lut (.I0(GND_net), .I1(n11262[14]), .I2(GND_net), 
            .I3(n52399), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_17 (.CI(n52399), .I0(n11262[14]), .I1(GND_net), 
            .CO(n52400));
    SB_LUT4 mult_16_add_1225_16_lut (.I0(GND_net), .I1(n11262[13]), .I2(n1096_adj_4830), 
            .I3(n52398), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_16 (.CI(n52398), .I0(n11262[13]), .I1(n1096_adj_4830), 
            .CO(n52399));
    SB_LUT4 mult_16_add_1225_15_lut (.I0(GND_net), .I1(n11262[12]), .I2(n1023_adj_4829), 
            .I3(n52397), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_15 (.CI(n52397), .I0(n11262[12]), .I1(n1023_adj_4829), 
            .CO(n52398));
    SB_LUT4 mult_16_add_1225_14_lut (.I0(GND_net), .I1(n11262[11]), .I2(n950_adj_4828), 
            .I3(n52396), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_14 (.CI(n52396), .I0(n11262[11]), .I1(n950_adj_4828), 
            .CO(n52397));
    SB_LUT4 mult_16_add_1225_13_lut (.I0(GND_net), .I1(n11262[10]), .I2(n877_adj_4827), 
            .I3(n52395), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_13 (.CI(n52395), .I0(n11262[10]), .I1(n877_adj_4827), 
            .CO(n52396));
    SB_LUT4 mult_16_add_1225_12_lut (.I0(GND_net), .I1(n11262[9]), .I2(n804_adj_4826), 
            .I3(n52394), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_12 (.CI(n52394), .I0(n11262[9]), .I1(n804_adj_4826), 
            .CO(n52395));
    SB_LUT4 mult_16_add_1225_11_lut (.I0(GND_net), .I1(n11262[8]), .I2(n731_adj_4822), 
            .I3(n52393), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_11 (.CI(n52393), .I0(n11262[8]), .I1(n731_adj_4822), 
            .CO(n52394));
    SB_LUT4 mult_16_add_1225_10_lut (.I0(GND_net), .I1(n11262[7]), .I2(n658_adj_4821), 
            .I3(n52392), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_10 (.CI(n52392), .I0(n11262[7]), .I1(n658_adj_4821), 
            .CO(n52393));
    SB_LUT4 mult_16_add_1225_9_lut (.I0(GND_net), .I1(n11262[6]), .I2(n585_adj_4819), 
            .I3(n52391), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_9 (.CI(n52391), .I0(n11262[6]), .I1(n585_adj_4819), 
            .CO(n52392));
    SB_LUT4 mult_16_add_1225_8_lut (.I0(GND_net), .I1(n11262[5]), .I2(n512_adj_4818), 
            .I3(n52390), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_8 (.CI(n52390), .I0(n11262[5]), .I1(n512_adj_4818), 
            .CO(n52391));
    SB_LUT4 mult_16_add_1225_7_lut (.I0(GND_net), .I1(n11262[4]), .I2(n439_adj_4815), 
            .I3(n52389), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_7 (.CI(n52389), .I0(n11262[4]), .I1(n439_adj_4815), 
            .CO(n52390));
    SB_LUT4 mult_16_add_1225_6_lut (.I0(GND_net), .I1(n11262[3]), .I2(n366_adj_4812), 
            .I3(n52388), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_6 (.CI(n52388), .I0(n11262[3]), .I1(n366_adj_4812), 
            .CO(n52389));
    SB_LUT4 mult_16_add_1225_5_lut (.I0(GND_net), .I1(n11262[2]), .I2(n293_adj_4810), 
            .I3(n52387), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_5 (.CI(n52387), .I0(n11262[2]), .I1(n293_adj_4810), 
            .CO(n52388));
    SB_LUT4 mult_16_add_1225_4_lut (.I0(GND_net), .I1(n11262[1]), .I2(n220_adj_4808), 
            .I3(n52386), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_4 (.CI(n52386), .I0(n11262[1]), .I1(n220_adj_4808), 
            .CO(n52387));
    SB_LUT4 mult_16_add_1225_3_lut (.I0(GND_net), .I1(n11262[0]), .I2(n147_adj_4807), 
            .I3(n52385), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_3 (.CI(n52385), .I0(n11262[0]), .I1(n147_adj_4807), 
            .CO(n52386));
    SB_LUT4 mult_16_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4806), .I2(n74_adj_4805), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_2 (.CI(GND_net), .I0(n5_adj_4806), .I1(n74_adj_4805), 
            .CO(n52385));
    SB_LUT4 add_4449_23_lut (.I0(GND_net), .I1(n12924[20]), .I2(GND_net), 
            .I3(n52384), .O(n11262[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4449_22_lut (.I0(GND_net), .I1(n12924[19]), .I2(GND_net), 
            .I3(n52383), .O(n11262[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_22 (.CI(n52383), .I0(n12924[19]), .I1(GND_net), 
            .CO(n52384));
    SB_LUT4 add_4449_21_lut (.I0(GND_net), .I1(n12924[18]), .I2(GND_net), 
            .I3(n52382), .O(n11262[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_21 (.CI(n52382), .I0(n12924[18]), .I1(GND_net), 
            .CO(n52383));
    SB_LUT4 add_4449_20_lut (.I0(GND_net), .I1(n12924[17]), .I2(GND_net), 
            .I3(n52381), .O(n11262[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_20 (.CI(n52381), .I0(n12924[17]), .I1(GND_net), 
            .CO(n52382));
    SB_LUT4 add_4449_19_lut (.I0(GND_net), .I1(n12924[16]), .I2(GND_net), 
            .I3(n52380), .O(n11262[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_19 (.CI(n52380), .I0(n12924[16]), .I1(GND_net), 
            .CO(n52381));
    SB_LUT4 add_4449_18_lut (.I0(GND_net), .I1(n12924[15]), .I2(GND_net), 
            .I3(n52379), .O(n11262[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_18 (.CI(n52379), .I0(n12924[15]), .I1(GND_net), 
            .CO(n52380));
    SB_LUT4 add_4449_17_lut (.I0(GND_net), .I1(n12924[14]), .I2(GND_net), 
            .I3(n52378), .O(n11262[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_17 (.CI(n52378), .I0(n12924[14]), .I1(GND_net), 
            .CO(n52379));
    SB_LUT4 add_4449_16_lut (.I0(GND_net), .I1(n12924[13]), .I2(n1099_adj_4804), 
            .I3(n52377), .O(n11262[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_16 (.CI(n52377), .I0(n12924[13]), .I1(n1099_adj_4804), 
            .CO(n52378));
    SB_LUT4 add_4449_15_lut (.I0(GND_net), .I1(n12924[12]), .I2(n1026_adj_4803), 
            .I3(n52376), .O(n11262[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_15 (.CI(n52376), .I0(n12924[12]), .I1(n1026_adj_4803), 
            .CO(n52377));
    SB_LUT4 add_4449_14_lut (.I0(GND_net), .I1(n12924[11]), .I2(n953_adj_4802), 
            .I3(n52375), .O(n11262[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_14 (.CI(n52375), .I0(n12924[11]), .I1(n953_adj_4802), 
            .CO(n52376));
    SB_LUT4 add_4449_13_lut (.I0(GND_net), .I1(n12924[10]), .I2(n880_adj_4801), 
            .I3(n52374), .O(n11262[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_13 (.CI(n52374), .I0(n12924[10]), .I1(n880_adj_4801), 
            .CO(n52375));
    SB_LUT4 add_4449_12_lut (.I0(GND_net), .I1(n12924[9]), .I2(n807_adj_4800), 
            .I3(n52373), .O(n11262[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_12 (.CI(n52373), .I0(n12924[9]), .I1(n807_adj_4800), 
            .CO(n52374));
    SB_LUT4 add_4449_11_lut (.I0(GND_net), .I1(n12924[8]), .I2(n734_adj_4799), 
            .I3(n52372), .O(n11262[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_11 (.CI(n52372), .I0(n12924[8]), .I1(n734_adj_4799), 
            .CO(n52373));
    SB_LUT4 add_4449_10_lut (.I0(GND_net), .I1(n12924[7]), .I2(n661_adj_4798), 
            .I3(n52371), .O(n11262[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_10 (.CI(n52371), .I0(n12924[7]), .I1(n661_adj_4798), 
            .CO(n52372));
    SB_LUT4 add_4449_9_lut (.I0(GND_net), .I1(n12924[6]), .I2(n588_adj_4797), 
            .I3(n52370), .O(n11262[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_9 (.CI(n52370), .I0(n12924[6]), .I1(n588_adj_4797), 
            .CO(n52371));
    SB_LUT4 add_4449_8_lut (.I0(GND_net), .I1(n12924[5]), .I2(n515_adj_4796), 
            .I3(n52369), .O(n11262[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_8 (.CI(n52369), .I0(n12924[5]), .I1(n515_adj_4796), 
            .CO(n52370));
    SB_LUT4 add_4449_7_lut (.I0(GND_net), .I1(n12924[4]), .I2(n442_adj_4793), 
            .I3(n52368), .O(n11262[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_7 (.CI(n52368), .I0(n12924[4]), .I1(n442_adj_4793), 
            .CO(n52369));
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n356[22]), .I1(n436[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4929));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4449_6_lut (.I0(GND_net), .I1(n12924[3]), .I2(n369_adj_4792), 
            .I3(n52367), .O(n11262[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_6 (.CI(n52367), .I0(n12924[3]), .I1(n369_adj_4792), 
            .CO(n52368));
    SB_LUT4 add_4449_5_lut (.I0(GND_net), .I1(n12924[2]), .I2(n296_adj_4790), 
            .I3(n52366), .O(n11262[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_5 (.CI(n52366), .I0(n12924[2]), .I1(n296_adj_4790), 
            .CO(n52367));
    SB_LUT4 add_4449_4_lut (.I0(GND_net), .I1(n12924[1]), .I2(n223_adj_4789), 
            .I3(n52365), .O(n11262[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_4 (.CI(n52365), .I0(n12924[1]), .I1(n223_adj_4789), 
            .CO(n52366));
    SB_LUT4 add_4449_3_lut (.I0(GND_net), .I1(n12924[0]), .I2(n150_adj_4788), 
            .I3(n52364), .O(n11262[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_3 (.CI(n52364), .I0(n12924[0]), .I1(n150_adj_4788), 
            .CO(n52365));
    SB_LUT4 add_4449_2_lut (.I0(GND_net), .I1(n8_adj_4787), .I2(n77), 
            .I3(GND_net), .O(n11262[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4449_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4449_2 (.CI(GND_net), .I0(n8_adj_4787), .I1(n77), .CO(n52364));
    SB_LUT4 add_4742_22_lut (.I0(GND_net), .I1(n14183[19]), .I2(GND_net), 
            .I3(n52363), .O(n12924[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4742_21_lut (.I0(GND_net), .I1(n14183[18]), .I2(GND_net), 
            .I3(n52362), .O(n12924[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_21 (.CI(n52362), .I0(n14183[18]), .I1(GND_net), 
            .CO(n52363));
    SB_LUT4 add_4742_20_lut (.I0(GND_net), .I1(n14183[17]), .I2(GND_net), 
            .I3(n52361), .O(n12924[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_20 (.CI(n52361), .I0(n14183[17]), .I1(GND_net), 
            .CO(n52362));
    SB_LUT4 add_4742_19_lut (.I0(GND_net), .I1(n14183[16]), .I2(GND_net), 
            .I3(n52360), .O(n12924[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_19 (.CI(n52360), .I0(n14183[16]), .I1(GND_net), 
            .CO(n52361));
    SB_LUT4 add_4742_18_lut (.I0(GND_net), .I1(n14183[15]), .I2(GND_net), 
            .I3(n52359), .O(n12924[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_18 (.CI(n52359), .I0(n14183[15]), .I1(GND_net), 
            .CO(n52360));
    SB_LUT4 add_4742_17_lut (.I0(GND_net), .I1(n14183[14]), .I2(GND_net), 
            .I3(n52358), .O(n12924[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_17 (.CI(n52358), .I0(n14183[14]), .I1(GND_net), 
            .CO(n52359));
    SB_LUT4 add_4742_16_lut (.I0(GND_net), .I1(n14183[13]), .I2(n1102), 
            .I3(n52357), .O(n12924[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_16 (.CI(n52357), .I0(n14183[13]), .I1(n1102), .CO(n52358));
    SB_LUT4 add_4742_15_lut (.I0(GND_net), .I1(n14183[12]), .I2(n1029), 
            .I3(n52356), .O(n12924[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_15 (.CI(n52356), .I0(n14183[12]), .I1(n1029), .CO(n52357));
    SB_LUT4 add_4742_14_lut (.I0(GND_net), .I1(n14183[11]), .I2(n956), 
            .I3(n52355), .O(n12924[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_14 (.CI(n52355), .I0(n14183[11]), .I1(n956), .CO(n52356));
    SB_LUT4 add_4742_13_lut (.I0(GND_net), .I1(n14183[10]), .I2(n883), 
            .I3(n52354), .O(n12924[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_13 (.CI(n52354), .I0(n14183[10]), .I1(n883), .CO(n52355));
    SB_LUT4 add_4742_12_lut (.I0(GND_net), .I1(n14183[9]), .I2(n810), 
            .I3(n52353), .O(n12924[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_12 (.CI(n52353), .I0(n14183[9]), .I1(n810), .CO(n52354));
    SB_LUT4 add_4742_11_lut (.I0(GND_net), .I1(n14183[8]), .I2(n737), 
            .I3(n52352), .O(n12924[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_11 (.CI(n52352), .I0(n14183[8]), .I1(n737), .CO(n52353));
    SB_LUT4 add_4742_10_lut (.I0(GND_net), .I1(n14183[7]), .I2(n664), 
            .I3(n52351), .O(n12924[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_10 (.CI(n52351), .I0(n14183[7]), .I1(n664), .CO(n52352));
    SB_LUT4 add_4742_9_lut (.I0(GND_net), .I1(n14183[6]), .I2(n591), .I3(n52350), 
            .O(n12924[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_9 (.CI(n52350), .I0(n14183[6]), .I1(n591), .CO(n52351));
    SB_LUT4 add_4742_8_lut (.I0(GND_net), .I1(n14183[5]), .I2(n518), .I3(n52349), 
            .O(n12924[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_8 (.CI(n52349), .I0(n14183[5]), .I1(n518), .CO(n52350));
    SB_LUT4 add_4742_7_lut (.I0(GND_net), .I1(n14183[4]), .I2(n445_adj_4783), 
            .I3(n52348), .O(n12924[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_7 (.CI(n52348), .I0(n14183[4]), .I1(n445_adj_4783), 
            .CO(n52349));
    SB_LUT4 add_4742_6_lut (.I0(GND_net), .I1(n14183[3]), .I2(n372_adj_4782), 
            .I3(n52347), .O(n12924[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_6 (.CI(n52347), .I0(n14183[3]), .I1(n372_adj_4782), 
            .CO(n52348));
    SB_LUT4 add_4742_5_lut (.I0(GND_net), .I1(n14183[2]), .I2(n299_adj_4781), 
            .I3(n52346), .O(n12924[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_5 (.CI(n52346), .I0(n14183[2]), .I1(n299_adj_4781), 
            .CO(n52347));
    SB_LUT4 add_4742_4_lut (.I0(GND_net), .I1(n14183[1]), .I2(n226_adj_4780), 
            .I3(n52345), .O(n12924[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_4 (.CI(n52345), .I0(n14183[1]), .I1(n226_adj_4780), 
            .CO(n52346));
    SB_LUT4 add_4742_3_lut (.I0(GND_net), .I1(n14183[0]), .I2(n153_adj_4779), 
            .I3(n52344), .O(n12924[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_3 (.CI(n52344), .I0(n14183[0]), .I1(n153_adj_4779), 
            .CO(n52345));
    SB_LUT4 add_4742_2_lut (.I0(GND_net), .I1(n11_adj_4778), .I2(n80), 
            .I3(GND_net), .O(n12924[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4742_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4742_2 (.CI(GND_net), .I0(n11_adj_4778), .I1(n80), .CO(n52344));
    SB_LUT4 add_4799_21_lut (.I0(GND_net), .I1(n15295[18]), .I2(GND_net), 
            .I3(n52343), .O(n14183[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4799_20_lut (.I0(GND_net), .I1(n15295[17]), .I2(GND_net), 
            .I3(n52342), .O(n14183[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_20 (.CI(n52342), .I0(n15295[17]), .I1(GND_net), 
            .CO(n52343));
    SB_LUT4 add_4799_19_lut (.I0(GND_net), .I1(n15295[16]), .I2(GND_net), 
            .I3(n52341), .O(n14183[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_19 (.CI(n52341), .I0(n15295[16]), .I1(GND_net), 
            .CO(n52342));
    SB_LUT4 add_4799_18_lut (.I0(GND_net), .I1(n15295[15]), .I2(GND_net), 
            .I3(n52340), .O(n14183[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_18 (.CI(n52340), .I0(n15295[15]), .I1(GND_net), 
            .CO(n52341));
    SB_LUT4 add_4799_17_lut (.I0(GND_net), .I1(n15295[14]), .I2(GND_net), 
            .I3(n52339), .O(n14183[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_17 (.CI(n52339), .I0(n15295[14]), .I1(GND_net), 
            .CO(n52340));
    SB_LUT4 add_4799_16_lut (.I0(GND_net), .I1(n15295[13]), .I2(n1105), 
            .I3(n52338), .O(n14183[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_16 (.CI(n52338), .I0(n15295[13]), .I1(n1105), .CO(n52339));
    SB_LUT4 add_4799_15_lut (.I0(GND_net), .I1(n15295[12]), .I2(n1032), 
            .I3(n52337), .O(n14183[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_15 (.CI(n52337), .I0(n15295[12]), .I1(n1032), .CO(n52338));
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n356[8]), .I1(n436[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4930));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4799_14_lut (.I0(GND_net), .I1(n15295[11]), .I2(n959), 
            .I3(n52336), .O(n14183[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_14 (.CI(n52336), .I0(n15295[11]), .I1(n959), .CO(n52337));
    SB_LUT4 add_4799_13_lut (.I0(GND_net), .I1(n15295[10]), .I2(n886), 
            .I3(n52335), .O(n14183[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_13 (.CI(n52335), .I0(n15295[10]), .I1(n886), .CO(n52336));
    SB_LUT4 add_4799_12_lut (.I0(GND_net), .I1(n15295[9]), .I2(n813), 
            .I3(n52334), .O(n14183[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_12 (.CI(n52334), .I0(n15295[9]), .I1(n813), .CO(n52335));
    SB_LUT4 add_4799_11_lut (.I0(GND_net), .I1(n15295[8]), .I2(n740), 
            .I3(n52333), .O(n14183[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_11 (.CI(n52333), .I0(n15295[8]), .I1(n740), .CO(n52334));
    SB_LUT4 add_4799_10_lut (.I0(GND_net), .I1(n15295[7]), .I2(n667), 
            .I3(n52332), .O(n14183[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_10 (.CI(n52332), .I0(n15295[7]), .I1(n667), .CO(n52333));
    SB_LUT4 add_4799_9_lut (.I0(GND_net), .I1(n15295[6]), .I2(n594), .I3(n52331), 
            .O(n14183[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_9 (.CI(n52331), .I0(n15295[6]), .I1(n594), .CO(n52332));
    SB_LUT4 add_4799_8_lut (.I0(GND_net), .I1(n15295[5]), .I2(n521), .I3(n52330), 
            .O(n14183[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_8 (.CI(n52330), .I0(n15295[5]), .I1(n521), .CO(n52331));
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n356[9]), .I1(n436[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4931));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4799_7_lut (.I0(GND_net), .I1(n15295[4]), .I2(n448_adj_4777), 
            .I3(n52329), .O(n14183[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_7 (.CI(n52329), .I0(n15295[4]), .I1(n448_adj_4777), 
            .CO(n52330));
    SB_LUT4 add_4799_6_lut (.I0(GND_net), .I1(n15295[3]), .I2(n375_adj_4776), 
            .I3(n52328), .O(n14183[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_6 (.CI(n52328), .I0(n15295[3]), .I1(n375_adj_4776), 
            .CO(n52329));
    SB_LUT4 add_4799_5_lut (.I0(GND_net), .I1(n15295[2]), .I2(n302_adj_4773), 
            .I3(n52327), .O(n14183[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_5 (.CI(n52327), .I0(n15295[2]), .I1(n302_adj_4773), 
            .CO(n52328));
    SB_LUT4 add_4799_4_lut (.I0(GND_net), .I1(n15295[1]), .I2(n229_adj_4772), 
            .I3(n52326), .O(n14183[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_4 (.CI(n52326), .I0(n15295[1]), .I1(n229_adj_4772), 
            .CO(n52327));
    SB_LUT4 add_4799_3_lut (.I0(GND_net), .I1(n15295[0]), .I2(n156_adj_4771), 
            .I3(n52325), .O(n14183[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_3 (.CI(n52325), .I0(n15295[0]), .I1(n156_adj_4771), 
            .CO(n52326));
    SB_LUT4 add_4799_2_lut (.I0(GND_net), .I1(n14_adj_4770), .I2(n83), 
            .I3(GND_net), .O(n14183[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4799_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4799_2 (.CI(GND_net), .I0(n14_adj_4770), .I1(n83), .CO(n52325));
    SB_LUT4 add_4850_20_lut (.I0(GND_net), .I1(n16271[17]), .I2(GND_net), 
            .I3(n52324), .O(n15295[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_19_lut (.I0(GND_net), .I1(n16271[16]), .I2(GND_net), 
            .I3(n52323), .O(n15295[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_19 (.CI(n52323), .I0(n16271[16]), .I1(GND_net), 
            .CO(n52324));
    SB_LUT4 add_4850_18_lut (.I0(GND_net), .I1(n16271[15]), .I2(GND_net), 
            .I3(n52322), .O(n15295[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_18 (.CI(n52322), .I0(n16271[15]), .I1(GND_net), 
            .CO(n52323));
    SB_LUT4 add_4850_17_lut (.I0(GND_net), .I1(n16271[14]), .I2(GND_net), 
            .I3(n52321), .O(n15295[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_17 (.CI(n52321), .I0(n16271[14]), .I1(GND_net), 
            .CO(n52322));
    SB_LUT4 add_4850_16_lut (.I0(GND_net), .I1(n16271[13]), .I2(n1108), 
            .I3(n52320), .O(n15295[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_16 (.CI(n52320), .I0(n16271[13]), .I1(n1108), .CO(n52321));
    SB_LUT4 add_4850_15_lut (.I0(GND_net), .I1(n16271[12]), .I2(n1035), 
            .I3(n52319), .O(n15295[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4850_15 (.CI(n52319), .I0(n16271[12]), .I1(n1035), .CO(n52320));
    SB_LUT4 add_4850_14_lut (.I0(GND_net), .I1(n16271[11]), .I2(n962), 
            .I3(n52318), .O(n15295[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_14 (.CI(n52318), .I0(n16271[11]), .I1(n962), .CO(n52319));
    SB_LUT4 add_4850_13_lut (.I0(GND_net), .I1(n16271[10]), .I2(n889), 
            .I3(n52317), .O(n15295[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_13 (.CI(n52317), .I0(n16271[10]), .I1(n889), .CO(n52318));
    SB_LUT4 add_4850_12_lut (.I0(GND_net), .I1(n16271[9]), .I2(n816), 
            .I3(n52316), .O(n15295[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_12 (.CI(n52316), .I0(n16271[9]), .I1(n816), .CO(n52317));
    SB_LUT4 add_4850_11_lut (.I0(GND_net), .I1(n16271[8]), .I2(n743), 
            .I3(n52315), .O(n15295[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_11 (.CI(n52315), .I0(n16271[8]), .I1(n743), .CO(n52316));
    SB_LUT4 add_4850_10_lut (.I0(GND_net), .I1(n16271[7]), .I2(n670), 
            .I3(n52314), .O(n15295[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_10 (.CI(n52314), .I0(n16271[7]), .I1(n670), .CO(n52315));
    SB_LUT4 add_4850_9_lut (.I0(GND_net), .I1(n16271[6]), .I2(n597), .I3(n52313), 
            .O(n15295[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_9 (.CI(n52313), .I0(n16271[6]), .I1(n597), .CO(n52314));
    SB_LUT4 add_4850_8_lut (.I0(GND_net), .I1(n16271[5]), .I2(n524), .I3(n52312), 
            .O(n15295[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_8 (.CI(n52312), .I0(n16271[5]), .I1(n524), .CO(n52313));
    SB_LUT4 add_4850_7_lut (.I0(GND_net), .I1(n16271[4]), .I2(n451_adj_4767), 
            .I3(n52311), .O(n15295[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_7 (.CI(n52311), .I0(n16271[4]), .I1(n451_adj_4767), 
            .CO(n52312));
    SB_LUT4 add_4850_6_lut (.I0(GND_net), .I1(n16271[3]), .I2(n378_adj_4766), 
            .I3(n52310), .O(n15295[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_6 (.CI(n52310), .I0(n16271[3]), .I1(n378_adj_4766), 
            .CO(n52311));
    SB_LUT4 add_4850_5_lut (.I0(GND_net), .I1(n16271[2]), .I2(n305_adj_4765), 
            .I3(n52309), .O(n15295[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_5 (.CI(n52309), .I0(n16271[2]), .I1(n305_adj_4765), 
            .CO(n52310));
    SB_LUT4 add_4850_4_lut (.I0(GND_net), .I1(n16271[1]), .I2(n232), .I3(n52308), 
            .O(n15295[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_4 (.CI(n52308), .I0(n16271[1]), .I1(n232), .CO(n52309));
    SB_LUT4 add_4850_3_lut (.I0(GND_net), .I1(n16271[0]), .I2(n159_adj_4762), 
            .I3(n52307), .O(n15295[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_3 (.CI(n52307), .I0(n16271[0]), .I1(n159_adj_4762), 
            .CO(n52308));
    SB_LUT4 add_4850_2_lut (.I0(GND_net), .I1(n17_adj_4761), .I2(n86), 
            .I3(GND_net), .O(n15295[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_2 (.CI(GND_net), .I0(n17_adj_4761), .I1(n86), .CO(n52307));
    SB_LUT4 add_4897_19_lut (.I0(GND_net), .I1(n17045[16]), .I2(GND_net), 
            .I3(n52306), .O(n16271[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4751));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4897_18_lut (.I0(GND_net), .I1(n17045[15]), .I2(GND_net), 
            .I3(n52305), .O(n16271[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_18 (.CI(n52305), .I0(n17045[15]), .I1(GND_net), 
            .CO(n52306));
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4897_17_lut (.I0(GND_net), .I1(n17045[14]), .I2(GND_net), 
            .I3(n52304), .O(n16271[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_17 (.CI(n52304), .I0(n17045[14]), .I1(GND_net), 
            .CO(n52305));
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n356[21]), .I1(n436[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4932));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4897_16_lut (.I0(GND_net), .I1(n17045[13]), .I2(n1111), 
            .I3(n52303), .O(n16271[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_16 (.CI(n52303), .I0(n17045[13]), .I1(n1111), .CO(n52304));
    SB_LUT4 add_4897_15_lut (.I0(GND_net), .I1(n17045[12]), .I2(n1038), 
            .I3(n52302), .O(n16271[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_15 (.CI(n52302), .I0(n17045[12]), .I1(n1038), .CO(n52303));
    SB_LUT4 add_4897_14_lut (.I0(GND_net), .I1(n17045[11]), .I2(n965), 
            .I3(n52301), .O(n16271[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_14 (.CI(n52301), .I0(n17045[11]), .I1(n965), .CO(n52302));
    SB_LUT4 add_4897_13_lut (.I0(GND_net), .I1(n17045[10]), .I2(n892), 
            .I3(n52300), .O(n16271[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_13 (.CI(n52300), .I0(n17045[10]), .I1(n892), .CO(n52301));
    SB_LUT4 add_4897_12_lut (.I0(GND_net), .I1(n17045[9]), .I2(n819), 
            .I3(n52299), .O(n16271[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_12 (.CI(n52299), .I0(n17045[9]), .I1(n819), .CO(n52300));
    SB_LUT4 add_4897_11_lut (.I0(GND_net), .I1(n17045[8]), .I2(n746), 
            .I3(n52298), .O(n16271[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_11 (.CI(n52298), .I0(n17045[8]), .I1(n746), .CO(n52299));
    SB_LUT4 add_4897_10_lut (.I0(GND_net), .I1(n17045[7]), .I2(n673), 
            .I3(n52297), .O(n16271[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_10 (.CI(n52297), .I0(n17045[7]), .I1(n673), .CO(n52298));
    SB_LUT4 add_4897_9_lut (.I0(GND_net), .I1(n17045[6]), .I2(n600), .I3(n52296), 
            .O(n16271[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_9 (.CI(n52296), .I0(n17045[6]), .I1(n600), .CO(n52297));
    SB_LUT4 add_4897_8_lut (.I0(GND_net), .I1(n17045[5]), .I2(n527), .I3(n52295), 
            .O(n16271[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_8 (.CI(n52295), .I0(n17045[5]), .I1(n527), .CO(n52296));
    SB_LUT4 add_4897_7_lut (.I0(GND_net), .I1(n17045[4]), .I2(n454_adj_4758), 
            .I3(n52294), .O(n16271[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_7 (.CI(n52294), .I0(n17045[4]), .I1(n454_adj_4758), 
            .CO(n52295));
    SB_LUT4 add_4897_6_lut (.I0(GND_net), .I1(n17045[3]), .I2(n381), .I3(n52293), 
            .O(n16271[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_6 (.CI(n52293), .I0(n17045[3]), .I1(n381), .CO(n52294));
    SB_LUT4 add_4897_5_lut (.I0(GND_net), .I1(n17045[2]), .I2(n308), .I3(n52292), 
            .O(n16271[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_5 (.CI(n52292), .I0(n17045[2]), .I1(n308), .CO(n52293));
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4750));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4897_4_lut (.I0(GND_net), .I1(n17045[1]), .I2(n235), .I3(n52291), 
            .O(n16271[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_4 (.CI(n52291), .I0(n17045[1]), .I1(n235), .CO(n52292));
    SB_LUT4 add_4897_3_lut (.I0(GND_net), .I1(n17045[0]), .I2(n162_adj_4755), 
            .I3(n52290), .O(n16271[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_3 (.CI(n52290), .I0(n17045[0]), .I1(n162_adj_4755), 
            .CO(n52291));
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4897_2_lut (.I0(GND_net), .I1(n20_adj_4753), .I2(n89), 
            .I3(GND_net), .O(n16271[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_2 (.CI(GND_net), .I0(n20_adj_4753), .I1(n89), .CO(n52290));
    SB_LUT4 add_4941_18_lut (.I0(GND_net), .I1(n17626[15]), .I2(GND_net), 
            .I3(n52289), .O(n17045[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4941_17_lut (.I0(GND_net), .I1(n17626[14]), .I2(GND_net), 
            .I3(n52288), .O(n17045[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_17 (.CI(n52288), .I0(n17626[14]), .I1(GND_net), 
            .CO(n52289));
    SB_LUT4 add_4941_16_lut (.I0(GND_net), .I1(n17626[13]), .I2(n1114), 
            .I3(n52287), .O(n17045[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_16 (.CI(n52287), .I0(n17626[13]), .I1(n1114), .CO(n52288));
    SB_LUT4 add_4941_15_lut (.I0(GND_net), .I1(n17626[12]), .I2(n1041), 
            .I3(n52286), .O(n17045[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_15 (.CI(n52286), .I0(n17626[12]), .I1(n1041), .CO(n52287));
    SB_LUT4 add_4941_14_lut (.I0(GND_net), .I1(n17626[11]), .I2(n968), 
            .I3(n52285), .O(n17045[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4941_14 (.CI(n52285), .I0(n17626[11]), .I1(n968), .CO(n52286));
    SB_LUT4 add_4941_13_lut (.I0(GND_net), .I1(n17626[10]), .I2(n895), 
            .I3(n52284), .O(n17045[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_13 (.CI(n52284), .I0(n17626[10]), .I1(n895), .CO(n52285));
    SB_LUT4 add_4941_12_lut (.I0(GND_net), .I1(n17626[9]), .I2(n822_adj_4748), 
            .I3(n52283), .O(n17045[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_12 (.CI(n52283), .I0(n17626[9]), .I1(n822_adj_4748), 
            .CO(n52284));
    SB_LUT4 add_4941_11_lut (.I0(GND_net), .I1(n17626[8]), .I2(n749_adj_4747), 
            .I3(n52282), .O(n17045[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_11 (.CI(n52282), .I0(n17626[8]), .I1(n749_adj_4747), 
            .CO(n52283));
    SB_LUT4 add_4941_10_lut (.I0(GND_net), .I1(n17626[7]), .I2(n676_adj_4746), 
            .I3(n52281), .O(n17045[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_10 (.CI(n52281), .I0(n17626[7]), .I1(n676_adj_4746), 
            .CO(n52282));
    SB_LUT4 add_4941_9_lut (.I0(GND_net), .I1(n17626[6]), .I2(n603_adj_4745), 
            .I3(n52280), .O(n17045[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_9 (.CI(n52280), .I0(n17626[6]), .I1(n603_adj_4745), 
            .CO(n52281));
    SB_LUT4 add_4941_8_lut (.I0(GND_net), .I1(n17626[5]), .I2(n530_adj_4744), 
            .I3(n52279), .O(n17045[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_8 (.CI(n52279), .I0(n17626[5]), .I1(n530_adj_4744), 
            .CO(n52280));
    SB_LUT4 add_4941_7_lut (.I0(GND_net), .I1(n17626[4]), .I2(n457_adj_4743), 
            .I3(n52278), .O(n17045[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_7 (.CI(n52278), .I0(n17626[4]), .I1(n457_adj_4743), 
            .CO(n52279));
    SB_LUT4 add_4941_6_lut (.I0(GND_net), .I1(n17626[3]), .I2(n384_adj_4741), 
            .I3(n52277), .O(n17045[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_6 (.CI(n52277), .I0(n17626[3]), .I1(n384_adj_4741), 
            .CO(n52278));
    SB_LUT4 add_4941_5_lut (.I0(GND_net), .I1(n17626[2]), .I2(n311_adj_4740), 
            .I3(n52276), .O(n17045[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_5 (.CI(n52276), .I0(n17626[2]), .I1(n311_adj_4740), 
            .CO(n52277));
    SB_LUT4 add_4941_4_lut (.I0(GND_net), .I1(n17626[1]), .I2(n238_adj_4738), 
            .I3(n52275), .O(n17045[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4941_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4941_4 (.CI(n52275), .I0(n17626[1]), .I1(n238_adj_4738), 
            .CO(n52276));
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4674));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n356[16]), .I1(n436[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4933));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n363), .I1(n436[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4934));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n356[18]), .I1(n436[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4935));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n356[13]), .I1(n436[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4936));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n356[14]), .I1(n436[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4937));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n356[15]), .I1(n436[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4938));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n356[10]), .I1(n436[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4939));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4665));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n356[11]), .I1(n436[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4940));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n356[12]), .I1(n436[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4941));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49127_4_lut (.I0(n21_adj_4939), .I1(n19_adj_4931), .I2(n17_adj_4930), 
            .I3(n9_adj_4703), .O(n66143));
    defparam i49127_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49115_4_lut (.I0(n27_adj_4936), .I1(n15_adj_4693), .I2(n13_adj_4705), 
            .I3(n11_adj_4704), .O(n66131));
    defparam i49115_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n436[7]), .I1(n436[16]), .I2(n33_adj_4933), 
            .I3(GND_net), .O(n12_adj_4942));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4734));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4733));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n436[5]), .I1(n436[6]), .I2(n13_adj_4705), 
            .I3(GND_net), .O(n10_adj_4943));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12_adj_4942), .I1(n436[17]), .I2(n35_adj_4934), 
            .I3(GND_net), .O(n30_adj_4944));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4730));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11813_3_lut (.I0(n356[1]), .I1(n436[1]), .I2(n9649), .I3(GND_net), 
            .O(n27546));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50022_4_lut (.I0(n13_adj_4705), .I1(n11_adj_4704), .I2(n9_adj_4703), 
            .I3(n66173), .O(n67038));
    defparam i50022_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i23425_4_lut (.I0(PWMLimit[1]), .I1(n61055), .I2(n27546), 
            .I3(n9647), .O(n1[1]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23425_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11808_3_lut (.I0(n356[2]), .I1(n436[2]), .I2(n9649), .I3(GND_net), 
            .O(n27541));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23424_4_lut (.I0(PWMLimit[2]), .I1(n61055), .I2(n27541), 
            .I3(n9647), .O(n1[2]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23424_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11803_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n9649), .I3(GND_net), 
            .O(n27536));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23423_4_lut (.I0(PWMLimit[3]), .I1(n61055), .I2(n27536), 
            .I3(n9647), .O(n1[3]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23423_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11798_3_lut (.I0(n356[4]), .I1(n436[4]), .I2(n9649), .I3(GND_net), 
            .O(n27531));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23422_4_lut (.I0(PWMLimit[4]), .I1(n61055), .I2(n27531), 
            .I3(n9647), .O(n1[4]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23422_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11793_3_lut (.I0(n356[5]), .I1(n436[5]), .I2(n9649), .I3(GND_net), 
            .O(n27526));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23421_4_lut (.I0(PWMLimit[5]), .I1(n61055), .I2(n27526), 
            .I3(n9647), .O(n1[5]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23421_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i50012_4_lut (.I0(n19_adj_4931), .I1(n17_adj_4930), .I2(n15_adj_4693), 
            .I3(n67038), .O(n67028));
    defparam i50012_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51056_4_lut (.I0(n25_adj_4941), .I1(n23_adj_4940), .I2(n21_adj_4939), 
            .I3(n67028), .O(n68072));
    defparam i51056_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50465_4_lut (.I0(n31_adj_4938), .I1(n29_adj_4937), .I2(n27_adj_4936), 
            .I3(n68072), .O(n67481));
    defparam i50465_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i11788_3_lut (.I0(n356[6]), .I1(n436[6]), .I2(n9649), .I3(GND_net), 
            .O(n27521));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51189_4_lut (.I0(n37_adj_4935), .I1(n35_adj_4934), .I2(n33_adj_4933), 
            .I3(n67481), .O(n68205));
    defparam i51189_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23420_4_lut (.I0(PWMLimit[6]), .I1(n61055), .I2(n27521), 
            .I3(n9647), .O(n1[6]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23420_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i50813_3_lut (.I0(n6_adj_4945), .I1(n436[10]), .I2(n21_adj_4939), 
            .I3(GND_net), .O(n67829));   // verilog/motorControl.v(54[23:39])
    defparam i50813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n436[9]), .I1(n436[21]), .I2(n43_adj_4932), 
            .I3(GND_net), .O(n16_adj_4946));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11783_3_lut (.I0(n356[7]), .I1(n436[7]), .I2(n9649), .I3(GND_net), 
            .O(n27516));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23419_4_lut (.I0(PWMLimit[7]), .I1(n61055), .I2(n27516), 
            .I3(n9647), .O(n1[7]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23419_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11778_3_lut (.I0(n356[8]), .I1(n436[8]), .I2(n9649), .I3(GND_net), 
            .O(n27511));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n436[4]), .I1(n436[8]), .I2(n17_adj_4930), 
            .I3(GND_net), .O(n8_adj_4947));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23418_4_lut (.I0(PWMLimit[8]), .I1(n61055), .I2(n27511), 
            .I3(n9647), .O(n1[8]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23418_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11773_3_lut (.I0(n356[9]), .I1(n436[9]), .I2(n9649), .I3(GND_net), 
            .O(n27506));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23417_4_lut (.I0(PWMLimit[9]), .I1(n61055), .I2(n27506), 
            .I3(n9647), .O(n1[9]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23417_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11768_3_lut (.I0(n356[10]), .I1(n436[10]), .I2(n9649), .I3(GND_net), 
            .O(n27501));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_4946), .I1(n436[22]), .I2(n45_adj_4929), 
            .I3(GND_net), .O(n24_adj_4948));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50814_3_lut (.I0(n67829), .I1(n436[11]), .I2(n23_adj_4940), 
            .I3(GND_net), .O(n67830));   // verilog/motorControl.v(54[23:39])
    defparam i50814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23416_4_lut (.I0(PWMLimit[10]), .I1(n61055), .I2(n27501), 
            .I3(n9647), .O(n1[10]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23416_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11763_3_lut (.I0(n356[11]), .I1(n436[11]), .I2(n9649), .I3(GND_net), 
            .O(n27496));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23415_4_lut (.I0(PWMLimit[11]), .I1(n61055), .I2(n27496), 
            .I3(n9647), .O(n1[11]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23415_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i49072_4_lut (.I0(n43_adj_4932), .I1(n25_adj_4941), .I2(n23_adj_4940), 
            .I3(n66143), .O(n66088));
    defparam i49072_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i11486_3_lut (.I0(n356[0]), .I1(n436[0]), .I2(n9649), .I3(GND_net), 
            .O(n27219));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50652_4_lut (.I0(n24_adj_4948), .I1(n8_adj_4947), .I2(n45_adj_4929), 
            .I3(n66082), .O(n67668));   // verilog/motorControl.v(54[23:39])
    defparam i50652_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i11758_3_lut (.I0(n356[12]), .I1(n436[12]), .I2(n9649), .I3(GND_net), 
            .O(n27491));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23414_4_lut (.I0(PWMLimit[12]), .I1(n61055), .I2(n27491), 
            .I3(n9647), .O(n1[12]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23414_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11753_3_lut (.I0(n356[13]), .I1(n436[13]), .I2(n9649), .I3(GND_net), 
            .O(n27486));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49650_3_lut (.I0(n67830), .I1(n436[12]), .I2(n25_adj_4941), 
            .I3(GND_net), .O(n66666));   // verilog/motorControl.v(54[23:39])
    defparam i49650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23413_4_lut (.I0(PWMLimit[13]), .I1(n61055), .I2(n27486), 
            .I3(n9647), .O(n1[13]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23413_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4638));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4637));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4636));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11748_3_lut (.I0(n356[14]), .I1(n436[14]), .I2(n9649), .I3(GND_net), 
            .O(n27481));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23412_4_lut (.I0(PWMLimit[14]), .I1(n61055), .I2(n27481), 
            .I3(n9647), .O(n1[14]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23412_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i23272_4_lut (.I0(PWMLimit[0]), .I1(n61055), .I2(n27219), 
            .I3(n9647), .O(n1[0]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23272_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_25_i4_4_lut (.I0(n436[0]), .I1(n436[1]), .I2(n356[1]), 
            .I3(n356[0]), .O(n4_adj_4949));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i11743_3_lut (.I0(n356[15]), .I1(n436[15]), .I2(n9649), .I3(GND_net), 
            .O(n27476));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23411_4_lut (.I0(PWMLimit[15]), .I1(n61055), .I2(n27476), 
            .I3(n9647), .O(n1[15]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23411_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11738_3_lut (.I0(n356[16]), .I1(n436[16]), .I2(n9649), .I3(GND_net), 
            .O(n27471));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23410_4_lut (.I0(PWMLimit[16]), .I1(n61055), .I2(n27471), 
            .I3(n9647), .O(n1[16]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23410_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11733_3_lut (.I0(n363), .I1(n436[17]), .I2(n9649), .I3(GND_net), 
            .O(n27466));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23408_4_lut (.I0(PWMLimit[17]), .I1(n61055), .I2(n27466), 
            .I3(n9647), .O(n1[17]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23408_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i50811_3_lut (.I0(n4_adj_4949), .I1(n436[13]), .I2(n27_adj_4936), 
            .I3(GND_net), .O(n67827));   // verilog/motorControl.v(54[23:39])
    defparam i50811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11728_3_lut (.I0(n356[18]), .I1(n436[18]), .I2(n9649), .I3(GND_net), 
            .O(n27461));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23407_4_lut (.I0(PWMLimit[18]), .I1(n61055), .I2(n27461), 
            .I3(n9647), .O(n1[18]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23407_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i50812_3_lut (.I0(n67827), .I1(n436[14]), .I2(n29_adj_4937), 
            .I3(GND_net), .O(n67828));   // verilog/motorControl.v(54[23:39])
    defparam i50812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49107_4_lut (.I0(n33_adj_4933), .I1(n31_adj_4938), .I2(n29_adj_4937), 
            .I3(n66131), .O(n66123));
    defparam i49107_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i11723_3_lut (.I0(n356[19]), .I1(n436[19]), .I2(n9649), .I3(GND_net), 
            .O(n27456));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23406_4_lut (.I0(PWMLimit[19]), .I1(n61055), .I2(n27456), 
            .I3(n9647), .O(n1[19]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23406_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11718_3_lut (.I0(n356[20]), .I1(n436[20]), .I2(n9649), .I3(GND_net), 
            .O(n27451));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23405_4_lut (.I0(PWMLimit[20]), .I1(n61055), .I2(n27451), 
            .I3(n9647), .O(n1[20]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23405_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i51161_4_lut (.I0(n30_adj_4944), .I1(n10_adj_4943), .I2(n35_adj_4934), 
            .I3(n66119), .O(n68177));   // verilog/motorControl.v(54[23:39])
    defparam i51161_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49652_3_lut (.I0(n67828), .I1(n436[15]), .I2(n31_adj_4938), 
            .I3(GND_net), .O(n66668));   // verilog/motorControl.v(54[23:39])
    defparam i49652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51296_4_lut (.I0(n66668), .I1(n68177), .I2(n35_adj_4934), 
            .I3(n66123), .O(n68312));   // verilog/motorControl.v(54[23:39])
    defparam i51296_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11713_3_lut (.I0(n356[21]), .I1(n436[21]), .I2(n9649), .I3(GND_net), 
            .O(n27446));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23404_4_lut (.I0(PWMLimit[21]), .I1(n61055), .I2(n27446), 
            .I3(n9647), .O(n1[21]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23404_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i51297_3_lut (.I0(n68312), .I1(n436[18]), .I2(n37_adj_4935), 
            .I3(GND_net), .O(n68313));   // verilog/motorControl.v(54[23:39])
    defparam i51297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11708_3_lut (.I0(n356[22]), .I1(n436[22]), .I2(n9649), .I3(GND_net), 
            .O(n27441));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23403_4_lut (.I0(PWMLimit[22]), .I1(n61055), .I2(n27441), 
            .I3(n9647), .O(n1[22]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23403_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51251_3_lut (.I0(n68313), .I1(n436[19]), .I2(n39_adj_4928), 
            .I3(GND_net), .O(n68267));   // verilog/motorControl.v(54[23:39])
    defparam i51251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49076_4_lut (.I0(n43_adj_4932), .I1(n41_adj_4927), .I2(n39_adj_4928), 
            .I3(n68205), .O(n66092));
    defparam i49076_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4634));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4633));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11703_3_lut (.I0(n356[23]), .I1(n436[23]), .I2(n9649), .I3(GND_net), 
            .O(n27436));   // verilog/motorControl.v(41[14] 61[8])
    defparam i11703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23402_4_lut (.I0(PWMLimit[23]), .I1(n61055), .I2(n27436), 
            .I3(n9647), .O(n1[23]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i23402_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i51134_4_lut (.I0(n66666), .I1(n67668), .I2(n45_adj_4929), 
            .I3(n66088), .O(n68150));   // verilog/motorControl.v(54[23:39])
    defparam i51134_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49658_3_lut (.I0(n68267), .I1(n436[20]), .I2(n41_adj_4927), 
            .I3(GND_net), .O(n66674));   // verilog/motorControl.v(54[23:39])
    defparam i49658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4632));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4631));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4630));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4628));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [11]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4564));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4563));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51136_4_lut (.I0(n66674), .I1(n68150), .I2(n45_adj_4929), 
            .I3(n66092), .O(n68152));   // verilog/motorControl.v(54[23:39])
    defparam i51136_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4627));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4626));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4625));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4562));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51137_3_lut (.I0(n68152), .I1(n356[23]), .I2(n436[23]), .I3(GND_net), 
            .O(n68153));   // verilog/motorControl.v(54[23:39])
    defparam i51137_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4561));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4326_3_lut (.I0(control_update), .I1(n409), .I2(n68153), 
            .I3(GND_net), .O(n9649));   // verilog/motorControl.v(20[7:21])
    defparam i4326_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4560));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4559));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(deadband[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4610));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4558));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4557));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[0]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4555));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[1]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4553));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[2]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4551));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4550));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(deadband[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4609));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4548));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4547));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(deadband[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4619));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4546));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4545));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49161_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(PWMLimit[9]), 
            .I3(n356[9]), .O(n66177));
    defparam i49161_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4544));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4543));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[3]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4541));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[4]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4539));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[5]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4537));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[6]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4535));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[7]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[8]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[9]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[10]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[11]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[12]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[13]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[14]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[15]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4522));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4521));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35189_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I2(\PID_CONTROLLER.integral_23__N_3715 [21]), .I3(\Ki[1] ), 
            .O(n20600[0]));   // verilog/motorControl.v(50[27:38])
    defparam i35189_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[16]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35191_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I2(\PID_CONTROLLER.integral_23__N_3715 [21]), .I3(\Ki[1] ), 
            .O(n50810));   // verilog/motorControl.v(50[27:38])
    defparam i35191_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(deadband[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4605));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4519));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[17]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4517));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4516));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[18]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35347_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I2(n4_adj_4951), .I3(n20536[1]), .O(n6_adj_4952));   // verilog/motorControl.v(50[27:38])
    defparam i35347_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_956 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I2(n4_adj_4951), .I3(n20536[1]), .O(n20476[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_956.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4514));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_957 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I2(n50958), .I3(n20536[0]), .O(n20476[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_957.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[19]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4512));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[20]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4510));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35339_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I2(n50958), .I3(n20536[0]), .O(n4_adj_4951));   // verilog/motorControl.v(50[27:38])
    defparam i35339_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4509));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35326_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3715 [18]), .I3(\Ki[1] ), 
            .O(n20476[0]));   // verilog/motorControl.v(50[27:38])
    defparam i35326_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i35328_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3715 [18]), .I3(\Ki[1] ), 
            .O(n50958));   // verilog/motorControl.v(50[27:38])
    defparam i35328_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4508));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4507));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4506));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[21]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4504));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4503));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4502));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_958 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(n4_adj_4953), .I3(n20576[1]), .O(n20536[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_958.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[22]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35309_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(n4_adj_4953), .I3(n20576[1]), .O(n6_adj_4954));   // verilog/motorControl.v(50[27:38])
    defparam i35309_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4500));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4499));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35301_3_lut_4_lut (.I0(n62_adj_4955), .I1(n131_adj_4956), .I2(n204_adj_4957), 
            .I3(n20576[0]), .O(n4_adj_4953));   // verilog/motorControl.v(50[27:38])
    defparam i35301_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4982[23]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_adj_959 (.I0(n62_adj_4955), .I1(n131_adj_4956), 
            .I2(n204_adj_4957), .I3(n20576[0]), .O(n20536[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_959.LUT_INIT = 16'h8778;
    SB_LUT4 i35252_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3715 [20]), .I3(\Ki[1] ), 
            .O(n50876));   // verilog/motorControl.v(50[27:38])
    defparam i35252_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4496));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35250_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3715 [20]), .I3(\Ki[1] ), 
            .O(n20576[0]));   // verilog/motorControl.v(50[27:38])
    defparam i35250_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4495));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4494));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4493));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4492));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18139_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25));   // verilog/motorControl.v(41[14] 61[8])
    defparam i18139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23670_1_lut (.I0(n356[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n39319));   // verilog/motorControl.v(50[18:38])
    defparam i23670_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[0]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n49[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49189_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(PWMLimit[7]), 
            .I3(n356[7]), .O(n66205));
    defparam i49189_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4490));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n49[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4488));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_960 (.I0(n20536[2]), .I1(n6_adj_4952), .I2(\Ki[4] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715 [18]), .O(n20476[3]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_960.LUT_INIT = 16'h9666;
    SB_LUT4 mult_17_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_4957));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_961 (.I0(n20600[0]), .I1(n50876), .I2(\Ki[2] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715 [20]), .O(n20576[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_961.LUT_INIT = 16'h9666;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_4956));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_4955));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n207[19]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i20_3_lut (.I0(n207[19]), .I1(IntegralLimit[19]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [19]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n207[18]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i19_3_lut (.I0(n207[18]), .I1(IntegralLimit[18]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [18]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_962 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3715 [23]), .O(n62030));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_962.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_963 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(\PID_CONTROLLER.integral_23__N_3715 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3715 [19]), .O(n62034));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_963.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_964 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I3(\PID_CONTROLLER.integral_23__N_3715 [21]), .O(n62032));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_964.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_965 (.I0(n62032), .I1(n50810), .I2(n62034), .I3(n62030), 
            .O(n62040));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i35263_4_lut (.I0(n20600[0]), .I1(\Ki[2] ), .I2(n50876), .I3(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .O(n4_adj_4960));   // verilog/motorControl.v(50[27:38])
    defparam i35263_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i35355_4_lut (.I0(n20536[2]), .I1(\Ki[4] ), .I2(n6_adj_4952), 
            .I3(\PID_CONTROLLER.integral_23__N_3715 [18]), .O(n8_adj_4961));   // verilog/motorControl.v(50[27:38])
    defparam i35355_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_966 (.I0(n6_adj_4954), .I1(n8_adj_4961), .I2(n4_adj_4960), 
            .I3(n62040), .O(n60196));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n49[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4598));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4487));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n49[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n363), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4567));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4962));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4486));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4963));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49157_3_lut_4_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(n356[2]), .O(n66173));   // verilog/motorControl.v(54[23:39])
    defparam i49157_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(GND_net), .O(n6_adj_4945));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[1]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4484));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4483));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[2]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4481));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[3]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4479));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[4]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4477));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4476));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n207[17]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i18_3_lut (.I0(n207[17]), .I1(IntegralLimit[17]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [17]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[5]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4474));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[6]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4472));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4471));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[7]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n49[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4964));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4965));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[8]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[9]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4966));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4967));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4968));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4969));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4970));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48971_4_lut (.I0(n21_adj_4711), .I1(n19_adj_4712), .I2(n17_adj_4714), 
            .I3(n9_adj_4706), .O(n65987));
    defparam i48971_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n306[0]));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n49[0]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[10]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n49[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[11]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48948_4_lut (.I0(n27_adj_4719), .I1(n15_adj_4709), .I2(n13_adj_4708), 
            .I3(n11_adj_4707), .O(n65964));
    defparam i48948_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[12]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[13]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n49[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4463));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[14]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4461));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[15]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[16]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[17]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[18]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[19]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[20]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155_adj_4607), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4453));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4452));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[21]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4450));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[22]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4981[23]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4446));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4445));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[0]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4443));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4442));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_4969), 
            .I3(GND_net), .O(n12_adj_4972));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_4708), 
            .I3(GND_net), .O(n10_adj_4973));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[1]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4441));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4440));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[2]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4438));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4437));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[3]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4435));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[4]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4434));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[5]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4433));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[6]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48584_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n65600));
    defparam i48584_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4432));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[7]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4431));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n49[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[8]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[9]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48631_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n65647));
    defparam i48631_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[10]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[11]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_4972), .I1(n130[17]), .I2(n35_adj_4970), 
            .I3(GND_net), .O(n30_adj_4974));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48898_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n65914));   // verilog/motorControl.v(47[21:44])
    defparam i48898_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_adj_4667));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49410_2_lut_4_lut (.I0(deadband[21]), .I1(n356[21]), .I2(deadband[9]), 
            .I3(n356[9]), .O(n66426));
    defparam i49410_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49017_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n66033));   // verilog/motorControl.v(45[12:34])
    defparam i49017_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[12]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_4975));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[13]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[14]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48582_3_lut_4_lut (.I0(deadband[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(deadband[2]), .O(n65598));   // verilog/motorControl.v(51[12:29])
    defparam i48582_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_4616));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49910_4_lut (.I0(n13_adj_4708), .I1(n11_adj_4707), .I2(n9_adj_4706), 
            .I3(n66033), .O(n66926));
    defparam i49910_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[15]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[16]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n49[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[17]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4980[18]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49243_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(PWMLimit[2]), .O(n66259));   // verilog/motorControl.v(52[14:29])
    defparam i49243_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_4844));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49902_4_lut (.I0(n19_adj_4712), .I1(n17_adj_4714), .I2(n15_adj_4709), 
            .I3(n66926), .O(n66918));
    defparam i49902_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35423_2_lut_4_lut (.I0(\Kp[0] ), .I1(n49[20]), .I2(\Kp[1] ), 
            .I3(n49[19]), .O(n20560[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35423_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i51034_4_lut (.I0(n25_adj_4717), .I1(n23_adj_4716), .I2(n21_adj_4711), 
            .I3(n66918), .O(n68050));
    defparam i51034_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4597));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50399_4_lut (.I0(n31_adj_4968), .I1(n29_adj_4967), .I2(n27_adj_4719), 
            .I3(n68050), .O(n67415));
    defparam i50399_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n49[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4596));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51183_4_lut (.I0(n37_adj_4965), .I1(n35_adj_4970), .I2(n33_adj_4969), 
            .I3(n67415), .O(n68199));
    defparam i51183_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43_adj_4963), 
            .I3(GND_net), .O(n16_adj_4976));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49428_2_lut_4_lut (.I0(deadband[16]), .I1(n356[16]), .I2(deadband[7]), 
            .I3(n356[7]), .O(n66444));
    defparam i49428_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50425_3_lut (.I0(n6_adj_4975), .I1(n130[10]), .I2(n21_adj_4711), 
            .I3(GND_net), .O(n67441));   // verilog/motorControl.v(45[12:34])
    defparam i50425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50426_3_lut (.I0(n67441), .I1(n130[11]), .I2(n23_adj_4716), 
            .I3(GND_net), .O(n67442));   // verilog/motorControl.v(45[12:34])
    defparam i50426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_4714), 
            .I3(GND_net), .O(n8_adj_4977));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_4976), .I1(n130[22]), .I2(n45_adj_4966), 
            .I3(GND_net), .O(n24_adj_4978));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48902_4_lut (.I0(n43_adj_4963), .I1(n25_adj_4717), .I2(n23_adj_4716), 
            .I3(n65987), .O(n65918));
    defparam i48902_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50636_4_lut (.I0(n24_adj_4978), .I1(n8_adj_4977), .I2(n45_adj_4966), 
            .I3(n65916), .O(n67652));   // verilog/motorControl.v(45[12:34])
    defparam i50636_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49610_3_lut (.I0(n67442), .I1(n130[12]), .I2(n25_adj_4717), 
            .I3(GND_net), .O(n66626));   // verilog/motorControl.v(45[12:34])
    defparam i49610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4979));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i50423_3_lut (.I0(n4_adj_4979), .I1(n130[13]), .I2(n27_adj_4719), 
            .I3(GND_net), .O(n67439));   // verilog/motorControl.v(45[12:34])
    defparam i50423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4595));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50424_3_lut (.I0(n67439), .I1(n130[14]), .I2(n29_adj_4967), 
            .I3(GND_net), .O(n67440));   // verilog/motorControl.v(45[12:34])
    defparam i50424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n49[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4594));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48938_4_lut (.I0(n33_adj_4969), .I1(n31_adj_4968), .I2(n29_adj_4967), 
            .I3(n65964), .O(n65954));
    defparam i48938_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51012_4_lut (.I0(n30_adj_4974), .I1(n10_adj_4973), .I2(n35_adj_4970), 
            .I3(n65950), .O(n68028));   // verilog/motorControl.v(45[12:34])
    defparam i51012_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49612_3_lut (.I0(n67440), .I1(n130[15]), .I2(n31_adj_4968), 
            .I3(GND_net), .O(n66628));   // verilog/motorControl.v(45[12:34])
    defparam i49612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51254_4_lut (.I0(n66628), .I1(n68028), .I2(n35_adj_4970), 
            .I3(n65954), .O(n68270));   // verilog/motorControl.v(45[12:34])
    defparam i51254_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51255_3_lut (.I0(n68270), .I1(n130[18]), .I2(n37_adj_4965), 
            .I3(GND_net), .O(n68271));   // verilog/motorControl.v(45[12:34])
    defparam i51255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51188_3_lut (.I0(n68271), .I1(n130[19]), .I2(n39_adj_4964), 
            .I3(GND_net), .O(n68204));   // verilog/motorControl.v(45[12:34])
    defparam i51188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48911_4_lut (.I0(n43_adj_4963), .I1(n41_adj_4962), .I2(n39_adj_4964), 
            .I3(n68199), .O(n65927));
    defparam i48911_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50941_4_lut (.I0(n66626), .I1(n67652), .I2(n45_adj_4966), 
            .I3(n65918), .O(n67957));   // verilog/motorControl.v(45[12:34])
    defparam i50941_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49618_3_lut (.I0(n68204), .I1(n130[20]), .I2(n41_adj_4962), 
            .I3(GND_net), .O(n66634));   // verilog/motorControl.v(45[12:34])
    defparam i49618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51120_4_lut (.I0(n66634), .I1(n67957), .I2(n45_adj_4966), 
            .I3(n65927), .O(n68136));   // verilog/motorControl.v(45[12:34])
    defparam i51120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50837_3_lut (.I0(n4_adj_4678), .I1(n356[13]), .I2(n27), .I3(GND_net), 
            .O(n67853));   // verilog/motorControl.v(51[12:29])
    defparam i50837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51121_3_lut (.I0(n68136), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155_adj_4607));   // verilog/motorControl.v(45[12:34])
    defparam i51121_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
