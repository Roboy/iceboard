// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu May 21 15:11:04 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    
    wire n36823;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n60331;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(351[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(359[15:20])
    
    wire pwm_setpoint_23__N_207, n12187, n12191, n6, n260, n12227, 
        n294, n298, n299, n300, n301, n302, n303, n304, n305, 
        n306, n307, n308, n309, n49650, n49763, n49649, n49762, 
        n15, n4928, n4927, n4926, n4925, n4924, n4923, n4922, 
        n4921, n4920, n4919, n4918, n4917, n4916, n59279;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n49761;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n61974, GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, 
        GLC_N_400, dti_N_404, n29999, RX_N_2, n66402, n1744, n1742;
    wire [31:0]motor_state_23__N_91;
    wire [32:0]encoder0_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        read_N_409, n1319, n61968, n49648, n49647, n68547, n49760, 
        n49646, n7, n6_adj_5676, n5, n4, n26, n19, n17, n16, 
        n15_adj_5677, n13, n11, n9, n8, n7_adj_5678, n6_adj_5679, 
        n5_adj_5680, n4_adj_5681, n1784, n1786, n1788, n1790, n1792, 
        n1794, n1796;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n1822, n1824;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [1:0]state;   // verilog/neopixel.v(16[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    
    wire n68473, n69135, n49759, n4915, n4914, n4913, n4912, n4911, 
        n4910, n61964, n625, n43396, n4940, n4937, n29989, n49903, 
        n49534, n69679, n61958, n49902, n29986, n29983, n61956, 
        n59130, n623;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n9_adj_5682, n25, n24, n8_adj_5683, n23, n22, n21, n20, 
        n49901, n26_adj_5684, n19_adj_5685, n17_adj_5686, n16_adj_5687, 
        n61954, n49758, n49757, n622, n621, n2, n14, n15_adj_5688, 
        n16_adj_5689, n17_adj_5690, n18, n19_adj_5691, n20_adj_5692, 
        n21_adj_5693, n22_adj_5694, n23_adj_5695, n24_adj_5696, n25_adj_5697, 
        n68384, n5774, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    
    wire n49756, n49755;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active, n68360, n68359, n49900, n49754;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n49899, n3470, n2820, n49898, 
        n29979, n49897, n49896, n25465, n2873, n49895, n25595, 
        n161, n49753, n68471, n68313, n4909, n4908, n4907, n15_adj_5698, 
        n29976, n49533, n49752, n49751, n49894, n6_adj_5699, n49645, 
        n49644, n49643, n49750, n61932, n49642, n49749, n50523, 
        n49641, n49640, n4_adj_5700, n68240, n49518, n49748, n49639, 
        n49638, n50522, n50521, n50520, n49747, n49746, n50519, 
        n49637, n50518, n50517, n49636, n50516, n49745, n49744, 
        n50515, n49532, n50514, n50513, n50512, n50511, n50510, 
        n50509, n49880, n49879, n50508, n50507, n50107, n50506, 
        n50505, n50504, n50106, n49531, n50503, n49878, n50502, 
        n49635, n49877, n49876, n50501, n50105, n50104, n49875, 
        n50500, n50499, n49874, n50103, n50102, n49873, n50498, 
        n50497, n50496, n49530, n50495, n50101, n50494, n50493, 
        n50100, n49872, n50492, n50491, n50490, n50489, n50099, 
        n50488, n50487, n50486, n50485, n49634, n50098, n50484, 
        n50097, n50483, n50482, n50096, n49633, n50481, n61926, 
        n50095, n50480, n50479, n50094, n50093, n50478, n50477, 
        n61924, n50476, n50475, n50474, n50092, n50473, n50472, 
        n50471, n50470, n50469, n49529, n49632, n50468, n50467, 
        n42792, n50466, n50465, n42845, n50464, n50463, n50462, 
        n50461, n61918, n50460, n61916, n50459, n61914, n50458, 
        n50457, n49517, n49631, n50456, n50455, n50454, n42890, 
        n50453, n42880, n68167, n68386, n68388, n68068, n61902, 
        n68067, n69673, n69667, n15_adj_5701, n11_adj_5702, n61896, 
        n25505, n25848, n67264, n61886, n12225, n32, n31, n50452, 
        n50451, n13_adj_5703, n67858, n67210, n61880, n61874, n62220, 
        n61864, n6_adj_5704, n61860, Kp_23__N_1389, n61854, n61852, 
        n43717, n30, n29, n28, n12189, n27, n26_adj_5705, n25_adj_5706, 
        n24_adj_5707, n23_adj_5708, n22_adj_5709, n21_adj_5710, n20_adj_5711, 
        n19_adj_5712, n18_adj_5713, n17_adj_5714, n16_adj_5715, n15_adj_5716, 
        n14_adj_5717, n13_adj_5718, n12, n11_adj_5719, n10, n9_adj_5720, 
        n8_adj_5721, n7_adj_5722, n6_adj_5723, \FRAME_MATCHER.i_31__N_2513 , 
        Kp_23__N_1748, n5_adj_5724, n50450, n43575, n43567, n67280, 
        n61836, n29912, n29900, n29879, n29878, n29877, n29876, 
        n29875, n29874, n29873, n29872, n29871, n29870, n29869, 
        n29868, n29867, n29866, n29865, n29864, n29863, n29862, 
        n29861, n29860, n29859, n29858, n29857, n29856, n29855, 
        n29854, n29853, n29852, n29851, n29850, n29849, n29848, 
        n29847, n29846, n29845, n29844, n29843, n29842, n29841, 
        n29840, n29839, n29838, n29837, n29836, n29835, n29834, 
        n29833, n29832, n29831, n29830, n29829, n29827, n29826, 
        n29825, n29824, n29823, n29822, n29821, n29820, n29819, 
        n29818, n29817, n29816, n29815, n29814, n29813, n29812, 
        n29811, n29810, n29809, n29808, n29807, n29805, n29802, 
        n29798, n29797, n29796, n43615, n43613, n43611, n43511, 
        n29767, n43605, n29764, n29760, n29759, n36852, n5_adj_5725, 
        n524, n523, n522, n521, n29758, n29757, n29756, n29755, 
        n29754, n29753, n29752, n29751, n29750, n29749, n29748, 
        n29747, n29746, n29745, n29744, n29743, n29742, n29739, 
        n29738, n29735, n29734, n29733, n29732, n29731, n29730, 
        n29729, n29725, n29721, n29718, n58170, n29714, n29707, 
        n29701, n29700, n29699, n29692, n29691, n29690, n43595, 
        n29683, n29677, n29676, n29675, n29673, n29672, n29671, 
        n29669, n43591, n29664, n29663, n29662, n29661, n29660, 
        n43589, n29656, n29655, n29654, n29653, n29652, n43587, 
        n43585, n29645, n29644, n43583, n29637, n29636, n29635, 
        n29632, n29628, n29624, n29621, n29618, n29609, n56536, 
        n56538, n56540, n29594, n56542, n53095, n29576, n29573, 
        n29570, n61830, n30_adj_5726, n68061, n23_adj_5727, n21_adj_5728, 
        n19_adj_5729, n59015, n520, n4_adj_5730, n3, n2_adj_5731, 
        n17_adj_5732, n16_adj_5733, n15_adj_5734, n13_adj_5735, n11_adj_5736, 
        n10_adj_5737, n9_adj_5738, n8_adj_5739, n7_adj_5740, n6_adj_5741, 
        n4_adj_5742, n25615, n69088, n61824, n61822, n67855, n67934, 
        n15_adj_5743, n58373, n7_adj_5744, n4_adj_5745, n4_adj_5746, 
        n67854, n59026, n50072, n10_adj_5747, n6_adj_5748, n50995, 
        n30549, n30548, n30547, n30546, n30545, n30544, n30543, 
        n519, n518, n516, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    
    wire n50071, n30538, n50994, n50993, n30534, n30533, n30529, 
        n155, n212, n213, n214, n219;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3715 ;
    
    wire n365, n379, n380, n405, n69661, n459, n460, n12185, 
        n61804, n30523, n30519, n43621, n30512, n26517, n43619, 
        n30506, n6_adj_5749, n30504, n30503, n50992, n30501, n30500, 
        n30499, n30498, n30497, n30496, n30495, n15_adj_5750, n11_adj_5751, 
        n30494, n30493, n30491;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, n30490, n30489, n30488, n50991, n30487, position_31__N_3827, 
        n50449, n50070, n30486, n30485, n30484, n30483, n30482, 
        n30481, n30480, n30479, n30478, n30477, n30476, n30475, 
        n30474, n30473, n50069, n50448, n50990;
    wire [1:0]a_new_adj_5965;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5753, n50447, position_31__N_3827_adj_5754, n61800, 
        n50068, n61798, n50446, n50989, n49630, n50445, n50067, 
        n50444;
    wire [7:0]data_adj_5978;   // verilog/eeprom.v(23[12:16])
    
    wire ready_prev, rw;
    wire [7:0]state_adj_5979;   // verilog/eeprom.v(27[11:16])
    
    wire n50066;
    wire [7:0]state_7__N_3916;
    
    wire n50443, n8_adj_5757, n30440, n61792, n30439, n30438, n30437, 
        n30436, n30435, n61788, n30434, n50065, n30433, n50064, 
        n50988, n50063, n30432, n30431, n30429, n30428, n30427, 
        n50442, n30426, n6617, n30425, n30424, n30423, n50441, 
        n58317, n30422, n30421, n30420, n30419, n30418, n50987, 
        n30417, n30415, n25477, n4906, n4905, n49528, n50440, 
        clk_out;
    wire [15:0]data_adj_5985;   // verilog/tli4970.v(27[14:18])
    
    wire n50986, n50439, n50438;
    wire [7:0]state_adj_5987;   // verilog/tli4970.v(29[13:18])
    
    wire n19_adj_5768, n18_adj_5769, n17_adj_5770, n4_adj_5771, n3_adj_5772, 
        n2_adj_5773, n58304, n50437, n50985, n50436, n30383, n30382, 
        n50435, n30381, n60222, n30380, n30378, n30372, n30371, 
        n50984, n50983, n50434, n30355, n30354, n50982, n50062, 
        n50981, n50433, n50432, n30353, n30352, n30351, n30350, 
        n30349, n30348, n30347, n12193, n12195, n12197, n12199, 
        n8_adj_5774, state_7__N_4317, n50431, n50430, n58294, n30343, 
        n30342, n16_adj_5775, n30336, n8_adj_5776, n58292, n50429, 
        n50980, n30317, n50061, n50979, n50978, n50977, n50976, 
        n30316, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n50975, n30314, n22917, n50974, n12201, n12203, n12205, 
        n12207, n12209, n12211, n12213, n12215, n50060, n50973, 
        n69640, n69637;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n12217, n12219, n12221, n12223, n29536, n15_adj_5777, n14_adj_5778, 
        n13_adj_5779, n12_adj_5780, n61768;
    wire [2:0]r_SM_Main_adj_5996;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5997;   // verilog/uart_tx.v(33[16:29])
    
    wire n50428, n30287, n58290, n50972, n50059, n50971, n50427, 
        n50970, n11_adj_5791, n10_adj_5792, n9_adj_5793, n50426, n8_adj_5794, 
        n7_adj_5795, n6_adj_5796, n30265, n43537;
    wire [7:0]state_adj_6010;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n61764, enable_slow_N_4211, n5_adj_5798, n50425, n66334, 
        n5_adj_5799, n36888, n50058, n49853;
    wire [7:0]state_7__N_4108;
    
    wire n50424, n50423, n6428, n3_adj_5800, n50422;
    wire [7:0]state_7__N_4124;
    
    wire n50969, n50968, n61762, n50421, n30251, n30246, n30245, 
        n30244, n30243, n30242, n8_adj_5801, n30241, n50967, n30240, 
        n58278, n29530, n50420, n30231, n30230, n29526, n29523, 
        n29520, n56568, n50419, n43541, n50966, n50418, n50417, 
        n61758, n49629, n50416, n50415, n50965, n50414, n49628, 
        n50413, n7455, n7454, n7453, n7452, n7451, n7450, n50412, 
        n828, n829, n830, n831, n832, n833, n861, n50411, n896, 
        n897, n898, n899, n900, n901, n927, n928, n929, n930, 
        n931, n932, n933, n939, n940, n941, n942, n943, n944, 
        n945, n946, n947, n948, n949, n950, n951, n952, n953, 
        n954, n955, n956, n957, n960, n995, n996, n997, n998, 
        n999, n1000, n1001, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n42305, n42304, n1059, n1093, n1094, 
        n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1125, 
        n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
        n1158, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
        n1200, n1201, n50410, n1224_adj_5802, n1225_adj_5803, n1226_adj_5804, 
        n1227_adj_5805, n1228_adj_5806, n1229_adj_5807, n1230_adj_5808, 
        n1231_adj_5809, n1232_adj_5810, n1233_adj_5811, n61746, n25_adj_5812, 
        n1257, n50409, n1291, n1292, n1293, n1294, n1295, n1296, 
        n1297, n1298, n1299, n1300, n1301, n50408, n50407, n1323, 
        n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
        n1332, n1333, n1356, n1391, n1392, n1393, n1394, n1395, 
        n1396, n1397, n1398, n1399, n1400, n1401, n50406, n50405, 
        n50404, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
        n1429, n1430, n1431, n1432, n1433, n1455, n490, n61740, 
        n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
        n1498, n1499, n1500, n1501, n1521, n1522, n1523, n1524, 
        n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
        n1533, n41755, n41756, n1554, n69063, n1589, n1590, n1591, 
        n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
        n1600, n1601, n1620, n1621, n1622, n1623, n1624, n1625, 
        n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
        n68592, n1653, n50403, n1687, n1688, n1689, n1690, n1691, 
        n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
        n1700, n1701, n61726, n1719, n1720, n1721, n1722, n1723, 
        n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
        n1732, n1733, n1752, n50402, n61720, n1787, n1788_adj_5813, 
        n1789, n1790_adj_5814, n1791, n1792_adj_5815, n1793, n1794_adj_5816, 
        n1795, n1796_adj_5817, n1797, n1798, n1799, n1800, n1801, 
        n1818, n1819, n1820, n1821, n1822_adj_5818, n1823, n1824_adj_5819, 
        n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
        n1833, n19_adj_5820, n1851, n20_adj_5821, n1885, n1886, 
        n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
        n1895, n1896, n1897, n1898, n1899, n1900, n1901, n61714, 
        n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
        n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
        n1933, n69092, n1950, n1985, n1986, n1987, n1988, n1989, 
        n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
        n1998, n1999, n2000, n2001, n2016, n2017, n2018, n2019, 
        n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
        n2028, n2029, n2030, n2031, n2032, n2033, n2049, n2084, 
        n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
        n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
        n2101, n2115, n2116, n2117, n2118, n2119, n2120, n2121, 
        n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
        n2130, n2131, n2132, n2133, n2148, n2182, n2183, n2184, 
        n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
        n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
        n2201, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
        n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
        n2229, n2230, n2231, n2232, n2233, n66937, n41114, n2247, 
        n31_adj_5822, n2282, n2283, n2284, n2285, n2286, n2287, 
        n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
        n2296, n2297, n2298, n2299, n2300, n2301, n2313, n2314, 
        n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
        n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
        n2331, n2332, n2333, n2346, n2381, n2382, n2383, n2384, 
        n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
        n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
        n2401, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
        n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
        n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2445, 
        n172, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
        n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
        n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2511, 
        n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
        n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, 
        n2528, n2529, n2530, n2531, n2532, n2533, n2544, n61700, 
        n417, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
        n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
        n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
        n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, 
        n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
        n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
        n2643, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
        n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
        n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
        n2701, n2709, n2710, n2711, n2712, n2713, n2714, n2715, 
        n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
        n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, 
        n2732, n2733, n2742, n57410, n106, n105, n58179, n91, 
        n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
        n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
        n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
        n2800, n2801, n2808, n2809, n2810, n2811, n2812, n2813, 
        n2814, n2815, n2816, n2817, n2818, n2819, n2820_adj_5823, 
        n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
        n2829, n2830, n2831, n2832, n2833, n2841, n58177, n61696, 
        n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
        n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
        n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
        n2900, n2901, n2907, n2908, n2909, n2910, n2911, n2912, 
        n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
        n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
        n2929, n2930, n2931, n2932, n2933, n2940, n58175, n2975, 
        n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
        n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
        n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
        n3000, n3001, n3006, n3007, n3008, n3009, n3010, n3011, 
        n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
        n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
        n3028, n3029, n3030, n3031, n3032, n3033, n68813, n3039, 
        n50401, n58173, n50400, n20203, n50399, n3074, n3075, 
        n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
        n3100, n3101, n3105, n3106, n3107, n3108, n3109, n3110, 
        n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
        n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
        n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3138, 
        n50398, n58169, n50397, n3173, n3174, n3175, n3176, n3177, 
        n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
        n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
        n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
        n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
        n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
        n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
        n3228, n3229, n3230, n3231, n3232, n3233, n50396, n3237, 
        n50395, n42725, n3272, n3273, n3274, n3275, n3276, n3277, 
        n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, 
        n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
        n3294, n3295, n3296, n3298, n3301, n68744, n61688, n50394, 
        n50393, n24_adj_5824, n50392, n27_adj_5825, n50391, n50390, 
        n50389, n50388, n50387, n62, n50386, n61680, n50385, n25480, 
        n50384, n28027, n50383, n27996, n50382, n49852, n61670, 
        n43, n45, n61664, n50381, n43398, n53024, n57879, n61658, 
        n50380, n50379, n27950, n43400, n30203, n50378, n30199, 
        n30196, n50377, n49851, n50376, n50375, n49516, n67947, 
        n50374, n30186, n50373, n49850, n61652, n25471, n61650, 
        n30183, n61648, n50372, n50371, n30180, n49849, n30177, 
        n27810, n30176, n61644, n49848, n30173, n50370, n59100, 
        n50369, n50030, n30170, n50368, n50367, n61980, n30167, 
        n27754, n25593, n50366, n49847, n56774, n27736, n50365, 
        n25590, n69775, n69769, n69034, n61634, n4_adj_5826, n69763, 
        n4_adj_5827, n30_adj_5828, n32_adj_5829, n4_adj_5830, n69757, 
        n69378, n27728, n27726, n27722, n50029, n50364, n50363, 
        n50028, n50362, n50361, n67946, n50360, n344, n20252, 
        n68593, n61628, n50359, n50358, n61622, n20204, n50357, 
        n50356, n20205, n61616, n50355, n50354, n61614, n20253, 
        n271, n50353, n50027, n49846, n50352, n27676, n50351, 
        n25612, n30154, n50026, n50350, n61608, n50025, n68060, 
        n61602, n50349, n50024, n56570, n198, n50348, n61596, 
        n30151, n50023, n50347, n50346, n61590, n27652, n50345, 
        n50344, n61582, n30148, n61580, n125, n50022, n50343, 
        n61576, n50342, n50341, n61568, n43_adj_5831, n69365, n37308, 
        n61566, n50340, n50339, n110, n61564, n35, n61562, n61560, 
        n38, n61558, n50338, n50021, n50337, n50336, n61556, n4_adj_5832, 
        n56, n53, n61554, n61552, n50335, n50020, n50019, n50018, 
        n50334, n61550, n50333, n61548, n61546, n50017, n61544, 
        n50332, n50331, n61542, n61538, n50330, n61530, n50329, 
        n50328, n61528, n61526, n57819, n50327, n50326, n61524, 
        n50325, n61518, n50324, n50323, n61512, n50322, n61506, 
        n61504, n50321, n50320, n61498, n61496, n50319, n50318, 
        n50317, n66774, n50316, n61484, n66772, n61478, n59370, 
        n50315, n50314, n66764, n61472, n66748, n61466, n49999, 
        n61460, n4_adj_5833, n6_adj_5834, n8_adj_5835, n9_adj_5836, 
        n50313, n4_adj_5837, n6_adj_5838, n8_adj_5839, n9_adj_5840, 
        n11_adj_5841, n13_adj_5842, n15_adj_5843, n69350, n61454, 
        n61452, n49998, n50312, n50311, n50310, n49997, n50309, 
        n59115, n50308, n50307, n50306, n50305, n49996, n50304, 
        n49995, n50303, n50302, n50301, n50300, n50299, n38_adj_5844, 
        n39, n40, n41, n42, n43_adj_5845, n44, n45_adj_5846, n29510, 
        n29508, n11610, n69751, n11579, n11577, n49834, n49833, 
        n50298, n50297, n57392, n61440, n60332, n53127, n43450, 
        n53215, n29192, n61434, n61428, n68809, n57425, n28464, 
        n57426, n61424, n28915, n28908, n28413, n28409, n57317, 
        n49994, n50296, n50295, n49993, n49992, n49991, n49832, 
        n50294, n50767, n50766, n61414, n60225, n50293, n50765, 
        n50292, n50764, n66607, n49831, n50763, n49990, n50762, 
        n69006, n50761, n49989, n50291, n49830, n50290, n50289, 
        n61412, n49988, n49829, n49828, n49987, n50288, n38_adj_5847, 
        n35_adj_5848, n61406, n34, n33, n56546, n32_adj_5849, n50287, 
        n31_adj_5850, n22792, n50286, n61400, n30144, n30141, n61396, 
        n4_adj_5851, n50285, n50284, n61390, n50283, n62096, n68059, 
        n61382, n66552, n50282, n50281, n49527, n50280, n50279, 
        n30138, n6_adj_5852, n30134, n30131, n30125, n30122, n30118, 
        n30115, n30112, n30108, n50278, n66548, n50277, n50276, 
        n61376, n21_adj_5853, n30105, n59018, n30102, n30099, n30096, 
        n30093, n43687, n30087, n43685, n30083, n30080, n30077, 
        n49822, n49821, n68740, n50275, n49820, n50274, n30068, 
        n43677, n30065, n30062, n25578, n30059, n50273, n61370, 
        n43671, n30055, n43669, n49819, n29477, n43667, n5_adj_5854, 
        n43663, n53678, n49818, n50272, n43655, n43651, n50271, 
        n50270, n50269, n49817, n50268, n50267, n50266, n50265, 
        n49816, n49815, n50264, n50263, n50262, n49814, n49813, 
        n50261, n49812, n50260, n57737, n50259, n49962, n49961, 
        n50258, n50257, n50256, n49960, n50255, n49959, n50254, 
        n50253, n50252, n49958, n50251, n49957, n2_adj_5855, n3_adj_5856, 
        n4_adj_5857, n5_adj_5858, n6_adj_5859, n7_adj_5860, n8_adj_5861, 
        n9_adj_5862, n10_adj_5863, n11_adj_5864, n12_adj_5865, n13_adj_5866, 
        n14_adj_5867, n15_adj_5868, n16_adj_5869, n17_adj_5870, n18_adj_5871, 
        n19_adj_5872, n20_adj_5873, n21_adj_5874, n22_adj_5875, n23_adj_5876, 
        n24_adj_5877, n25_adj_5878, n26_adj_5879, n27_adj_5880, n28_adj_5881, 
        n29_adj_5882, n30_adj_5883, n31_adj_5884, n32_adj_5885, n49420, 
        n50250, n50249, n49526, n50248, n50247, n49525, n50246, 
        n66520, n49515, n50245, n49956, n49955, n50244, n50243, 
        n50242, n50241, n50240, n50239, n50238, n50237, n49954, 
        n49953, n50236, n49952, n49951, n50235, n50234, n50233, 
        n50232, n50231, n50230, n50229, n50228, n50227, n50226, 
        n49514, n50225, n50224, n50223, n50222, n49524, n50221, 
        n50220, n50219, n50218, n50217, n50216, n50215, n50214, 
        n50213, n66510, n49523, n50212, n50211, n50210, n50209, 
        n50208, n50207, n50206, n50205, n66508, n50204, n50203, 
        n50202, n50201, n50200, n50199, n50198, n50197, n50196, 
        n50195, n50194, n50193, n50192, n50191, n50190, n50189, 
        n50188, n69333, n49513, n49522, n49512, n49935, n49934, 
        n49521, n49933, n49520, n62794, n49932, n49931, n49930, 
        n49929, n49928, n49927, n49926, n49779, n62090, n49925, 
        n66483, n49778, n49777, n49776, n49775, n49774, n49773, 
        n66470, n49772, n111, n49519, n49771, n49511, n49770, 
        n49541, n49769, n50165, n49768, n49767, n49540, n50164, 
        n49539, n50163, n49538, n50162, n49537, n49536, n13_adj_5886, 
        n15_adj_5887, n19_adj_5888, n23_adj_5889, n27_adj_5890, n31_adj_5891, 
        n59, n61, n50161, n49766, n49470, n50160, n33793, n25600, 
        n50159, n20969, n33801, n49765, n20965, n49764, n20283, 
        n62084, n63007, n62082, n57685, n29471, n29474, n69745, 
        n62076, n62072, n62070, n62068, n69303, n59056, n52186, 
        n11642, n10_adj_5892, n25564, n50158, n50157, n50156, n50155, 
        n50154, n68974, n50153, n50152, n53222, n69691, n50151, 
        n63154, n52054, n57336, n50150, n69739, n50149, n25587, 
        n69297, n49535, n25583, n52011, n62060, n6_adj_5893, n68948, 
        n69733, n62046, n61170, n6_adj_5894, n62040, n61154, n65782, 
        n65775, n61138, n69727, n5_adj_5895, n61122, n55644, n24_adj_5896, 
        n17_adj_5897, n25_adj_5898, n68081, n61106, n69225, n65740, 
        n65737, n67758, n55740, n61090, n61074, n68521, n61058, 
        n58171, n67766, n57499, n4_adj_5899, n67774, n57625, n12_adj_5900, 
        n69721, n57657, n69206, n4_adj_5901, n5_adj_5902, n67324, 
        n57990, n58117, n57956, n63008, n6_adj_5903, n68915, n14_adj_5904, 
        n10_adj_5905, n59034, n60151, n25_adj_5906, n15_adj_5907, 
        n14_adj_5908, n58132, n14_adj_5909, n13_adj_5910, n22_adj_5911, 
        n69715, n57862, n6_adj_5912, n62574, n62578, n62582, n69184, 
        n62792, n62790, n4_adj_5913, n67358, n69974, n59013, n60224, 
        n56368, n56398, n56402, n56406, n56410, n8_adj_5914, n56414, 
        n7_adj_5915, n56418, n56422, n59080, n56430, n56434, n56438, 
        n56442, n56446, n56450, n57340, n56454, n56458, n56462, 
        n57836, n56466, n56470, n56474, n56478, n9_adj_5916, n7_adj_5917, 
        n65611, n56534, n59684, n57437, n8_adj_5918, n56566, n12_adj_5919, 
        n56604, n65589, n65588, n56636, n69709, n56662, n7_adj_5920, 
        n65579, n65578, n56678, n69160, n63155, n56690, n57424, 
        n62647, n7_adj_5921, n62929, n62927, n62926, n62923, n69703, 
        n23_adj_5922, n6_adj_5923, n65564, n60507, n59153, n59095, 
        n60298, n67374, n59118, n68881, n69697, n69808, n69685, 
        n7_adj_5924, n68554, n68553, n68548;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5696));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n50289), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n27652), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i53364_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69092));
    defparam i53364_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4124[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .GND_net(GND_net), .state({state}), .bit_ctr({Open_0, Open_1, 
            Open_2, bit_ctr[1:0]}), .timer({timer}), .neopxl_color({neopxl_color}), 
            .n23(n23_adj_5922), .n43567(n43567), .n27950(n27950), .n29707(n29707), 
            .n111(n111), .VCC_net(VCC_net), .n30355(n30355), .n30354(n30354), 
            .n30353(n30353), .n30352(n30352), .n30351(n30351), .n30350(n30350), 
            .n30349(n30349), .n30348(n30348), .n30347(n30347), .n30342(n30342), 
            .n30251(n30251), .n5(n5_adj_5902), .NEOPXL_c(NEOPXL_c), .n25(n25_adj_5906), 
            .LED_c(LED_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_CARRY encoder0_position_30__I_0_add_1704_4 (.CI(n50289), .I0(n2532), 
            .I1(GND_net), .CO(n50290));
    SB_LUT4 i15726_3_lut (.I0(\data_in_frame[0] [7]), .I1(rx_data[7]), .I2(n7_adj_5921), 
            .I3(GND_net), .O(n29802));   // verilog/coms.v(130[12] 305[6])
    defparam i15726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n50288), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53085_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68813));
    defparam i53085_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(n36888), .I1(Ki[0]), .I2(GND_net), .I3(GND_net), 
            .O(n53));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53575_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69303));
    defparam i53575_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i835_3_lut (.I0(n1224_adj_5802), .I1(n1291), 
            .I2(n1257), .I3(GND_net), .O(n1323));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i835_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27728), 
            .D(n1219), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i53016_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68744));
    defparam i53016_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53012_1_lut (.I0(n43717), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68740));
    defparam i53012_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5890));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5888));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5889));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5886));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n3225), .I1(n27_adj_5890), .I2(n3292), .I3(n3237), 
            .O(n61528));
    defparam i1_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5887));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1980 (.I0(n3223), .I1(n19_adj_5888), .I2(n3290), 
            .I3(n3237), .O(n61524));
    defparam i1_4_lut_adj_1980.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1981 (.I0(n3227), .I1(n13_adj_5886), .I2(n3294), 
            .I3(n3237), .O(n61526));
    defparam i1_4_lut_adj_1981.LUT_INIT = 16'heefc;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n65588), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5854));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i50241_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n65578));
    defparam i50241_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_4_lut_adj_1982 (.I0(n3221), .I1(n23_adj_5889), .I2(n3288), 
            .I3(n3237), .O(n61530));
    defparam i1_4_lut_adj_1982.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1983 (.I0(n65578), .I1(n5_adj_5854), .I2(n65579), 
            .I3(n3237), .O(n53678));
    defparam i1_4_lut_adj_1983.LUT_INIT = 16'h88c0;
    SB_LUT4 i1_4_lut_adj_1984 (.I0(n61526), .I1(n61524), .I2(n15_adj_5887), 
            .I3(n61528), .O(n61538));
    defparam i1_4_lut_adj_1984.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5891));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1985 (.I0(n31_adj_5891), .I1(n61538), .I2(n53678), 
            .I3(n61530), .O(n61542));
    defparam i1_4_lut_adj_1985.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1986 (.I0(n3219), .I1(n61542), .I2(n3286), .I3(n3237), 
            .O(n61544));
    defparam i1_4_lut_adj_1986.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1987 (.I0(n3218), .I1(n61544), .I2(n3285), .I3(n3237), 
            .O(n61546));
    defparam i1_4_lut_adj_1987.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1988 (.I0(n3217), .I1(n61546), .I2(n3284), .I3(n3237), 
            .O(n61548));
    defparam i1_4_lut_adj_1988.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1989 (.I0(n3216), .I1(n61548), .I2(n3283), .I3(n3237), 
            .O(n61550));
    defparam i1_4_lut_adj_1989.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1990 (.I0(n3215), .I1(n61550), .I2(n3282), .I3(n3237), 
            .O(n61552));
    defparam i1_4_lut_adj_1990.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1991 (.I0(n3214), .I1(n61552), .I2(n3281), .I3(n3237), 
            .O(n61554));
    defparam i1_4_lut_adj_1991.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1992 (.I0(n3213), .I1(n61554), .I2(n3280), .I3(n3237), 
            .O(n61556));
    defparam i1_4_lut_adj_1992.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1993 (.I0(n3212), .I1(n61556), .I2(n3279), .I3(n3237), 
            .O(n61558));
    defparam i1_4_lut_adj_1993.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1994 (.I0(n3211), .I1(n61558), .I2(n3278), .I3(n3237), 
            .O(n61560));
    defparam i1_4_lut_adj_1994.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1995 (.I0(n3210), .I1(n61560), .I2(n3277), .I3(n3237), 
            .O(n61562));
    defparam i1_4_lut_adj_1995.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1996 (.I0(n3209), .I1(n61562), .I2(n3276), .I3(n3237), 
            .O(n61564));
    defparam i1_4_lut_adj_1996.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1997 (.I0(n3208), .I1(n61564), .I2(n3275), .I3(n3237), 
            .O(n61566));
    defparam i1_4_lut_adj_1997.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1998 (.I0(n3207), .I1(n61566), .I2(n3274), .I3(n3237), 
            .O(n61568));
    defparam i1_4_lut_adj_1998.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53015_4_lut (.I0(n61), .I1(n62647), .I2(n59), .I3(n61568), 
            .O(n43717));
    defparam i53015_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42499_3_lut (.I0(encoder0_position[27]), .I1(n58175), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut (.I0(dti_counter[0]), .I1(n14_adj_5904), .I2(n10_adj_5905), 
            .I3(dti_counter[3]), .O(n22917));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29610_4_lut (.I0(n520), .I1(n931), .I2(n932), .I3(n933), 
            .O(n43585));
    defparam i29610_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27728), 
            .D(n1218), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27728), 
            .D(n1217), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27728), 
            .D(n1216), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27728), 
            .D(n1215), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27728), 
            .D(n1214), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27728), 
            .D(n1213), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27728), 
            .D(n1212), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27728), 
            .D(n1211), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27728), 
            .D(n1210), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27728), 
            .D(n1209), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27728), 
            .D(n1208), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53558_2_lut (.I0(n22917), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i53558_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1999 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n61696));
    defparam i1_2_lut_adj_1999.LUT_INIT = 16'h8888;
    SB_LUT4 n11579_bdd_4_lut (.I0(n11579), .I1(current[15]), .I2(duty[22]), 
            .I3(n11577), .O(n69775));
    defparam n11579_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69775_bdd_4_lut (.I0(n69775), .I1(duty[19]), .I2(n4909), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[19]));
    defparam n69775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_4310_i10_3_lut (.I0(encoder0_position[9]), .I1(n23_adj_5708), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11579_bdd_4_lut_53989 (.I0(n11579), .I1(current[15]), .I2(duty[21]), 
            .I3(n11577), .O(n69769));
    defparam n11579_bdd_4_lut_53989.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69769_bdd_4_lut (.I0(n69769), .I1(duty[18]), .I2(n4910), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[18]));
    defparam n69769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i14_3_lut (.I0(encoder0_position[13]), .I1(n19_adj_5712), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11579_bdd_4_lut_53984 (.I0(n11579), .I1(current[15]), .I2(duty[20]), 
            .I3(n11577), .O(n69763));
    defparam n11579_bdd_4_lut_53984.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69763_bdd_4_lut (.I0(n69763), .I1(duty[17]), .I2(n4911), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[17]));
    defparam n69763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53979 (.I0(n11579), .I1(current[15]), .I2(duty[19]), 
            .I3(n11577), .O(n69757));
    defparam n11579_bdd_4_lut_53979.LUT_INIT = 16'he4aa;
    SB_LUT4 n69757_bdd_4_lut (.I0(n69757), .I1(duty[16]), .I2(n4912), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[16]));
    defparam n69757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i1_3_lut (.I0(encoder0_position[0]), .I1(n32), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2000 (.I0(n3228), .I1(n3216), .I2(n3224), .I3(n3227), 
            .O(n62068));
    defparam i1_4_lut_adj_2000.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2001 (.I0(n3217), .I1(n3222), .I2(n3226), .I3(n3218), 
            .O(n62070));
    defparam i1_4_lut_adj_2001.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2002 (.I0(n3221), .I1(n3225), .I2(GND_net), .I3(GND_net), 
            .O(n62060));
    defparam i1_2_lut_adj_2002.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut (.I0(n62068), .I1(n3223), .I2(n3220), .I3(GND_net), 
            .O(n62072));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2003 (.I0(n62060), .I1(n3215), .I2(n62070), .I3(n3219), 
            .O(n62076));
    defparam i1_4_lut_adj_2003.LUT_INIT = 16'hfffe;
    SB_LUT4 i29712_4_lut (.I0(n957), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n43687));
    defparam i29712_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2004 (.I0(n3213), .I1(n3214), .I2(n62076), .I3(n62072), 
            .O(n62082));
    defparam i1_4_lut_adj_2004.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2005 (.I0(n3229), .I1(n62082), .I2(n43687), .I3(n3230), 
            .O(n62084));
    defparam i1_4_lut_adj_2005.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2006 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n62084), 
            .O(n62090));
    defparam i1_4_lut_adj_2006.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2007 (.I0(n927), .I1(n61696), .I2(n928), .I3(n43585), 
            .O(n960));
    defparam i1_4_lut_adj_2007.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_2008 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n62090), 
            .O(n62096));
    defparam i1_4_lut_adj_2008.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53047_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n62096), 
            .O(n3237));
    defparam i53047_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29614_3_lut (.I0(n521), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n43589));
    defparam i29614_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i42494_3_lut (.I0(n3), .I1(n7451), .I2(n58170), .I3(GND_net), 
            .O(n58171));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i2_3_lut (.I0(encoder0_position[1]), .I1(n31), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2009 (.I0(n3121), .I1(n3128), .I2(n3127), .I3(n3126), 
            .O(n61454));
    defparam i1_4_lut_adj_2009.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2010 (.I0(n3124), .I1(n3123), .I2(n3125), .I3(n3122), 
            .O(n61452));
    defparam i1_4_lut_adj_2010.LUT_INIT = 16'hfffe;
    SB_LUT4 i29567_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n43541));
    defparam i29567_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2011 (.I0(n3119), .I1(n61452), .I2(n61454), .I3(n3120), 
            .O(n61460));
    defparam i1_4_lut_adj_2011.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2012 (.I0(n3129), .I1(n43541), .I2(n3130), .I3(n3131), 
            .O(n59118));
    defparam i1_4_lut_adj_2012.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2013 (.I0(n59118), .I1(n3117), .I2(n3118), .I3(n61460), 
            .O(n61466));
    defparam i1_4_lut_adj_2013.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2014 (.I0(n3114), .I1(n3115), .I2(n3116), .I3(n61466), 
            .O(n61472));
    defparam i1_4_lut_adj_2014.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2015 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n61472), 
            .O(n61478));
    defparam i1_4_lut_adj_2015.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2016 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n61478), 
            .O(n61484));
    defparam i1_4_lut_adj_2016.LUT_INIT = 16'hfffe;
    SB_LUT4 i53118_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n61484), 
            .O(n3138));
    defparam i53118_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2017 (.I0(n1029), .I1(n43589), .I2(n1030), .I3(n1031), 
            .O(n59018));
    defparam i1_4_lut_adj_2017.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42495_3_lut (.I0(encoder0_position[29]), .I1(n58171), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i3_3_lut (.I0(encoder0_position[2]), .I1(n30), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53653_4_lut (.I0(n1026), .I1(n59018), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i53653_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53081_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68809));
    defparam i53081_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2018 (.I0(n3021), .I1(n3022), .I2(n3025), .I3(n3023), 
            .O(n61954));
    defparam i1_4_lut_adj_2018.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2019 (.I0(n3028), .I1(n3017), .I2(n3024), .I3(n3020), 
            .O(n61956));
    defparam i1_4_lut_adj_2019.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2020 (.I0(n3026), .I1(n3019), .I2(n3018), .I3(n3027), 
            .O(n61958));
    defparam i1_4_lut_adj_2020.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2021 (.I0(n3016), .I1(n61958), .I2(n61956), .I3(n61954), 
            .O(n61964));
    defparam i1_4_lut_adj_2021.LUT_INIT = 16'hfffe;
    SB_LUT4 i29563_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n43537));
    defparam i29563_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_2022 (.I0(n3014), .I1(n3015), .I2(n61964), .I3(GND_net), 
            .O(n61968));
    defparam i1_3_lut_adj_2022.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2023 (.I0(n3029), .I1(n43537), .I2(n3030), .I3(n3031), 
            .O(n59153));
    defparam i1_4_lut_adj_2023.LUT_INIT = 16'ha080;
    SB_LUT4 n11579_bdd_4_lut_53974 (.I0(n11579), .I1(current[15]), .I2(duty[18]), 
            .I3(n11577), .O(n69751));
    defparam n11579_bdd_4_lut_53974.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_2024 (.I0(n3012), .I1(n3013), .I2(n59153), .I3(n61968), 
            .O(n61974));
    defparam i1_4_lut_adj_2024.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2025 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n61974), 
            .O(n61980));
    defparam i1_4_lut_adj_2025.LUT_INIT = 16'hfffe;
    SB_LUT4 i53084_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n61980), 
            .O(n3039));
    defparam i53084_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29688_4_lut (.I0(n522), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n43663));
    defparam i29688_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2026 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n61688));
    defparam i1_3_lut_adj_2026.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1919_3_lut (.I0(n2820_adj_5823), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225_adj_5803));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2027 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n61700));
    defparam i1_2_lut_adj_2027.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i836_3_lut (.I0(n1225_adj_5803), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i4_3_lut (.I0(encoder0_position[3]), .I1(n29), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53153_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68881));
    defparam i53153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_2028 (.I0(n2925), .I1(n2924), .I2(n2927), .I3(GND_net), 
            .O(n61644));
    defparam i1_3_lut_adj_2028.LUT_INIT = 16'hfefe;
    SB_LUT4 i53572_4_lut (.I0(n61700), .I1(n1125), .I2(n61688), .I3(n43663), 
            .O(n1158));
    defparam i53572_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i29694_4_lut (.I0(n954), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n43669));
    defparam i29694_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2029 (.I0(n2921), .I1(n61644), .I2(n2923), .I3(n2928), 
            .O(n61648));
    defparam i1_4_lut_adj_2029.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2030 (.I0(n2926), .I1(n2922), .I2(GND_net), .I3(GND_net), 
            .O(n61896));
    defparam i1_2_lut_adj_2030.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2031 (.I0(n2929), .I1(n61648), .I2(n43669), .I3(n2930), 
            .O(n61650));
    defparam i1_4_lut_adj_2031.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2032 (.I0(n2918), .I1(n2920), .I2(n2919), .I3(n61896), 
            .O(n61652));
    defparam i1_4_lut_adj_2032.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2033 (.I0(n2916), .I1(n2917), .I2(n61652), .I3(n61650), 
            .O(n61658));
    defparam i1_4_lut_adj_2033.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2034 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n61658), 
            .O(n61664));
    defparam i1_4_lut_adj_2034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2035 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n61664), 
            .O(n61670));
    defparam i1_4_lut_adj_2035.LUT_INIT = 16'hfffe;
    SB_LUT4 i53156_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n61670), 
            .O(n2940));
    defparam i53156_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1840_3_lut (.I0(n2709), .I1(n2776), 
            .I2(n2742), .I3(GND_net), .O(n2808));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_3 (.CI(n50288), .I0(n2533), 
            .I1(VCC_net), .CO(n50289));
    SB_LUT4 encoder0_position_30__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n50288));
    SB_LUT4 encoder0_position_30__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_24_lut (.I0(n69006), .I1(n2412), 
            .I2(VCC_net), .I3(n50287), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n50286), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_23 (.CI(n50286), .I0(n2413), 
            .I1(VCC_net), .CO(n50287));
    SB_LUT4 encoder0_position_30__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n50285), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_22 (.CI(n50285), .I0(n2414), 
            .I1(VCC_net), .CO(n50286));
    SB_LUT4 encoder0_position_30__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n50284), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820_adj_5823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_21 (.CI(n50284), .I0(n2415), 
            .I1(VCC_net), .CO(n50285));
    SB_LUT4 encoder0_position_30__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n50283), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i5_3_lut (.I0(encoder0_position[4]), .I1(n28), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1637_20 (.CI(n50283), .I0(n2416), 
            .I1(VCC_net), .CO(n50284));
    SB_LUT4 encoder0_position_30__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n50282), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53187_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68915));
    defparam i53187_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_19 (.CI(n50282), .I0(n2417), 
            .I1(VCC_net), .CO(n50283));
    SB_LUT4 n69751_bdd_4_lut (.I0(n69751), .I1(duty[15]), .I2(n4913), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[15]));
    defparam n69751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_2036 (.I0(n2827), .I1(n2819), .I2(n2826), .I3(n2820_adj_5823), 
            .O(n61914));
    defparam i1_4_lut_adj_2036.LUT_INIT = 16'hfffe;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n50281), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2037 (.I0(n2828), .I1(n2818), .I2(n2825), .I3(n2823), 
            .O(n61916));
    defparam i1_4_lut_adj_2037.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2038 (.I0(n61914), .I1(n2822), .I2(n2821), .I3(GND_net), 
            .O(n61918));
    defparam i1_3_lut_adj_2038.LUT_INIT = 16'hfefe;
    SB_LUT4 i29696_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n43671));
    defparam i29696_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2039 (.I0(n2816), .I1(n2817), .I2(n61918), .I3(n61916), 
            .O(n61924));
    defparam i1_4_lut_adj_2039.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2040 (.I0(n2829), .I1(n61924), .I2(n43671), .I3(n2830), 
            .O(n61926));
    defparam i1_4_lut_adj_2040.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2041 (.I0(n2814), .I1(n2812), .I2(n2815), .I3(n2824), 
            .O(n59279));
    defparam i1_4_lut_adj_2041.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2042 (.I0(n59279), .I1(n2811), .I2(n2813), .I3(n61926), 
            .O(n61932));
    defparam i1_4_lut_adj_2042.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1637_18 (.CI(n50281), .I0(n2418), 
            .I1(VCC_net), .CO(n50282));
    SB_LUT4 i53190_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n61932), 
            .O(n2841));
    defparam i53190_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53969 (.I0(n11579), .I1(current[15]), .I2(duty[17]), 
            .I3(n11577), .O(n69745));
    defparam n11579_bdd_4_lut_53969.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n50280), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_17 (.CI(n50280), .I0(n2419), 
            .I1(VCC_net), .CO(n50281));
    SB_LUT4 encoder0_position_30__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n50279), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_16 (.CI(n50279), .I0(n2420), 
            .I1(VCC_net), .CO(n50280));
    SB_LUT4 encoder0_position_30__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n50278), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_15 (.CI(n50278), .I0(n2421), 
            .I1(VCC_net), .CO(n50279));
    SB_LUT4 encoder0_position_30__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n50277), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_14 (.CI(n50277), .I0(n2422), 
            .I1(VCC_net), .CO(n50278));
    SB_LUT4 encoder0_position_30__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n50276), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut (.I0(hall1), .I1(hall2), .I2(n20965), .I3(GND_net), 
            .O(n4_adj_5913));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 encoder0_position_30__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1034_15_lut (.I0(n69333), .I1(n1521), 
            .I2(VCC_net), .I3(n49999), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n49998), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_13 (.CI(n50276), .I0(n2423), 
            .I1(VCC_net), .CO(n50277));
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_30__I_0_add_1034_14 (.CI(n49998), .I0(n1522), 
            .I1(VCC_net), .CO(n49999));
    SB_LUT4 encoder0_position_30__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n50275), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n49997), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_13 (.CI(n49997), .I0(n1523), 
            .I1(VCC_net), .CO(n49998));
    SB_LUT4 encoder0_position_30__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n49996), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_12 (.CI(n50275), .I0(n2424), 
            .I1(VCC_net), .CO(n50276));
    SB_CARRY encoder0_position_30__I_0_add_1034_12 (.CI(n49996), .I0(n1524), 
            .I1(VCC_net), .CO(n49997));
    SB_LUT4 encoder0_position_30__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n50274), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4310_i6_3_lut (.I0(encoder0_position[5]), .I1(n27), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_11 (.CI(n50274), .I0(n2425), 
            .I1(VCC_net), .CO(n50275));
    SB_LUT4 encoder0_position_30__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n49995), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n50273), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i53220_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68948));
    defparam i53220_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_10 (.CI(n50273), .I0(n2426), 
            .I1(VCC_net), .CO(n50274));
    SB_LUT4 i29646_3_lut (.I0(n952), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n43621));
    defparam i29646_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n50272), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n69745_bdd_4_lut (.I0(n69745), .I1(duty[14]), .I2(n4914), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[14]));
    defparam n69745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_2043 (.I0(n2724), .I1(n2728), .I2(n2725), .I3(GND_net), 
            .O(n61424));
    defparam i1_3_lut_adj_2043.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2044 (.I0(n2720), .I1(n61424), .I2(n2726), .I3(n2722), 
            .O(n61428));
    defparam i1_4_lut_adj_2044.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2045 (.I0(n2729), .I1(n43621), .I2(n2730), .I3(n2731), 
            .O(n59095));
    defparam i1_4_lut_adj_2045.LUT_INIT = 16'ha080;
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 i1_4_lut_adj_2046 (.I0(n2717), .I1(n2718), .I2(n59095), .I3(n61428), 
            .O(n61434));
    defparam i1_4_lut_adj_2046.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2047 (.I0(n2719), .I1(n2721), .I2(n2723), .I3(n2727), 
            .O(n61602));
    defparam i1_4_lut_adj_2047.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2048 (.I0(n2713), .I1(n2715), .I2(n2716), .I3(n61434), 
            .O(n61440));
    defparam i1_4_lut_adj_2048.LUT_INIT = 16'hfffe;
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_1034_11 (.CI(n49995), .I0(n1525), 
            .I1(VCC_net), .CO(n49996));
    SB_LUT4 i1_4_lut_adj_2049 (.I0(n2710), .I1(n2712), .I2(n2714), .I3(n61602), 
            .O(n61608));
    defparam i1_4_lut_adj_2049.LUT_INIT = 16'hfffe;
    SB_LUT4 i53223_4_lut (.I0(n2711), .I1(n61608), .I2(n61440), .I3(n2709), 
            .O(n2742));
    defparam i53223_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n49994), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53964 (.I0(n11579), .I1(current[15]), .I2(duty[16]), 
            .I3(n11577), .O(n69739));
    defparam n11579_bdd_4_lut_53964.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_9 (.CI(n50272), .I0(n2427), 
            .I1(VCC_net), .CO(n50273));
    SB_CARRY encoder0_position_30__I_0_add_1034_10 (.CI(n49994), .I0(n1526), 
            .I1(VCC_net), .CO(n49995));
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n50271), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n49993), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1034_9 (.CI(n49993), .I0(n1527), 
            .I1(VCC_net), .CO(n49994));
    SB_CARRY encoder0_position_30__I_0_add_1637_8 (.CI(n50271), .I0(n2428), 
            .I1(VCC_net), .CO(n50272));
    SB_LUT4 encoder0_position_30__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69739_bdd_4_lut (.I0(n69739), .I1(duty[13]), .I2(n4915), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[13]));
    defparam n69739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n49992), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n50270), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_8 (.CI(n49992), .I0(n1528), 
            .I1(VCC_net), .CO(n49993));
    SB_LUT4 encoder0_position_30__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n49991), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_7 (.CI(n49991), .I0(n1529), 
            .I1(GND_net), .CO(n49992));
    SB_LUT4 encoder0_position_30__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28329_3_lut (.I0(current[11]), .I1(data_adj_5985[11]), .I2(n27736), 
            .I3(GND_net), .O(n30417));
    defparam i28329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16342_3_lut (.I0(current[10]), .I1(data_adj_5985[10]), .I2(n27736), 
            .I3(GND_net), .O(n30418));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16343_3_lut (.I0(current[9]), .I1(data_adj_5985[9]), .I2(n27736), 
            .I3(GND_net), .O(n30419));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16344_3_lut (.I0(current[8]), .I1(data_adj_5985[8]), .I2(n27736), 
            .I3(GND_net), .O(n30420));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16345_3_lut (.I0(current[7]), .I1(data_adj_5985[7]), .I2(n27736), 
            .I3(GND_net), .O(n30421));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16346_3_lut (.I0(current[6]), .I1(data_adj_5985[6]), .I2(n27736), 
            .I3(GND_net), .O(n30422));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16347_3_lut (.I0(current[5]), .I1(data_adj_5985[5]), .I2(n27736), 
            .I3(GND_net), .O(n30423));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i7_3_lut (.I0(encoder0_position[6]), .I1(n26_adj_5705), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53335_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69063));
    defparam i53335_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_2050 (.I0(n2627), .I1(n2623), .I2(GND_net), .I3(GND_net), 
            .O(n62040));
    defparam i1_2_lut_adj_2050.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2051 (.I0(n2621), .I1(n2618), .I2(n2624), .I3(n2620), 
            .O(n60332));
    defparam i1_4_lut_adj_2051.LUT_INIT = 16'hfffe;
    SB_LUT4 i29644_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n43619));
    defparam i29644_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16348_3_lut (.I0(current[4]), .I1(data_adj_5985[4]), .I2(n27736), 
            .I3(GND_net), .O(n30424));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16349_3_lut (.I0(current[3]), .I1(data_adj_5985[3]), .I2(n27736), 
            .I3(GND_net), .O(n30425));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16350_3_lut (.I0(current[2]), .I1(data_adj_5985[2]), .I2(n27736), 
            .I3(GND_net), .O(n30426));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16351_3_lut (.I0(current[1]), .I1(data_adj_5985[1]), .I2(n27736), 
            .I3(GND_net), .O(n30427));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2052 (.I0(n2617), .I1(n2619), .I2(n62040), .I3(n2625), 
            .O(n62046));
    defparam i1_4_lut_adj_2052.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2053 (.I0(n2629), .I1(n43619), .I2(n2630), .I3(n2631), 
            .O(n59130));
    defparam i1_4_lut_adj_2053.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2054 (.I0(n60332), .I1(n2628), .I2(n2626), .I3(n2622), 
            .O(n61880));
    defparam i1_4_lut_adj_2054.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1637_7 (.CI(n50270), .I0(n2429), 
            .I1(GND_net), .CO(n50271));
    SB_LUT4 i1_4_lut_adj_2055 (.I0(n2616), .I1(n2615), .I2(n59130), .I3(n62046), 
            .O(n60331));
    defparam i1_4_lut_adj_2055.LUT_INIT = 16'hfffe;
    SB_LUT4 i16356_3_lut (.I0(baudrate[31]), .I1(data_adj_5978[7]), .I2(n28027), 
            .I3(GND_net), .O(n30432));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2056 (.I0(n2613), .I1(n2614), .I2(n60331), .I3(n61880), 
            .O(n61886));
    defparam i1_4_lut_adj_2056.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n50269), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n49990), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16357_3_lut (.I0(baudrate[30]), .I1(data_adj_5978[6]), .I2(n28027), 
            .I3(GND_net), .O(n30433));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16357_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1637_6 (.CI(n50269), .I0(n2430), 
            .I1(GND_net), .CO(n50270));
    SB_CARRY encoder0_position_30__I_0_add_1034_6 (.CI(n49990), .I0(n1530), 
            .I1(GND_net), .CO(n49991));
    SB_LUT4 encoder0_position_30__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n50268), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_5 (.CI(n50268), .I0(n2431), 
            .I1(VCC_net), .CO(n50269));
    SB_LUT4 encoder0_position_30__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n49989), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16358_3_lut (.I0(baudrate[29]), .I1(data_adj_5978[5]), .I2(n28027), 
            .I3(GND_net), .O(n30434));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16359_3_lut (.I0(baudrate[28]), .I1(data_adj_5978[4]), .I2(n28027), 
            .I3(GND_net), .O(n30435));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53338_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n61886), 
            .O(n2643));
    defparam i53338_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16360_3_lut (.I0(baudrate[27]), .I1(data_adj_5978[3]), .I2(n28027), 
            .I3(GND_net), .O(n30436));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16361_3_lut (.I0(baudrate[26]), .I1(data_adj_5978[2]), .I2(n28027), 
            .I3(GND_net), .O(n30437));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16362_3_lut (.I0(baudrate[25]), .I1(data_adj_5978[1]), .I2(n28027), 
            .I3(GND_net), .O(n30438));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16362_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1034_5 (.CI(n49989), .I0(n1531), 
            .I1(VCC_net), .CO(n49990));
    SB_LUT4 encoder0_position_30__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n50267), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_4 (.CI(n50267), .I0(n2432), 
            .I1(GND_net), .CO(n50268));
    SB_LUT4 encoder0_position_30__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n50266), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n49988), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_3 (.CI(n50266), .I0(n2433), 
            .I1(VCC_net), .CO(n50267));
    SB_LUT4 encoder0_position_30__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_4 (.CI(n49988), .I0(n1532), 
            .I1(GND_net), .CO(n49989));
    SB_CARRY encoder0_position_30__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n50266));
    SB_LUT4 encoder0_position_30__I_0_add_1570_23_lut (.I0(n68974), .I1(n2313), 
            .I2(VCC_net), .I3(n50265), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n50264), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_22 (.CI(n50264), .I0(n2314), 
            .I1(VCC_net), .CO(n50265));
    SB_LUT4 encoder0_position_30__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n50263), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_21 (.CI(n50263), .I0(n2315), 
            .I1(VCC_net), .CO(n50264));
    SB_LUT4 encoder0_position_30__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16364_3_lut (.I0(baudrate[24]), .I1(data_adj_5978[0]), .I2(n28027), 
            .I3(GND_net), .O(n30440));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n50262), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_20 (.CI(n50262), .I0(n2316), 
            .I1(VCC_net), .CO(n50263));
    SB_LUT4 encoder0_position_30__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n49987), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15688_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n7_adj_5921), 
            .I3(GND_net), .O(n29764));   // verilog/coms.v(130[12] 305[6])
    defparam i15688_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53959 (.I0(n11579), .I1(current[15]), .I2(duty[15]), 
            .I3(n11577), .O(n69733));
    defparam n11579_bdd_4_lut_53959.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n50261), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_19 (.CI(n50261), .I0(n2317), 
            .I1(VCC_net), .CO(n50262));
    SB_LUT4 encoder0_position_30__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n50260), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5695));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_18 (.CI(n50260), .I0(n2318), 
            .I1(VCC_net), .CO(n50261));
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5694));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5693));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5692));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5691));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1034_3 (.CI(n49987), .I0(n1533), 
            .I1(VCC_net), .CO(n49988));
    SB_LUT4 encoder0_position_30__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n50259), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_17 (.CI(n50259), .I0(n2319), 
            .I1(VCC_net), .CO(n50260));
    SB_LUT4 i15663_3_lut (.I0(\data_in_frame[0] [2]), .I1(rx_data[2]), .I2(n7_adj_5921), 
            .I3(GND_net), .O(n29739));   // verilog/coms.v(130[12] 305[6])
    defparam i15663_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n49987));
    SB_LUT4 encoder0_position_30__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n50258), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_16 (.CI(n50258), .I0(n2320), 
            .I1(VCC_net), .CO(n50259));
    SB_LUT4 encoder0_position_30__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n50257), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5690));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_15 (.CI(n50257), .I0(n2321), 
            .I1(VCC_net), .CO(n50258));
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5689));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5688));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n50256), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_14 (.CI(n50256), .I0(n2322), 
            .I1(VCC_net), .CO(n50257));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69733_bdd_4_lut (.I0(n69733), .I1(duty[12]), .I2(n4916), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[12]));
    defparam n69733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53954 (.I0(n11579), .I1(current[11]), .I2(duty[14]), 
            .I3(n11577), .O(n69727));
    defparam n11579_bdd_4_lut_53954.LUT_INIT = 16'he4aa;
    SB_LUT4 i53306_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69034));
    defparam i53306_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2057 (.I0(n2525), .I1(n2526), .I2(n2524), .I3(n2523), 
            .O(n61496));
    defparam i1_4_lut_adj_2057.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2058 (.I0(n2522), .I1(n2528), .I2(n2527), .I3(GND_net), 
            .O(n61498));
    defparam i1_3_lut_adj_2058.LUT_INIT = 16'hfefe;
    SB_LUT4 i29702_4_lut (.I0(n950), .I1(n2531), .I2(n2532), .I3(n2533), 
            .O(n43677));
    defparam i29702_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2059 (.I0(n2520), .I1(n2521), .I2(n61498), .I3(n61496), 
            .O(n61504));
    defparam i1_4_lut_adj_2059.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2060 (.I0(n2529), .I1(n61504), .I2(n43677), .I3(n2530), 
            .O(n61506));
    defparam i1_4_lut_adj_2060.LUT_INIT = 16'heccc;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15824_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n61106), 
            .I3(n27_adj_5825), .O(n29900));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15824_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n69727_bdd_4_lut (.I0(n69727), .I1(duty[11]), .I2(n4917), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[11]));
    defparam n69727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n50255), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2061 (.I0(n2517), .I1(n2518), .I2(n61506), .I3(n2519), 
            .O(n61512));
    defparam i1_4_lut_adj_2061.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1570_13 (.CI(n50255), .I0(n2323), 
            .I1(VCC_net), .CO(n50256));
    SB_LUT4 i1_4_lut_adj_2062 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n61512), 
            .O(n61518));
    defparam i1_4_lut_adj_2062.LUT_INIT = 16'hfffe;
    SB_LUT4 i53309_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n61518), 
            .O(n2544));
    defparam i53309_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i53278_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69006));
    defparam i53278_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53246_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68974));
    defparam i53246_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16397_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .I2(control_update), .I3(GND_net), .O(n30473));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53432_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69160));
    defparam i53432_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16398_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I2(control_update), .I3(GND_net), .O(n30474));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16399_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .I2(control_update), .I3(GND_net), .O(n30475));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53407_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69135));
    defparam i53407_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53360_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69088));
    defparam i53360_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53456_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69184));
    defparam i53456_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16400_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I2(control_update), .I3(GND_net), .O(n30476));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53478_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69206));
    defparam i53478_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22787_3_lut (.I0(n212), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(n36823));
    defparam i22787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22788_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n36823), 
            .I2(control_update), .I3(GND_net), .O(n30477));   // verilog/motorControl.v(20[7:21])
    defparam i22788_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n50254), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22817_3_lut (.I0(n213), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(n36852));
    defparam i22817_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1570_12 (.CI(n50254), .I0(n2324), 
            .I1(VCC_net), .CO(n50255));
    SB_LUT4 i53497_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69225));
    defparam i53497_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22818_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n36852), 
            .I2(control_update), .I3(GND_net), .O(n30478));   // verilog/motorControl.v(20[7:21])
    defparam i22818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11579_bdd_4_lut_53949 (.I0(n11579), .I1(current[10]), .I2(duty[13]), 
            .I3(n11577), .O(n69721));
    defparam n11579_bdd_4_lut_53949.LUT_INIT = 16'he4aa;
    SB_LUT4 i22854_3_lut (.I0(n214), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(n36888));
    defparam i22854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53605_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69333));
    defparam i53605_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n50253), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n69721_bdd_4_lut (.I0(n69721), .I1(duty[10]), .I2(n4918), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[10]));
    defparam n69721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_1570_11 (.CI(n50253), .I0(n2325), 
            .I1(VCC_net), .CO(n50254));
    SB_LUT4 encoder0_position_30__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n50252), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53622_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69350));
    defparam i53622_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_10 (.CI(n50252), .I0(n2326), 
            .I1(VCC_net), .CO(n50253));
    SB_LUT4 i22855_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n36888), 
            .I2(control_update), .I3(GND_net), .O(n30479));   // verilog/motorControl.v(20[7:21])
    defparam i22855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n50251), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53637_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69365));
    defparam i53637_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_9 (.CI(n50251), .I0(n2327), 
            .I1(VCC_net), .CO(n50252));
    SB_LUT4 i53569_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69297));
    defparam i53569_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[22] [7]), .I1(n8_adj_5801), .I2(n43396), 
            .I3(n57336), .O(n56398));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i53650_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69378));
    defparam i53650_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16404_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(control_update), .I3(GND_net), .O(n30480));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16405_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(control_update), .I3(GND_net), .O(n30481));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16406_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(control_update), .I3(GND_net), .O(n30482));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n50250), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_8 (.CI(n50250), .I0(n2328), 
            .I1(VCC_net), .CO(n50251));
    SB_LUT4 i16407_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(control_update), .I3(GND_net), .O(n30483));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22497_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(control_update), .I3(GND_net), .O(n30484));   // verilog/motorControl.v(20[7:21])
    defparam i22497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16409_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(control_update), .I3(GND_net), .O(n30485));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16410_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(control_update), .I3(GND_net), .O(n30486));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n50249), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_7 (.CI(n50249), .I0(n2329), 
            .I1(GND_net), .CO(n50250));
    SB_LUT4 encoder0_position_30__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n50248), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11579_bdd_4_lut_53944 (.I0(n11579), .I1(current[9]), .I2(duty[12]), 
            .I3(n11577), .O(n69715));
    defparam n11579_bdd_4_lut_53944.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1570_6 (.CI(n50248), .I0(n2330), 
            .I1(GND_net), .CO(n50249));
    SB_LUT4 i16411_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(control_update), .I3(GND_net), .O(n30487));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16412_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(control_update), .I3(GND_net), .O(n30488));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n50247), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_5 (.CI(n50247), .I0(n2331), 
            .I1(VCC_net), .CO(n50248));
    SB_LUT4 n69715_bdd_4_lut (.I0(n69715), .I1(duty[9]), .I2(n4919), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n69715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i42496_3_lut (.I0(n4_adj_5730), .I1(n7452), .I2(n58170), .I3(GND_net), 
            .O(n58173));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16413_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(control_update), .I3(GND_net), .O(n30489));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16415_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(control_update), .I3(GND_net), .O(n30491));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16417_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(control_update), .I3(GND_net), .O(n30493));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16418_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(control_update), .I3(GND_net), .O(n30494));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16419_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(control_update), .I3(GND_net), .O(n30495));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n50246), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16420_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(control_update), .I3(GND_net), .O(n30496));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16421_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(control_update), .I3(GND_net), .O(n30497));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut (.I0(hall2), .I1(commutation_state_7__N_27[2]), .I2(GND_net), 
            .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i16430_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n57425), .I3(GND_net), .O(n30506));   // verilog/coms.v(130[12] 305[6])
    defparam i16430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2063 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_2063.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2820), .O(n25_adj_5898));   // verilog/TinyFPGA_B.v(376[7:11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 i16436_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n57425), .I3(GND_net), .O(n30512));   // verilog/coms.v(130[12] 305[6])
    defparam i16436_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1438_3_lut (.I0(n2115), .I1(n2182), 
            .I2(n2148), .I3(GND_net), .O(n2214));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14826_2_lut (.I0(n27676), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14826_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52880_4_lut (.I0(commutation_state[1]), .I1(n22917), .I2(dti), 
            .I3(commutation_state[2]), .O(n27676));
    defparam i52880_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i16443_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n20965), .I3(n4_adj_5913), .O(n30519));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i16443_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i29616_3_lut (.I0(n523), .I1(n1232_adj_5810), .I2(n1233_adj_5811), 
            .I3(GND_net), .O(n43591));
    defparam i29616_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_30__I_0_add_1570_4 (.CI(n50246), .I0(n2332), 
            .I1(GND_net), .CO(n50247));
    SB_LUT4 i15401_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n57425), .I3(GND_net), .O(n29477));   // verilog/coms.v(130[12] 305[6])
    defparam i15401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n50245), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_3 (.CI(n50245), .I0(n2333), 
            .I1(VCC_net), .CO(n50246));
    SB_LUT4 encoder0_position_30__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n49521), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n50245));
    SB_LUT4 i15836_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n61058), 
            .I3(n27_adj_5825), .O(n29912));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15836_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1503_22_lut (.I0(n69160), .I1(n2214), 
            .I2(VCC_net), .I3(n50244), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n50243), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16447_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[0]), 
            .I2(n10_adj_5892), .I3(n25600), .O(n30523));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16447_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_1503_21 (.CI(n50243), .I0(n2215), 
            .I1(VCC_net), .CO(n50244));
    SB_LUT4 encoder0_position_30__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n50242), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_20 (.CI(n50242), .I0(n2216), 
            .I1(VCC_net), .CO(n50243));
    SB_LUT4 encoder0_position_30__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n50241), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_19 (.CI(n50241), .I0(n2217), 
            .I1(VCC_net), .CO(n50242));
    SB_LUT4 encoder0_position_30__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n50240), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_14_lut (.I0(n69350), .I1(n1422), 
            .I2(VCC_net), .I3(n49962), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n49961), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4310_i12_3_lut (.I0(encoder0_position[11]), .I1(n21_adj_5710), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_967_13 (.CI(n49961), .I0(n1423), 
            .I1(VCC_net), .CO(n49962));
    SB_LUT4 encoder0_position_30__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n49960), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_12 (.CI(n49960), .I0(n1424), 
            .I1(VCC_net), .CO(n49961));
    SB_CARRY encoder0_position_30__I_0_add_1503_18 (.CI(n50240), .I0(n2218), 
            .I1(VCC_net), .CO(n50241));
    SB_LUT4 encoder0_position_30__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n50239), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n49959), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_17 (.CI(n50239), .I0(n2219), 
            .I1(VCC_net), .CO(n50240));
    SB_CARRY encoder0_position_30__I_0_add_967_11 (.CI(n49959), .I0(n1425), 
            .I1(VCC_net), .CO(n49960));
    SB_LUT4 encoder0_position_30__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n49958), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n50238), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_16 (.CI(n50238), .I0(n2220), 
            .I1(VCC_net), .CO(n50239));
    SB_LUT4 i16453_3_lut (.I0(n58373), .I1(r_Bit_Index[0]), .I2(n27996), 
            .I3(GND_net), .O(n30529));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16453_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_30__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n50237), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_10 (.CI(n49958), .I0(n1426), 
            .I1(VCC_net), .CO(n49959));
    SB_LUT4 encoder0_position_30__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n49957), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4310_i13_3_lut (.I0(encoder0_position[12]), .I1(n20_adj_5711), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_967_9 (.CI(n49957), .I0(n1427), 
            .I1(VCC_net), .CO(n49958));
    SB_LUT4 encoder0_position_30__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1503_15 (.CI(n50237), .I0(n2221), 
            .I1(VCC_net), .CO(n50238));
    SB_LUT4 i16457_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n61138), 
            .I3(n27_adj_5825), .O(n30533));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16457_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15638_3_lut (.I0(\data_in_frame[22] [6]), .I1(rx_data[6]), 
            .I2(n43396), .I3(GND_net), .O(n29714));   // verilog/coms.v(130[12] 305[6])
    defparam i15638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16458_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n7_adj_5921), 
            .I3(GND_net), .O(n30534));   // verilog/coms.v(130[12] 305[6])
    defparam i16458_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15398_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n57425), .I3(GND_net), .O(n29474));   // verilog/coms.v(130[12] 305[6])
    defparam i15398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53939 (.I0(n11579), .I1(current[8]), .I2(duty[11]), 
            .I3(n11577), .O(n69709));
    defparam n11579_bdd_4_lut_53939.LUT_INIT = 16'he4aa;
    SB_LUT4 i16462_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[0]), .I2(n11_adj_5751), 
            .I3(state_7__N_4317), .O(n30538));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16462_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30_4_lut (.I0(state_7__N_3916[0]), .I1(n25471), .I2(state_adj_5979[1]), 
            .I3(n57392), .O(n12_adj_5919));   // verilog/eeprom.v(35[8] 81[4])
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12_adj_5919), .I1(n65782), .I2(state_adj_5979[0]), 
            .I3(state_adj_5979[2]), .O(n56570));   // verilog/eeprom.v(35[8] 81[4])
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n49956), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i584_2_lut (.I0(n1319), .I1(n42725), .I2(GND_net), .I3(GND_net), 
            .O(n2820));   // verilog/TinyFPGA_B.v(383[18] 385[12])
    defparam i584_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50238_4_lut (.I0(data_ready), .I1(n6617), .I2(n24_adj_5896), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n65737));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i50238_4_lut.LUT_INIT = 16'hdccc;
    SB_CARRY encoder0_position_30__I_0_add_967_8 (.CI(n49956), .I0(n1428), 
            .I1(VCC_net), .CO(n49957));
    SB_LUT4 i50870_2_lut (.I0(n24_adj_5896), .I1(n6617), .I2(GND_net), 
            .I3(GND_net), .O(n65740));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i50870_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n49955), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n50236), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49_4_lut (.I0(n65740), .I1(n65737), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5912), .O(n55644));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_CARRY encoder0_position_30__I_0_add_1503_14 (.CI(n50236), .I0(n2222), 
            .I1(VCC_net), .CO(n50237));
    SB_CARRY encoder0_position_30__I_0_add_967_7 (.CI(n49955), .I0(n1429), 
            .I1(GND_net), .CO(n49956));
    SB_LUT4 encoder0_position_30__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n50235), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_13 (.CI(n50235), .I0(n2223), 
            .I1(VCC_net), .CO(n50236));
    SB_LUT4 encoder0_position_30__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n50234), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28323_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5701), .I3(n15), .O(n42304));
    defparam i28323_4_lut.LUT_INIT = 16'hf535;
    SB_CARRY encoder0_position_30__I_0_add_1503_12 (.CI(n50234), .I0(n2224), 
            .I1(VCC_net), .CO(n50235));
    SB_LUT4 encoder0_position_30__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n49954), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15395_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n57425), .I3(GND_net), .O(n29471));   // verilog/coms.v(130[12] 305[6])
    defparam i15395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n50233), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_11 (.CI(n50233), .I0(n2225), 
            .I1(VCC_net), .CO(n50234));
    SB_LUT4 encoder0_position_30__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n50232), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n69709_bdd_4_lut (.I0(n69709), .I1(duty[8]), .I2(n4920), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n69709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i42497_3_lut (.I0(encoder0_position[28]), .I1(n58173), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42497_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1503_10 (.CI(n50232), .I0(n2226), 
            .I1(VCC_net), .CO(n50233));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n49779), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_6 (.CI(n49954), .I0(n1430), 
            .I1(GND_net), .CO(n49955));
    SB_LUT4 encoder0_position_30__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n50231), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_9 (.CI(n50231), .I0(n2227), 
            .I1(VCC_net), .CO(n50232));
    SB_LUT4 encoder0_position_30__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n50230), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n49953), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_8 (.CI(n50230), .I0(n2228), 
            .I1(VCC_net), .CO(n50231));
    SB_LUT4 encoder0_position_30__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n50229), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n49513), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_5 (.CI(n49953), .I0(n1431), 
            .I1(VCC_net), .CO(n49954));
    SB_CARRY encoder0_position_30__I_0_add_1503_7 (.CI(n50229), .I0(n2229), 
            .I1(GND_net), .CO(n50230));
    SB_LUT4 encoder0_position_30__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n50228), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_13 (.CI(n49521), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n49522));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n49778), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n49952), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n49778), .I0(GND_net), .I1(n2), 
            .CO(n49779));
    SB_CARRY encoder0_position_30__I_0_add_1503_6 (.CI(n50228), .I0(n2230), 
            .I1(GND_net), .CO(n50229));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n49777), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n50227), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11579_bdd_4_lut_53934 (.I0(n11579), .I1(current[7]), .I2(duty[10]), 
            .I3(n11577), .O(n69703));
    defparam n11579_bdd_4_lut_53934.LUT_INIT = 16'he4aa;
    SB_LUT4 n69703_bdd_4_lut (.I0(n69703), .I1(duty[7]), .I2(n4921), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n69703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11579_bdd_4_lut_53929 (.I0(n11579), .I1(current[6]), .I2(duty[9]), 
            .I3(n11577), .O(n69697));
    defparam n11579_bdd_4_lut_53929.LUT_INIT = 16'he4aa;
    SB_LUT4 n69697_bdd_4_lut (.I0(n69697), .I1(duty[6]), .I2(n4922), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n69697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11579_bdd_4_lut_53924 (.I0(n11579), .I1(current[5]), .I2(duty[8]), 
            .I3(n11577), .O(n69691));
    defparam n11579_bdd_4_lut_53924.LUT_INIT = 16'he4aa;
    SB_LUT4 n69691_bdd_4_lut (.I0(n69691), .I1(duty[5]), .I2(n4923), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n69691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53919 (.I0(n11579), .I1(current[4]), .I2(duty[7]), 
            .I3(n11577), .O(n69685));
    defparam n11579_bdd_4_lut_53919.LUT_INIT = 16'he4aa;
    SB_LUT4 n69685_bdd_4_lut (.I0(n69685), .I1(duty[4]), .I2(n4924), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n69685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226_adj_5804));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53914 (.I0(n11579), .I1(current[3]), .I2(duty[6]), 
            .I3(n11577), .O(n69679));
    defparam n11579_bdd_4_lut_53914.LUT_INIT = 16'he4aa;
    SB_LUT4 n69679_bdd_4_lut (.I0(n69679), .I1(duty[3]), .I2(n4925), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n69679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i837_3_lut (.I0(n1226_adj_5804), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53909 (.I0(n11579), .I1(current[2]), .I2(duty[5]), 
            .I3(n11577), .O(n69673));
    defparam n11579_bdd_4_lut_53909.LUT_INIT = 16'he4aa;
    SB_LUT4 n69673_bdd_4_lut (.I0(n69673), .I1(duty[2]), .I2(n4926), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n69673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53904 (.I0(n11579), .I1(current[1]), .I2(duty[4]), 
            .I3(n11577), .O(n69667));
    defparam n11579_bdd_4_lut_53904.LUT_INIT = 16'he4aa;
    SB_LUT4 n69667_bdd_4_lut (.I0(n69667), .I1(duty[1]), .I2(n4927), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n69667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53899 (.I0(n11579), .I1(current[0]), .I2(duty[3]), 
            .I3(n11577), .O(n69661));
    defparam n11579_bdd_4_lut_53899.LUT_INIT = 16'he4aa;
    SB_LUT4 n69661_bdd_4_lut (.I0(n69661), .I1(duty[0]), .I2(n4928), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n69661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_967_4 (.CI(n49952), .I0(n1432), 
            .I1(GND_net), .CO(n49953));
    SB_LUT4 encoder0_position_30__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n49951), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_3 (.CI(n49951), .I0(n1433), 
            .I1(VCC_net), .CO(n49952));
    SB_LUT4 encoder0_position_30__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_5 (.CI(n50227), .I0(n2231), 
            .I1(VCC_net), .CO(n50228));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n49777), .I0(GND_net), .I1(n14), 
            .CO(n49778));
    SB_LUT4 encoder0_position_30__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n50226), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n49951));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5688), 
            .I3(n49776), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_4 (.CI(n50226), .I0(n2232), 
            .I1(GND_net), .CO(n50227));
    SB_CARRY unary_minus_16_add_3_12 (.CI(n49776), .I0(GND_net), .I1(n15_adj_5688), 
            .CO(n49777));
    SB_LUT4 encoder0_position_30__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n50225), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_3 (.CI(n50225), .I0(n2233), 
            .I1(VCC_net), .CO(n50226));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5689), 
            .I3(n49775), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n50225));
    SB_LUT4 encoder0_position_30__I_0_add_1436_21_lut (.I0(GND_net), .I1(n2115), 
            .I2(VCC_net), .I3(n50224), .O(n2182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n49775), .I0(GND_net), .I1(n16_adj_5689), 
            .CO(n49776));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5690), 
            .I3(n49774), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n50223), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_20 (.CI(n50223), .I0(n2116), 
            .I1(VCC_net), .CO(n50224));
    SB_LUT4 encoder0_position_30__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n50222), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n49774), .I0(GND_net), .I1(n17_adj_5690), 
            .CO(n49775));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n49773), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_19 (.CI(n50222), .I0(n2117), 
            .I1(VCC_net), .CO(n50223));
    SB_LUT4 encoder0_position_30__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n50221), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_18 (.CI(n50221), .I0(n2118), 
            .I1(VCC_net), .CO(n50222));
    SB_LUT4 encoder0_position_30__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n50220), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n49773), .I0(GND_net), .I1(n18), 
            .CO(n49774));
    SB_CARRY encoder0_position_30__I_0_add_1436_17 (.CI(n50220), .I0(n2119), 
            .I1(VCC_net), .CO(n50221));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5691), 
            .I3(n49772), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n50219), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n49772), .I0(GND_net), .I1(n19_adj_5691), 
            .CO(n49773));
    SB_CARRY encoder0_position_30__I_0_add_1436_16 (.CI(n50219), .I0(n2120), 
            .I1(VCC_net), .CO(n50220));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5692), 
            .I3(n49771), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n49771), .I0(GND_net), .I1(n20_adj_5692), 
            .CO(n49772));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5693), 
            .I3(n49770), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n50218), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_15 (.CI(n50218), .I0(n2121), 
            .I1(VCC_net), .CO(n50219));
    SB_LUT4 encoder0_position_30__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n50217), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n49770), .I0(GND_net), .I1(n21_adj_5693), 
            .CO(n49771));
    SB_LUT4 i42610_2_lut_3_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n57410), 
            .I2(n8_adj_5801), .I3(GND_net), .O(n58294));
    defparam i42610_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_30__I_0_add_1436_14 (.CI(n50217), .I0(n2122), 
            .I1(VCC_net), .CO(n50218));
    SB_LUT4 encoder0_position_30__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n50216), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5694), 
            .I3(n49769), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_13 (.CI(n50216), .I0(n2123), 
            .I1(VCC_net), .CO(n50217));
    SB_LUT4 encoder0_position_30__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n50215), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_12 (.CI(n50215), .I0(n2124), 
            .I1(VCC_net), .CO(n50216));
    SB_LUT4 encoder0_position_30__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n50214), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_11 (.CI(n50214), .I0(n2125), 
            .I1(VCC_net), .CO(n50215));
    SB_LUT4 encoder0_position_30__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n50213), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n49769), .I0(GND_net), .I1(n22_adj_5694), 
            .CO(n49770));
    SB_CARRY encoder0_position_30__I_0_add_1436_10 (.CI(n50213), .I0(n2126), 
            .I1(VCC_net), .CO(n50214));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5695), 
            .I3(n49768), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n50212), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_9 (.CI(n50212), .I0(n2127), 
            .I1(VCC_net), .CO(n50213));
    SB_LUT4 encoder0_position_30__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n50211), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_8 (.CI(n50211), .I0(n2128), 
            .I1(VCC_net), .CO(n50212));
    SB_LUT4 i1_4_lut_adj_2064 (.I0(n1229_adj_5807), .I1(n43591), .I2(n1230_adj_5808), 
            .I3(n1231_adj_5809), .O(n59015));
    defparam i1_4_lut_adj_2064.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n50210), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_7 (.CI(n50210), .I0(n2129), 
            .I1(GND_net), .CO(n50211));
    SB_CARRY unary_minus_16_add_3_4 (.CI(n49768), .I0(GND_net), .I1(n23_adj_5695), 
            .CO(n49769));
    SB_LUT4 encoder0_position_30__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n50209), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_13_lut (.I0(n69303), .I1(n1323), 
            .I2(VCC_net), .I3(n49935), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1436_6 (.CI(n50209), .I0(n2130), 
            .I1(GND_net), .CO(n50210));
    SB_LUT4 encoder0_position_30__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n49934), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n50208), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_5 (.CI(n50208), .I0(n2131), 
            .I1(VCC_net), .CO(n50209));
    SB_LUT4 encoder0_position_30__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n50207), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_12 (.CI(n49934), .I0(n1324), 
            .I1(VCC_net), .CO(n49935));
    SB_CARRY encoder0_position_30__I_0_add_1436_4 (.CI(n50207), .I0(n2132), 
            .I1(GND_net), .CO(n50208));
    SB_LUT4 encoder0_position_30__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n49933), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n50206), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_3 (.CI(n50206), .I0(n2133), 
            .I1(VCC_net), .CO(n50207));
    SB_LUT4 encoder0_position_30__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n50206));
    SB_LUT4 encoder0_position_30__I_0_add_1369_20_lut (.I0(n69092), .I1(n2016), 
            .I2(VCC_net), .I3(n50205), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n50204), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_19 (.CI(n50204), .I0(n2017), 
            .I1(VCC_net), .CO(n50205));
    SB_LUT4 encoder0_position_30__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n50203), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_18 (.CI(n50203), .I0(n2018), 
            .I1(VCC_net), .CO(n50204));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5696), 
            .I3(n49767), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n50202), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_11 (.CI(n49933), .I0(n1325), 
            .I1(VCC_net), .CO(n49934));
    SB_CARRY encoder0_position_30__I_0_add_1369_17 (.CI(n50202), .I0(n2019), 
            .I1(VCC_net), .CO(n50203));
    SB_CARRY unary_minus_16_add_3_3 (.CI(n49767), .I0(GND_net), .I1(n24_adj_5696), 
            .CO(n49768));
    SB_LUT4 encoder0_position_30__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n49932), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n50201), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_16 (.CI(n50201), .I0(n2020), 
            .I1(VCC_net), .CO(n50202));
    SB_LUT4 encoder0_position_30__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n50200), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n43450), .I1(GND_net), .I2(n25_adj_5697), 
            .I3(VCC_net), .O(n65589)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_900_10 (.CI(n49932), .I0(n1326), 
            .I1(VCC_net), .CO(n49933));
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5697), 
            .CO(n49767));
    SB_LUT4 encoder0_position_30__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n49931), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_15 (.CI(n50200), .I0(n2021), 
            .I1(VCC_net), .CO(n50201));
    SB_LUT4 encoder0_position_30__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n50199), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_14 (.CI(n50199), .I0(n2022), 
            .I1(VCC_net), .CO(n50200));
    SB_LUT4 encoder0_position_30__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n50198), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_9 (.CI(n49931), .I0(n1327), 
            .I1(VCC_net), .CO(n49932));
    SB_CARRY encoder0_position_30__I_0_add_1369_13 (.CI(n50198), .I0(n2023), 
            .I1(VCC_net), .CO(n50199));
    SB_LUT4 encoder0_position_30__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n50197), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5773), .I3(n49766), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_12 (.CI(n50197), .I0(n2024), 
            .I1(VCC_net), .CO(n50198));
    SB_LUT4 encoder0_position_30__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n50196), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5772), .I3(n49765), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n49930), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_11 (.CI(n50196), .I0(n2025), 
            .I1(VCC_net), .CO(n50197));
    SB_LUT4 encoder0_position_30__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n50195), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_10 (.CI(n50195), .I0(n2026), 
            .I1(VCC_net), .CO(n50196));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n49765), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5772), .CO(n49766));
    SB_LUT4 encoder0_position_30__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n50194), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5771), .I3(n49764), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_8 (.CI(n49930), .I0(n1328), 
            .I1(VCC_net), .CO(n49931));
    SB_LUT4 encoder0_position_30__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n49929), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_9 (.CI(n50194), .I0(n2027), 
            .I1(VCC_net), .CO(n50195));
    SB_CARRY encoder0_position_30__I_0_add_900_7 (.CI(n49929), .I0(n1329), 
            .I1(GND_net), .CO(n49930));
    SB_LUT4 encoder0_position_30__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n50193), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_8 (.CI(n50193), .I0(n2028), 
            .I1(VCC_net), .CO(n50194));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n49764), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5771), .CO(n49765));
    SB_LUT4 encoder0_position_30__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n50192), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n49928), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_6 (.CI(n49928), .I0(n1330), 
            .I1(GND_net), .CO(n49929));
    SB_LUT4 encoder0_position_30__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n49927), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_5 (.CI(n49927), .I0(n1331), 
            .I1(VCC_net), .CO(n49928));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5799), .I3(n49763), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1172_3_lut (.I0(n1721), .I1(n1788_adj_5813), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1369_7 (.CI(n50192), .I0(n2029), 
            .I1(GND_net), .CO(n50193));
    SB_LUT4 encoder0_position_30__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n50191), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut_adj_2065 (.I0(\data_out_frame[21] [0]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5894));
    defparam i1_2_lut_adj_2065.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n25_adj_5812), .I1(n53095), .I2(n57836), .I3(n6_adj_5894), 
            .O(n52011));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n49926), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_6 (.CI(n50191), .I0(n2030), 
            .I1(GND_net), .CO(n50192));
    SB_CARRY encoder0_position_30__I_0_add_900_4 (.CI(n49926), .I0(n1332), 
            .I1(GND_net), .CO(n49927));
    SB_LUT4 encoder0_position_30__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n49925), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_3 (.CI(n49925), .I0(n1333), 
            .I1(VCC_net), .CO(n49926));
    SB_LUT4 encoder0_position_30__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n50190), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_5 (.CI(n50190), .I0(n2031), 
            .I1(VCC_net), .CO(n50191));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n49763), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5799), .CO(n49764));
    SB_LUT4 encoder0_position_30__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n50189), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_4 (.CI(n50189), .I0(n2032), 
            .I1(GND_net), .CO(n50190));
    SB_LUT4 encoder0_position_30__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n50188), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_2_lut (.I0(GND_net), .I1(n524), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_2 (.CI(VCC_net), .I0(n524), 
            .I1(GND_net), .CO(n49925));
    SB_CARRY encoder0_position_30__I_0_add_1369_3 (.CI(n50188), .I0(n2033), 
            .I1(VCC_net), .CO(n50189));
    SB_LUT4 encoder0_position_30__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n50188));
    SB_LUT4 i52939_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42725), .I3(GND_net), .O(n27728));
    defparam i52939_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i50306_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n65611));
    defparam i50306_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i28877_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42725), .I3(GND_net), .O(n42845));
    defparam i28877_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5796), .I3(n49762), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n49762), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5796), .CO(n49763));
    SB_LUT4 i6565_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6565_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i6567_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6567_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5795), .I3(n49761), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n49761), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5795), .CO(n49762));
    SB_LUT4 i6569_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i6569_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i6571_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i6571_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5741));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5737));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5794), .I3(n49760), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5739));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n49760), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5794), .CO(n49761));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5793), .I3(n49759), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n49759), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5793), .CO(n49760));
    SB_LUT4 i23916_3_lut_4_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30383));
    defparam i23916_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16306_3_lut_4_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30382));   // verilog/coms.v(130[12] 305[6])
    defparam i16306_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16304_3_lut_4_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30380));   // verilog/coms.v(130[12] 305[6])
    defparam i16304_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5792), .I3(n49758), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut_adj_2066 (.I0(n260), .I1(n62792), .I2(duty[23]), 
            .I3(n22_adj_5911), .O(n11577));
    defparam i1_4_lut_4_lut_adj_2066.LUT_INIT = 16'h1505;
    SB_LUT4 i1_2_lut_adj_2067 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5812));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_2067.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n49758), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5792), .CO(n49759));
    SB_LUT4 encoder0_position_30__I_0_add_1302_19_lut (.I0(n69088), .I1(n1917), 
            .I2(VCC_net), .I3(n50165), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n50164), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_18 (.CI(n50164), .I0(n1918), 
            .I1(VCC_net), .CO(n50165));
    SB_LUT4 encoder0_position_30__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n50163), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_17 (.CI(n50163), .I0(n1919), 
            .I1(VCC_net), .CO(n50164));
    SB_LUT4 encoder0_position_30__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n50162), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_16 (.CI(n50162), .I0(n1920), 
            .I1(VCC_net), .CO(n50163));
    SB_LUT4 encoder0_position_30__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n50161), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_15 (.CI(n50161), .I0(n1921), 
            .I1(VCC_net), .CO(n50162));
    SB_LUT4 encoder0_position_30__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n50160), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5791), .I3(n49757), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n49757), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5791), .CO(n49758));
    SB_CARRY encoder0_position_30__I_0_add_1302_14 (.CI(n50160), .I0(n1922), 
            .I1(VCC_net), .CO(n50161));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5780), .I3(n49756), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16302_3_lut_4_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30378));   // verilog/coms.v(130[12] 305[6])
    defparam i16302_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n50159), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n3470), .I2(n161), 
            .I3(\FRAME_MATCHER.i [4]), .O(n91));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_CARRY encoder0_position_30__I_0_add_1302_13 (.CI(n50159), .I0(n1923), 
            .I1(VCC_net), .CO(n50160));
    SB_LUT4 i15444_3_lut_4_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(reset), .I3(n105), .O(n29520));   // verilog/coms.v(130[12] 305[6])
    defparam i15444_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15447_3_lut_4_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(reset), .I3(n105), .O(n29523));   // verilog/coms.v(130[12] 305[6])
    defparam i15447_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15450_3_lut_4_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(reset), .I3(n105), .O(n29526));   // verilog/coms.v(130[12] 305[6])
    defparam i15450_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15454_3_lut_4_lut (.I0(\data_in_frame[16] [6]), .I1(rx_data[6]), 
            .I2(reset), .I3(n105), .O(n29530));   // verilog/coms.v(130[12] 305[6])
    defparam i15454_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_30__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n50158), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_12 (.CI(n50158), .I0(n1924), 
            .I1(VCC_net), .CO(n50159));
    SB_LUT4 encoder0_position_30__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n50157), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n49756), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5780), .CO(n49757));
    SB_CARRY encoder0_position_30__I_0_add_1302_11 (.CI(n50157), .I0(n1925), 
            .I1(VCC_net), .CO(n50158));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n50156), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_10 (.CI(n50156), .I0(n1926), 
            .I1(VCC_net), .CO(n50157));
    SB_LUT4 i11_2_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n25848));   // verilog/coms.v(100[12:26])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n50155), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_9 (.CI(n50155), .I0(n1927), 
            .I1(VCC_net), .CO(n50156));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5779), .I3(n49755), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42606_2_lut_3_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n57410), 
            .I2(n8_adj_5774), .I3(GND_net), .O(n58290));
    defparam i42606_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15799_3_lut_4_lut (.I0(deadband[6]), .I1(\data_in_frame[16] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29875));   // verilog/coms.v(130[12] 305[6])
    defparam i15799_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15798_3_lut_4_lut (.I0(deadband[7]), .I1(\data_in_frame[16] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29874));   // verilog/coms.v(130[12] 305[6])
    defparam i15798_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15797_3_lut_4_lut (.I0(deadband[8]), .I1(\data_in_frame[15] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29873));   // verilog/coms.v(130[12] 305[6])
    defparam i15797_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n50154), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15796_3_lut_4_lut (.I0(deadband[9]), .I1(\data_in_frame[15] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29872));   // verilog/coms.v(130[12] 305[6])
    defparam i15796_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n49755), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5779), .CO(n49756));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5778), .I3(n49754), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_8 (.CI(n50154), .I0(n1928), 
            .I1(VCC_net), .CO(n50155));
    SB_LUT4 i50820_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n66548));
    defparam i50820_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_30__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n50153), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_7 (.CI(n50153), .I0(n1929), 
            .I1(GND_net), .CO(n50154));
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_833_12_lut (.I0(GND_net), .I1(n1224_adj_5802), 
            .I2(VCC_net), .I3(n49903), .O(n1291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15795_3_lut_4_lut (.I0(deadband[10]), .I1(\data_in_frame[15] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29871));   // verilog/coms.v(130[12] 305[6])
    defparam i15795_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225_adj_5803), 
            .I2(VCC_net), .I3(n49902), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_11 (.CI(n49902), .I0(n1225_adj_5803), 
            .I1(VCC_net), .CO(n49903));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n49754), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5778), .CO(n49755));
    SB_LUT4 encoder0_position_30__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226_adj_5804), 
            .I2(VCC_net), .I3(n49901), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5777), .I3(n49753), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n50152), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_6 (.CI(n50152), .I0(n1930), 
            .I1(GND_net), .CO(n50153));
    SB_LUT4 encoder0_position_30__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n50151), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1174_3_lut (.I0(n1723), .I1(n1790_adj_5814), 
            .I2(n1752), .I3(GND_net), .O(n1822_adj_5818));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1241_3_lut (.I0(n1822_adj_5818), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n49753), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5777), .CO(n49754));
    SB_CARRY encoder0_position_30__I_0_add_833_10 (.CI(n49901), .I0(n1226_adj_5804), 
            .I1(VCC_net), .CO(n49902));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5775), .I3(n49752), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227_adj_5805), 
            .I2(VCC_net), .I3(n49900), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_5 (.CI(n50151), .I0(n1931), 
            .I1(VCC_net), .CO(n50152));
    SB_LUT4 i15794_3_lut_4_lut (.I0(deadband[11]), .I1(\data_in_frame[15] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29870));   // verilog/coms.v(130[12] 305[6])
    defparam i15794_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n50150), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15793_3_lut_4_lut (.I0(deadband[12]), .I1(\data_in_frame[15] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29869));   // verilog/coms.v(130[12] 305[6])
    defparam i15793_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_833_9 (.CI(n49900), .I0(n1227_adj_5805), 
            .I1(VCC_net), .CO(n49901));
    SB_LUT4 i15792_3_lut_4_lut (.I0(deadband[13]), .I1(\data_in_frame[15] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29868));   // verilog/coms.v(130[12] 305[6])
    defparam i15792_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15791_3_lut_4_lut (.I0(deadband[14]), .I1(\data_in_frame[15] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29867));   // verilog/coms.v(130[12] 305[6])
    defparam i15791_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15790_3_lut_4_lut (.I0(deadband[15]), .I1(\data_in_frame[15] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29866));   // verilog/coms.v(130[12] 305[6])
    defparam i15790_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_1302_4 (.CI(n50150), .I0(n1932), 
            .I1(GND_net), .CO(n50151));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n49752), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5775), .CO(n49753));
    SB_LUT4 encoder0_position_30__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n50149), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_3 (.CI(n50149), .I0(n1933), 
            .I1(VCC_net), .CO(n50150));
    SB_LUT4 i15789_3_lut_4_lut (.I0(deadband[16]), .I1(\data_in_frame[14] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29865));   // verilog/coms.v(130[12] 305[6])
    defparam i15789_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15788_3_lut_4_lut (.I0(deadband[17]), .I1(\data_in_frame[14] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29864));   // verilog/coms.v(130[12] 305[6])
    defparam i15788_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15787_3_lut_4_lut (.I0(deadband[18]), .I1(\data_in_frame[14] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29863));   // verilog/coms.v(130[12] 305[6])
    defparam i15787_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15786_3_lut_4_lut (.I0(deadband[19]), .I1(\data_in_frame[14] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29862));   // verilog/coms.v(130[12] 305[6])
    defparam i15786_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228_adj_5806), 
            .I2(VCC_net), .I3(n49899), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15785_3_lut_4_lut (.I0(deadband[20]), .I1(\data_in_frame[14] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29861));   // verilog/coms.v(130[12] 305[6])
    defparam i15785_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15784_3_lut_4_lut (.I0(deadband[21]), .I1(\data_in_frame[14] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29860));   // verilog/coms.v(130[12] 305[6])
    defparam i15784_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n50149));
    SB_LUT4 i15783_3_lut_4_lut (.I0(deadband[22]), .I1(\data_in_frame[14] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29859));   // verilog/coms.v(130[12] 305[6])
    defparam i15783_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_833_8 (.CI(n49899), .I0(n1228_adj_5806), 
            .I1(VCC_net), .CO(n49900));
    SB_LUT4 i15782_3_lut_4_lut (.I0(deadband[23]), .I1(\data_in_frame[14] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29858));   // verilog/coms.v(130[12] 305[6])
    defparam i15782_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i42608_2_lut_3_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n57410), 
            .I2(n8_adj_5757), .I3(GND_net), .O(n58292));
    defparam i42608_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15781_3_lut_4_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29857));   // verilog/coms.v(130[12] 305[6])
    defparam i15781_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15780_3_lut_4_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29856));   // verilog/coms.v(130[12] 305[6])
    defparam i15780_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15779_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29855));   // verilog/coms.v(130[12] 305[6])
    defparam i15779_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5770), .I3(n49751), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n49751), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5770), .CO(n49752));
    SB_LUT4 i15778_3_lut_4_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29854));   // verilog/coms.v(130[12] 305[6])
    defparam i15778_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFF read_197 (.Q(state_7__N_3916[0]), .C(clk16MHz), .D(n60507));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i15777_3_lut_4_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29853));   // verilog/coms.v(130[12] 305[6])
    defparam i15777_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15776_3_lut_4_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29852));   // verilog/coms.v(130[12] 305[6])
    defparam i15776_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15775_3_lut_4_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29851));   // verilog/coms.v(130[12] 305[6])
    defparam i15775_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229_adj_5807), 
            .I2(GND_net), .I3(n49898), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_7 (.CI(n49898), .I0(n1229_adj_5807), 
            .I1(GND_net), .CO(n49899));
    SB_LUT4 encoder0_position_30__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230_adj_5808), 
            .I2(GND_net), .I3(n49897), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5769), .I3(n49750), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n49750), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5769), .CO(n49751));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5768), .I3(n49749), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n49749), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5768), .CO(n49750));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n49748), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_4310_i11_3_lut (.I0(encoder0_position[10]), .I1(n22_adj_5709), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53881 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n69637));
    defparam byte_transmit_counter_0__bdd_4_lut_53881.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_adj_2068 (.I0(n1225_adj_5803), .I1(n1226_adj_5804), 
            .I2(n1227_adj_5805), .I3(GND_net), .O(n61714));
    defparam i1_3_lut_adj_2068.LUT_INIT = 16'hfefe;
    SB_LUT4 i53640_4_lut (.I0(n1224_adj_5802), .I1(n61714), .I2(n1228_adj_5806), 
            .I3(n59015), .O(n1257));
    defparam i53640_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n69637_bdd_4_lut (.I0(n69637), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n69640));
    defparam n69637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5679));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50780_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n66508));
    defparam i50780_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15774_3_lut_4_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29850));   // verilog/coms.v(130[12] 305[6])
    defparam i15774_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227_adj_5805));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29612_3_lut (.I0(n524), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n43587));
    defparam i29612_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2069 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n61680));
    defparam i1_4_lut_adj_2069.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2070 (.I0(n1329), .I1(n43587), .I2(n1330), .I3(n1331), 
            .O(n59013));
    defparam i1_4_lut_adj_2070.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53590_4_lut (.I0(n59013), .I1(n1323), .I2(n1324), .I3(n61680), 
            .O(n1356));
    defparam i53590_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n49748), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n49749));
    SB_CARRY encoder0_position_30__I_0_add_833_6 (.CI(n49897), .I0(n1230_adj_5808), 
            .I1(GND_net), .CO(n49898));
    SB_LUT4 encoder0_position_30__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231_adj_5809), 
            .I2(VCC_net), .I3(n49896), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_5 (.CI(n49896), .I0(n1231_adj_5809), 
            .I1(VCC_net), .CO(n49897));
    SB_LUT4 i15773_3_lut_4_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29849));   // verilog/coms.v(130[12] 305[6])
    defparam i15773_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i838_3_lut (.I0(n1227_adj_5805), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29608_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n43583));
    defparam i29608_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_2_lut_adj_2071 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n61720));
    defparam i1_2_lut_adj_2071.LUT_INIT = 16'heeee;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2072 (.I0(n1429), .I1(n43583), .I2(n1430), .I3(n1431), 
            .O(n59026));
    defparam i1_4_lut_adj_2072.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2073 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n61720), 
            .O(n61726));
    defparam i1_4_lut_adj_2073.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i53625_4_lut (.I0(n1423), .I1(n1422), .I2(n61726), .I3(n59026), 
            .O(n1455));
    defparam i53625_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_2_lut_adj_2074 (.I0(n1527), .I1(n1528), .I2(GND_net), .I3(GND_net), 
            .O(n61406));
    defparam i1_2_lut_adj_2074.LUT_INIT = 16'heeee;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29676_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n43651));
    defparam i29676_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2075 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n61406), 
            .O(n61412));
    defparam i1_4_lut_adj_2075.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2076 (.I0(n1529), .I1(n61412), .I2(n43651), .I3(n1530), 
            .O(n61414));
    defparam i1_4_lut_adj_2076.LUT_INIT = 16'heccc;
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i53608_4_lut (.I0(n1522), .I1(n1521), .I2(n61414), .I3(n1523), 
            .O(n1554));
    defparam i53608_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i15772_3_lut_4_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29848));   // verilog/coms.v(130[12] 305[6])
    defparam i15772_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232_adj_5810), 
            .I2(GND_net), .I3(n49895), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22520_3_lut_4_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29847));
    defparam i22520_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i29600_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n43575));
    defparam i29600_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_2077 (.I0(n1629), .I1(n43575), .I2(n1630), .I3(n1631), 
            .O(n59034));
    defparam i1_4_lut_adj_2077.LUT_INIT = 16'ha080;
    SB_LUT4 i22521_3_lut_4_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29846));
    defparam i22521_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15769_3_lut_4_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29845));   // verilog/coms.v(130[12] 305[6])
    defparam i15769_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15768_3_lut_4_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29844));   // verilog/coms.v(130[12] 305[6])
    defparam i15768_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15767_3_lut_4_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29843));   // verilog/coms.v(130[12] 305[6])
    defparam i15767_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15766_3_lut_4_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29842));   // verilog/coms.v(130[12] 305[6])
    defparam i15766_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27728), 
            .D(n1238), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 mux_4310_i21_3_lut (.I0(encoder0_position[20]), .I1(n12), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_2078 (.I0(\data_in_frame[22] [5]), .I1(n8_adj_5801), 
            .I2(n43396), .I3(n57340), .O(n56402));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2078.LUT_INIT = 16'ha3a0;
    SB_LUT4 mux_4310_i15_3_lut (.I0(encoder0_position[14]), .I1(n18_adj_5713), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27728), 
            .D(n1237), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27728), 
            .D(n1236), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27728), 
            .D(n1235), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27728), 
            .D(n1234), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27728), 
            .D(n1233), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27728), 
            .D(n1232), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27728), 
            .D(n1231), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27728), 
            .D(n1230), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27728), 
            .D(n1229), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27728), 
            .D(n1228), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27728), 
            .D(n1227), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27728), 
            .D(n1226), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27728), 
            .D(n1225), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27728), 
            .D(n1224), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27728), 
            .D(n1223), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27728), 
            .D(n1222), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27728), 
            .D(n1221), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27728), 
            .D(n1220), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n58169));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n49747), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i845_3_lut (.I0(n523), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5855), .I3(n50995), .O(n2_adj_5731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5856), .I3(n50994), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_4 (.CI(n49895), .I0(n1232_adj_5810), 
            .I1(GND_net), .CO(n49896));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_32 (.CI(n50994), 
            .I0(GND_net), .I1(n3_adj_5856), .CO(n50995));
    SB_LUT4 encoder0_position_30__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233_adj_5811), 
            .I2(VCC_net), .I3(n49894), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n49747), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n49748));
    SB_CARRY encoder0_position_30__I_0_add_833_3 (.CI(n49894), .I0(n1233_adj_5811), 
            .I1(VCC_net), .CO(n49895));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5857), .I3(n50993), .O(n4_adj_5730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_31 (.CI(n50993), 
            .I0(GND_net), .I1(n4_adj_5857), .CO(n50994));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5858), .I3(n50992), .O(n5_adj_5725)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_30 (.CI(n50992), 
            .I0(GND_net), .I1(n5_adj_5858), .CO(n50993));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5859), .I3(n50991), .O(n6_adj_5723)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_29 (.CI(n50991), 
            .I0(GND_net), .I1(n6_adj_5859), .CO(n50992));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5860), .I3(n50990), .O(n7_adj_5722)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2079 (.I0(n1624), .I1(n1626), .I2(n1627), .I3(n1628), 
            .O(n61740));
    defparam i1_4_lut_adj_2079.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_28 (.CI(n50990), 
            .I0(GND_net), .I1(n7_adj_5860), .CO(n50991));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5861), .I3(n50989), .O(n8_adj_5721)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_27 (.CI(n50989), 
            .I0(GND_net), .I1(n8_adj_5861), .CO(n50990));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5862), .I3(n50988), .O(n9_adj_5720)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_26 (.CI(n50988), 
            .I0(GND_net), .I1(n9_adj_5862), .CO(n50989));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5863), .I3(n50987), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_25 (.CI(n50987), 
            .I0(GND_net), .I1(n10_adj_5863), .CO(n50988));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5864), .I3(n50986), .O(n11_adj_5719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_24 (.CI(n50986), 
            .I0(GND_net), .I1(n11_adj_5864), .CO(n50987));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5865), .I3(n50985), .O(n12)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_23 (.CI(n50985), 
            .I0(GND_net), .I1(n12_adj_5865), .CO(n50986));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5866), .I3(n50984), .O(n13_adj_5718)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_22 (.CI(n50984), 
            .I0(GND_net), .I1(n13_adj_5866), .CO(n50985));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5867), .I3(n50983), .O(n14_adj_5717)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n49746), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n49746), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n49747));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_21 (.CI(n50983), 
            .I0(GND_net), .I1(n14_adj_5867), .CO(n50984));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5868), .I3(n50982), .O(n15_adj_5716)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_20 (.CI(n50982), 
            .I0(GND_net), .I1(n15_adj_5868), .CO(n50983));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5869), .I3(n50981), .O(n16_adj_5715)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_2_lut (.I0(GND_net), .I1(n523), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_19 (.CI(n50981), 
            .I0(GND_net), .I1(n16_adj_5869), .CO(n50982));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5870), .I3(n50980), .O(n17_adj_5714)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_18 (.CI(n50980), 
            .I0(GND_net), .I1(n17_adj_5870), .CO(n50981));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5871), .I3(n50979), .O(n18_adj_5713)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_17 (.CI(n50979), 
            .I0(GND_net), .I1(n18_adj_5871), .CO(n50980));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5872), .I3(n50978), .O(n19_adj_5712)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_16 (.CI(n50978), 
            .I0(GND_net), .I1(n19_adj_5872), .CO(n50979));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5873), .I3(n50977), .O(n20_adj_5711)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_15 (.CI(n50977), 
            .I0(GND_net), .I1(n20_adj_5873), .CO(n50978));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5874), .I3(n50976), .O(n21_adj_5710)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_14 (.CI(n50976), 
            .I0(GND_net), .I1(n21_adj_5874), .CO(n50977));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5875), .I3(n50975), .O(n22_adj_5709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_13 (.CI(n50975), 
            .I0(GND_net), .I1(n22_adj_5875), .CO(n50976));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5876), .I3(n50974), .O(n23_adj_5708)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_12 (.CI(n50974), 
            .I0(GND_net), .I1(n23_adj_5876), .CO(n50975));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5877), .I3(n50973), .O(n24_adj_5707)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_11 (.CI(n50973), 
            .I0(GND_net), .I1(n24_adj_5877), .CO(n50974));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5878), .I3(n50972), .O(n25_adj_5706)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_10 (.CI(n50972), 
            .I0(GND_net), .I1(n25_adj_5878), .CO(n50973));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5879), .I3(n50971), .O(n26_adj_5705)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_9 (.CI(n50971), 
            .I0(GND_net), .I1(n26_adj_5879), .CO(n50972));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5880), .I3(n50970), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_8 (.CI(n50970), 
            .I0(GND_net), .I1(n27_adj_5880), .CO(n50971));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5881), .I3(n50969), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_7 (.CI(n50969), 
            .I0(GND_net), .I1(n28_adj_5881), .CO(n50970));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5882), .I3(n50968), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_6 (.CI(n50968), 
            .I0(GND_net), .I1(n29_adj_5882), .CO(n50969));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5883), .I3(n50967), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_5 (.CI(n50967), 
            .I0(GND_net), .I1(n30_adj_5883), .CO(n50968));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5884), .I3(n50966), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_4 (.CI(n50966), 
            .I0(GND_net), .I1(n31_adj_5884), .CO(n50967));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5885), .I3(n50965), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_3 (.CI(n50965), 
            .I0(GND_net), .I1(n32_adj_5885), .CO(n50966));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n50965));
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFESR dti_counter_1937__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n27810), 
            .D(n44), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n27810), 
            .D(n43_adj_5845), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n27810), 
            .D(n42), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n27810), 
            .D(n41), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n27810), 
            .D(n40), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n27810), 
            .D(n39), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n27810), 
            .D(n38_adj_5844), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5885));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2080 (.I0(n1623), .I1(n1621), .I2(n59034), .I3(n1625), 
            .O(n60222));
    defparam i1_4_lut_adj_2080.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5884));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5883));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_833_2 (.CI(VCC_net), .I0(n523), 
            .I1(GND_net), .CO(n49894));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5882));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5881));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n49745), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dti_counter_1937__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n27810), 
            .D(n45_adj_5846), .R(n29192));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5880));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n49745), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n49746));
    SB_LUT4 i53500_4_lut (.I0(n1620), .I1(n60222), .I2(n1622), .I3(n61740), 
            .O(n1653));
    defparam i53500_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i22868_3_lut_4_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29841));
    defparam i22868_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5879));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5878));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5877));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5876));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5875));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2081 (.I0(n1728), .I1(n1726), .I2(n1727), .I3(GND_net), 
            .O(n61390));
    defparam i1_3_lut_adj_2081.LUT_INIT = 16'hfefe;
    SB_LUT4 i29620_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n43595));
    defparam i29620_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2082 (.I0(n1723), .I1(n1724), .I2(n61390), .I3(n1725), 
            .O(n61396));
    defparam i1_4_lut_adj_2082.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2083 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n61746));
    defparam i1_2_lut_adj_2083.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_2084 (.I0(n61746), .I1(n1722), .I2(n61396), .I3(n43595), 
            .O(n61400));
    defparam i1_4_lut_adj_2084.LUT_INIT = 16'hfefc;
    SB_LUT4 i53481_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n61400), 
            .O(n1752));
    defparam i53481_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5874));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2085 (.I0(n1825), .I1(n1826), .I2(n1828), .I3(n1827), 
            .O(n61758));
    defparam i1_4_lut_adj_2085.LUT_INIT = 16'hfffe;
    SB_LUT4 i29692_4_lut (.I0(n943), .I1(n1831), .I2(n1832), .I3(n1833), 
            .O(n43667));
    defparam i29692_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5873));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5872));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_2086 (.I0(n1823), .I1(n1824_adj_5819), .I2(n61758), 
            .I3(GND_net), .O(n61762));
    defparam i1_3_lut_adj_2086.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_2087 (.I0(n1820), .I1(n1821), .I2(n1822_adj_5818), 
            .I3(GND_net), .O(n61768));
    defparam i1_3_lut_adj_2087.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2088 (.I0(n1829), .I1(n61762), .I2(n43667), .I3(n1830), 
            .O(n61764));
    defparam i1_4_lut_adj_2088.LUT_INIT = 16'heccc;
    SB_LUT4 i53459_4_lut (.I0(n1818), .I1(n61764), .I2(n61768), .I3(n1819), 
            .O(n1851));
    defparam i53459_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2089 (.I0(n1926), .I1(n1928), .I2(n1925), .I3(n1927), 
            .O(n61370));
    defparam i1_4_lut_adj_2089.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29537_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n43511));
    defparam i29537_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2090 (.I0(n1922), .I1(n1923), .I2(n61370), .I3(n1924), 
            .O(n61376));
    defparam i1_4_lut_adj_2090.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2091 (.I0(n1929), .I1(n43511), .I2(n1930), .I3(n1931), 
            .O(n59056));
    defparam i1_4_lut_adj_2091.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2092 (.I0(n1920), .I1(n59056), .I2(n1921), .I3(n61376), 
            .O(n61382));
    defparam i1_4_lut_adj_2092.LUT_INIT = 16'hfffe;
    SB_LUT4 i53363_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n61382), 
            .O(n1950));
    defparam i53363_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2093 (.I0(n2024), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n61792));
    defparam i1_2_lut_adj_2093.LUT_INIT = 16'heeee;
    SB_LUT4 i29630_4_lut (.I0(n945), .I1(n2031), .I2(n2032), .I3(n2033), 
            .O(n43605));
    defparam i29630_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 mux_4310_i16_3_lut (.I0(encoder0_position[15]), .I1(n17_adj_5714), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1180_3_lut (.I0(n1729), .I1(n1796_adj_5817), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2094 (.I0(n2021), .I1(n2027), .I2(n61792), .I3(n2025), 
            .O(n61798));
    defparam i1_4_lut_adj_2094.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2095 (.I0(n2029), .I1(n61798), .I2(n43605), .I3(n2030), 
            .O(n61800));
    defparam i1_4_lut_adj_2095.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_30__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5871));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5870));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_2096 (.I0(n2022), .I1(n2023), .I2(n2028), .I3(GND_net), 
            .O(n61874));
    defparam i1_3_lut_adj_2096.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2097 (.I0(n61874), .I1(n2019), .I2(n61800), .I3(n2020), 
            .O(n61804));
    defparam i1_4_lut_adj_2097.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53386_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n61804), 
            .O(n2049));
    defparam i53386_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i17_3_lut (.I0(encoder0_position[16]), .I1(n16_adj_5715), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22830_3_lut_4_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29840));
    defparam i22830_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5869));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5868));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42500_3_lut (.I0(n6_adj_5723), .I1(n7454), .I2(n58170), .I3(GND_net), 
            .O(n58177));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42500_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n55644));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i42501_3_lut (.I0(encoder0_position[26]), .I1(n58177), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22799_3_lut_4_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29839));
    defparam i22799_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30519));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5867));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5866));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5865));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5864));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_1937_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n50767), .O(n38_adj_5844)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_1937_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n50766), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_8 (.CI(n50766), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n50767));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n49744), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n49744), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n49745));
    SB_LUT4 encoder0_position_30__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228_adj_5806));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_1937_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n50765), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_7 (.CI(n50765), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n50766));
    SB_LUT4 dti_counter_1937_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n50764), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_6 (.CI(n50764), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n50765));
    SB_LUT4 dti_counter_1937_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n50763), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_5 (.CI(n50763), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n50764));
    SB_LUT4 dti_counter_1937_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n50762), .O(n43_adj_5845)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i839_3_lut (.I0(n1228_adj_5806), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_1937_add_4_4 (.CI(n50762), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n50763));
    SB_LUT4 dti_counter_1937_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n50761), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_3 (.CI(n50761), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n50762));
    SB_LUT4 dti_counter_1937_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45_adj_5846)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n50761));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5863));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5862));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5861));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5860));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i27765_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5701), .I3(n15), .O(n41755));
    defparam i27765_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 mux_4310_i18_3_lut (.I0(encoder0_position[17]), .I1(n15_adj_5716), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5859));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5858));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5857));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
           .D(n17_adj_5897));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15762_3_lut_4_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29838));   // verilog/coms.v(130[12] 305[6])
    defparam i15762_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15761_3_lut_4_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29837));   // verilog/coms.v(130[12] 305[6])
    defparam i15761_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15760_3_lut_4_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29836));   // verilog/coms.v(130[12] 305[6])
    defparam i15760_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_2098 (.I0(n2126), .I1(n2125), .I2(GND_net), .I3(GND_net), 
            .O(n61576));
    defparam i1_2_lut_adj_2098.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25), .CO(n49744));
    SB_LUT4 mux_4310_i19_3_lut (.I0(encoder0_position[18]), .I1(n14_adj_5717), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i20_3_lut (.I0(encoder0_position[19]), .I1(n13_adj_5718), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i913_3_lut (.I0(n524), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15759_3_lut_4_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29835));   // verilog/coms.v(130[12] 305[6])
    defparam i15759_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i22_3_lut (.I0(encoder0_position[21]), .I1(n11_adj_5719), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i777_3_lut (.I0(n522), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233_adj_5811));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i844_3_lut (.I0(n1233_adj_5811), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5856));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15758_3_lut_4_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29834));   // verilog/coms.v(130[12] 305[6])
    defparam i15758_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15757_3_lut_4_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29833));   // verilog/coms.v(130[12] 305[6])
    defparam i15757_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15756_3_lut_4_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29832));   // verilog/coms.v(130[12] 305[6])
    defparam i15756_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16175_4_lut_4_lut (.I0(n27950), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n30251));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16175_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5855));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_2099 (.I0(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I1(Ki[1]), .I2(GND_net), .I3(GND_net), .O(n110));
    defparam i1_2_lut_adj_2099.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_2100 (.I0(state_adj_5979[2]), .I1(state_adj_5979[1]), 
            .I2(state_adj_5979[0]), .I3(n42792), .O(n56368));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_2100.LUT_INIT = 16'ha8e8;
    SB_LUT4 i15552_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[1]), .I2(n6), 
            .I3(n25583), .O(n29628));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15552_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15559_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[2]), .I2(n6), 
            .I3(n25590), .O(n29635));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15559_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15560_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[3]), .I2(n6), 
            .I3(n25578), .O(n29636));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15560_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15755_3_lut_4_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29831));   // verilog/coms.v(130[12] 305[6])
    defparam i15755_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[15] [7]), .I1(n57685), .I2(n57990), 
            .I3(\data_in_frame[16] [1]), .O(n32_adj_5849));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[16] [4]), .I1(Kp_23__N_1389), 
            .I2(n57862), .I3(n57625), .O(n31_adj_5850));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[13] [6]), 
            .I2(n53215), .I3(n52054), .O(n35_adj_5848));
    defparam i15_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut (.I0(n57737), .I1(n57499), .I2(n57657), .I3(\data_in_frame[16] [6]), 
            .O(n34));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_3_lut (.I0(n35_adj_5848), .I1(n31_adj_5850), .I2(n32_adj_5849), 
            .I3(GND_net), .O(n38_adj_5847));
    defparam i18_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_2101 (.I0(n26517), .I1(n58117), .I2(\data_in_frame[16] [0]), 
            .I3(n57956), .O(n33));
    defparam i13_4_lut_adj_2101.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15561_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[4]), .I2(n6_adj_5749), 
            .I3(n25615), .O(n29637));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15561_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15569_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[5]), .I2(n6_adj_5749), 
            .I3(n25583), .O(n29645));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15569_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15754_3_lut_4_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29830));   // verilog/coms.v(130[12] 305[6])
    defparam i15754_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15576_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[6]), .I2(n6_adj_5749), 
            .I3(n25590), .O(n29652));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15576_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15753_3_lut_4_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29829));   // verilog/coms.v(130[12] 305[6])
    defparam i15753_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15577_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[7]), .I2(n6_adj_5749), 
            .I3(n25578), .O(n29653));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15577_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15578_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[8]), .I2(n5_adj_5724), 
            .I3(n25587), .O(n29654));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15578_4_lut.LUT_INIT = 16'hccca;
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n55740));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i15751_3_lut_4_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29827));   // verilog/coms.v(130[12] 305[6])
    defparam i15751_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15579_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[9]), .I2(n6_adj_5748), 
            .I3(n25583), .O(n29655));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15579_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15750_3_lut_4_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29826));   // verilog/coms.v(130[12] 305[6])
    defparam i15750_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4_4_lut_adj_2102 (.I0(n53024), .I1(\data_in_frame[12] [4]), 
            .I2(n57819), .I3(n6_adj_5704), .O(n59684));
    defparam i4_4_lut_adj_2102.LUT_INIT = 16'h6996;
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n49520), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_2103 (.I0(n52186), .I1(n58132), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5903));
    defparam i1_2_lut_adj_2103.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_2104 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [0]), 
            .I2(n57879), .I3(n6_adj_5903), .O(n53127));
    defparam i4_4_lut_adj_2104.LUT_INIT = 16'h6996;
    SB_LUT4 i15580_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[10]), .I2(n5_adj_5798), 
            .I3(n25587), .O(n29656));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15580_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15586_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n22792), .I3(GND_net), .O(n29662));   // verilog/coms.v(130[12] 305[6])
    defparam i15586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(n62220), .I2(control_mode[7]), 
            .I3(control_mode[5]), .O(n25465));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15749_3_lut_4_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29825));   // verilog/coms.v(130[12] 305[6])
    defparam i15749_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15593_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(control_update), .I3(GND_net), .O(n29669));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15748_3_lut_4_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29824));   // verilog/coms.v(130[12] 305[6])
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15747_3_lut_4_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29823));   // verilog/coms.v(130[12] 305[6])
    defparam i15747_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15746_3_lut_4_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29822));   // verilog/coms.v(130[12] 305[6])
    defparam i15746_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15595_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[11]), .I2(n6_adj_5748), 
            .I3(n25578), .O(n29671));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15595_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15596_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[12]), .I2(n42880), 
            .I3(n25615), .O(n29672));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15596_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15745_3_lut_4_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29821));   // verilog/coms.v(130[12] 305[6])
    defparam i15745_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15744_3_lut_4_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29820));   // verilog/coms.v(130[12] 305[6])
    defparam i15744_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY add_151_12 (.CI(n49520), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n49521));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n49541), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2105 (.I0(state_adj_5979[2]), .I1(data_ready), 
            .I2(n3_adj_5800), .I3(n25612), .O(n56774));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_2105.LUT_INIT = 16'hcca8;
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n49540), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15599_3_lut (.I0(current[0]), .I1(data_adj_5985[0]), .I2(n27736), 
            .I3(GND_net), .O(n29675));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15600_4_lut (.I0(rw), .I1(state_adj_5979[1]), .I2(state_adj_5979[2]), 
            .I3(n5774), .O(n29676));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15600_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i15601_3_lut (.I0(CS_c), .I1(state_adj_5987[0]), .I2(state_adj_5987[1]), 
            .I3(GND_net), .O(n29677));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15601_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i29710_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n43685));
    defparam i29710_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i53710_4_lut (.I0(n15_adj_5750), .I1(clk_out), .I2(state_adj_5987[0]), 
            .I3(state_adj_5987[1]), .O(n9_adj_5916));   // verilog/tli4970.v(35[10] 68[6])
    defparam i53710_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 encoder0_position_30__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15743_3_lut_4_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29819));   // verilog/coms.v(130[12] 305[6])
    defparam i15743_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27728), 
            .D(n1239), .R(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i15607_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(n57392), .I3(state_7__N_4108[0]), 
            .O(n29683));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15607_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_4_lut_adj_2106 (.I0(n2122), .I1(n2128), .I2(n61576), .I3(n2127), 
            .O(n61580));
    defparam i1_4_lut_adj_2106.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_766_11_lut (.I0(n69297), .I1(n1125), 
            .I2(VCC_net), .I3(n49880), .O(n1224_adj_5802)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n49879), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_10 (.CI(n49879), .I0(n1126), 
            .I1(VCC_net), .CO(n49880));
    SB_LUT4 encoder0_position_30__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n49878), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_18_lut (.I0(GND_net), .I1(n1818), 
            .I2(VCC_net), .I3(n50107), .O(n1885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n27676), .D(GHC_N_391), 
            .R(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n27676), .D(GHB_N_377), 
            .R(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n27676), .D(GHA_N_355), 
            .R(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n50106), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5924), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n27676), .D(GLA_N_372), 
            .R(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[25]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[24]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n27676), .D(GLB_N_386), 
            .R(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n27676), .D(GLC_N_400), 
            .R(n28908));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_30__I_0_add_1235_17 (.CI(n50106), .I0(n1819), 
            .I1(VCC_net), .CO(n50107));
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_30__I_0_add_766_9 (.CI(n49878), .I0(n1127), 
            .I1(VCC_net), .CO(n49879));
    SB_LUT4 encoder0_position_30__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n50105), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_2107 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57819));
    defparam i1_2_lut_adj_2107.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1235_16 (.CI(n50105), .I0(n1820), 
            .I1(VCC_net), .CO(n50106));
    SB_LUT4 encoder0_position_30__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n49877), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_8 (.CI(n49877), .I0(n1128), 
            .I1(VCC_net), .CO(n49878));
    SB_LUT4 encoder0_position_30__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n50104), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_15 (.CI(n50104), .I0(n1821), 
            .I1(VCC_net), .CO(n50105));
    SB_LUT4 encoder0_position_30__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822_adj_5818), 
            .I2(VCC_net), .I3(n50103), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n49876), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_14 (.CI(n50103), .I0(n1822_adj_5818), 
            .I1(VCC_net), .CO(n50104));
    SB_CARRY add_151_5 (.CI(n49513), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n49514));
    SB_LUT4 encoder0_position_30__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n50102), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_13 (.CI(n50102), .I0(n1823), 
            .I1(VCC_net), .CO(n50103));
    SB_LUT4 encoder0_position_30__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824_adj_5819), 
            .I2(VCC_net), .I3(n50101), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_7 (.CI(n49876), .I0(n1129), 
            .I1(GND_net), .CO(n49877));
    SB_CARRY encoder0_position_30__I_0_add_1235_12 (.CI(n50101), .I0(n1824_adj_5819), 
            .I1(VCC_net), .CO(n50102));
    SB_LUT4 add_2510_25_lut (.I0(n69378), .I1(n2_adj_5855), .I2(n1059), 
            .I3(n50523), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n50100), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2510_24_lut (.I0(n69297), .I1(n2_adj_5855), .I2(n1158), 
            .I3(n50522), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_24 (.CI(n50522), .I0(n2_adj_5855), .I1(n1158), .CO(n50523));
    SB_LUT4 add_2510_23_lut (.I0(n69365), .I1(n2_adj_5855), .I2(n1257), 
            .I3(n50521), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1235_11 (.CI(n50100), .I0(n1825), 
            .I1(VCC_net), .CO(n50101));
    SB_CARRY add_2510_23 (.CI(n50521), .I0(n2_adj_5855), .I1(n1257), .CO(n50522));
    SB_LUT4 add_2510_22_lut (.I0(n69303), .I1(n2_adj_5855), .I2(n1356), 
            .I3(n50520), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n50099), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n49875), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_22 (.CI(n50520), .I0(n2_adj_5855), .I1(n1356), .CO(n50521));
    SB_LUT4 add_2510_21_lut (.I0(n69350), .I1(n2_adj_5855), .I2(n1455), 
            .I3(n50519), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_21 (.CI(n50519), .I0(n2_adj_5855), .I1(n1455), .CO(n50520));
    SB_CARRY encoder0_position_30__I_0_add_1235_10 (.CI(n50099), .I0(n1826), 
            .I1(VCC_net), .CO(n50100));
    SB_LUT4 add_2510_20_lut (.I0(n69333), .I1(n2_adj_5855), .I2(n1554), 
            .I3(n50518), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_20 (.CI(n50518), .I0(n2_adj_5855), .I1(n1554), .CO(n50519));
    SB_LUT4 encoder0_position_30__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n50098), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_9 (.CI(n50098), .I0(n1827), 
            .I1(VCC_net), .CO(n50099));
    SB_LUT4 add_2510_19_lut (.I0(n69225), .I1(n2_adj_5855), .I2(n1653), 
            .I3(n50517), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n49519), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_19 (.CI(n50517), .I0(n2_adj_5855), .I1(n1653), .CO(n50518));
    SB_LUT4 add_2510_18_lut (.I0(n69206), .I1(n2_adj_5855), .I2(n1752), 
            .I3(n50516), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n50097), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_18 (.CI(n50516), .I0(n2_adj_5855), .I1(n1752), .CO(n50517));
    SB_LUT4 add_2510_17_lut (.I0(n69184), .I1(n2_adj_5855), .I2(n1851), 
            .I3(n50515), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1235_8 (.CI(n50097), .I0(n1828), 
            .I1(VCC_net), .CO(n50098));
    SB_CARRY add_2510_17 (.CI(n50515), .I0(n2_adj_5855), .I1(n1851), .CO(n50516));
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n49512), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2510_16_lut (.I0(n69088), .I1(n2_adj_5855), .I2(n1950), 
            .I3(n50514), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_16 (.CI(n50514), .I0(n2_adj_5855), .I1(n1950), .CO(n50515));
    SB_LUT4 encoder0_position_30__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n50096), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2510_15_lut (.I0(n69092), .I1(n2_adj_5855), .I2(n2049), 
            .I3(n50513), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_15 (.CI(n50513), .I0(n2_adj_5855), .I1(n2049), .CO(n50514));
    SB_LUT4 add_2510_14_lut (.I0(n69135), .I1(n2_adj_5855), .I2(n2148), 
            .I3(n50512), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_14 (.CI(n50512), .I0(n2_adj_5855), .I1(n2148), .CO(n50513));
    SB_LUT4 add_2510_13_lut (.I0(n69160), .I1(n2_adj_5855), .I2(n2247), 
            .I3(n50511), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_13 (.CI(n50511), .I0(n2_adj_5855), .I1(n2247), .CO(n50512));
    SB_CARRY encoder0_position_30__I_0_add_1235_7 (.CI(n50096), .I0(n1829), 
            .I1(GND_net), .CO(n50097));
    SB_LUT4 i15615_4_lut (.I0(CS_MISO_c), .I1(data_adj_5985[15]), .I2(n42880), 
            .I3(n25578), .O(n29691));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15615_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_30__I_0_add_766_6 (.CI(n49875), .I0(n1130), 
            .I1(GND_net), .CO(n49876));
    SB_LUT4 add_2510_12_lut (.I0(n68974), .I1(n2_adj_5855), .I2(n2346), 
            .I3(n50510), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_12 (.CI(n50510), .I0(n2_adj_5855), .I1(n2346), .CO(n50511));
    SB_LUT4 encoder0_position_30__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n49874), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n50095), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_6 (.CI(n50095), .I0(n1830), 
            .I1(GND_net), .CO(n50096));
    SB_LUT4 add_2510_11_lut (.I0(n69006), .I1(n2_adj_5855), .I2(n2445), 
            .I3(n50509), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_151_32 (.CI(n49540), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n49541));
    SB_CARRY add_151_11 (.CI(n49519), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n49520));
    SB_CARRY add_2510_11 (.CI(n50509), .I0(n2_adj_5855), .I1(n2445), .CO(n50510));
    SB_LUT4 add_2510_10_lut (.I0(n69034), .I1(n2_adj_5855), .I2(n2544), 
            .I3(n50508), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_10 (.CI(n50508), .I0(n2_adj_5855), .I1(n2544), .CO(n50509));
    SB_CARRY encoder0_position_30__I_0_add_766_5 (.CI(n49874), .I0(n1131), 
            .I1(VCC_net), .CO(n49875));
    SB_LUT4 add_2510_9_lut (.I0(n69063), .I1(n2_adj_5855), .I2(n2643), 
            .I3(n50507), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n49539), .O(n1210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n49539), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n49540));
    SB_LUT4 encoder0_position_30__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n49873), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n50094), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_9 (.CI(n50507), .I0(n2_adj_5855), .I1(n2643), .CO(n50508));
    SB_LUT4 add_2510_8_lut (.I0(n68948), .I1(n2_adj_5855), .I2(n2742), 
            .I3(n50506), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_8 (.CI(n50506), .I0(n2_adj_5855), .I1(n2742), .CO(n50507));
    SB_LUT4 add_2510_7_lut (.I0(n68915), .I1(n2_adj_5855), .I2(n2841), 
            .I3(n50505), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1235_5 (.CI(n50094), .I0(n1831), 
            .I1(VCC_net), .CO(n50095));
    SB_CARRY encoder0_position_30__I_0_add_766_4 (.CI(n49873), .I0(n1132), 
            .I1(GND_net), .CO(n49874));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n49538), .O(n1211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n49872), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_3 (.CI(n49872), .I0(n1133), 
            .I1(VCC_net), .CO(n49873));
    SB_LUT4 encoder0_position_30__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n50093), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_7 (.CI(n50505), .I0(n2_adj_5855), .I1(n2841), .CO(n50506));
    SB_LUT4 add_2510_6_lut (.I0(n68881), .I1(n2_adj_5855), .I2(n2940), 
            .I3(n50504), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_6 (.CI(n50504), .I0(n2_adj_5855), .I1(n2940), .CO(n50505));
    SB_LUT4 add_2510_5_lut (.I0(n68809), .I1(n2_adj_5855), .I2(n3039), 
            .I3(n50503), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_1235_4 (.CI(n50093), .I0(n1832), 
            .I1(GND_net), .CO(n50094));
    SB_LUT4 encoder0_position_30__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n50092), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_3 (.CI(n50092), .I0(n1833), 
            .I1(VCC_net), .CO(n50093));
    SB_LUT4 encoder0_position_30__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_5 (.CI(n50503), .I0(n2_adj_5855), .I1(n3039), .CO(n50504));
    SB_CARRY encoder0_position_30__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n50092));
    SB_LUT4 encoder0_position_30__I_0_add_766_2_lut (.I0(GND_net), .I1(n522), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2510_4_lut (.I0(n68813), .I1(n2_adj_5855), .I2(n3138), 
            .I3(n50502), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_766_2 (.CI(VCC_net), .I0(n522), 
            .I1(GND_net), .CO(n49872));
    SB_CARRY add_2510_4 (.CI(n50502), .I0(n2_adj_5855), .I1(n3138), .CO(n50503));
    SB_LUT4 add_2510_3_lut (.I0(n68744), .I1(n2_adj_5855), .I2(n3237), 
            .I3(n50501), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_3 (.CI(n50501), .I0(n2_adj_5855), .I1(n3237), .CO(n50502));
    SB_LUT4 add_2510_2_lut (.I0(n68740), .I1(n2_adj_5855), .I2(n43717), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_2 (.CI(VCC_net), .I0(n2_adj_5855), .I1(n43717), 
            .CO(n50501));
    SB_LUT4 encoder0_position_30__I_0_add_2173_33_lut (.I0(n68744), .I1(n3204), 
            .I2(VCC_net), .I3(n50500), .O(n62647)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n50499), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_32 (.CI(n50499), .I0(n3205), 
            .I1(VCC_net), .CO(n50500));
    SB_LUT4 encoder0_position_30__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n50498), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_31 (.CI(n50498), .I0(n3206), 
            .I1(VCC_net), .CO(n50499));
    SB_LUT4 encoder0_position_30__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n50497), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_30 (.CI(n50497), .I0(n3207), 
            .I1(VCC_net), .CO(n50498));
    SB_LUT4 encoder0_position_30__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n50496), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_29 (.CI(n50496), .I0(n3208), 
            .I1(VCC_net), .CO(n50497));
    SB_LUT4 encoder0_position_30__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n50495), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_28 (.CI(n50495), .I0(n3209), 
            .I1(VCC_net), .CO(n50496));
    SB_LUT4 encoder0_position_30__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n50494), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_27 (.CI(n50494), .I0(n3210), 
            .I1(VCC_net), .CO(n50495));
    SB_LUT4 encoder0_position_30__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n50493), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_26 (.CI(n50493), .I0(n3211), 
            .I1(VCC_net), .CO(n50494));
    SB_LUT4 encoder0_position_30__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n50492), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_25 (.CI(n50492), .I0(n3212), 
            .I1(VCC_net), .CO(n50493));
    SB_LUT4 encoder0_position_30__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n50491), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_24 (.CI(n50491), .I0(n3213), 
            .I1(VCC_net), .CO(n50492));
    SB_LUT4 encoder0_position_30__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n50490), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_23 (.CI(n50490), .I0(n3214), 
            .I1(VCC_net), .CO(n50491));
    SB_LUT4 encoder0_position_30__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n50489), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_22 (.CI(n50489), .I0(n3215), 
            .I1(VCC_net), .CO(n50490));
    SB_LUT4 encoder0_position_30__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n50488), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_21 (.CI(n50488), .I0(n3216), 
            .I1(VCC_net), .CO(n50489));
    SB_LUT4 encoder0_position_30__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n50487), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_20 (.CI(n50487), .I0(n3217), 
            .I1(VCC_net), .CO(n50488));
    SB_LUT4 encoder0_position_30__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n50486), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_19 (.CI(n50486), .I0(n3218), 
            .I1(VCC_net), .CO(n50487));
    SB_LUT4 encoder0_position_30__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n50485), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_18 (.CI(n50485), .I0(n3219), 
            .I1(VCC_net), .CO(n50486));
    SB_LUT4 encoder0_position_30__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n50484), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_17 (.CI(n50484), .I0(n3220), 
            .I1(VCC_net), .CO(n50485));
    SB_LUT4 encoder0_position_30__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n50483), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_16 (.CI(n50483), .I0(n3221), 
            .I1(VCC_net), .CO(n50484));
    SB_LUT4 encoder0_position_30__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n50482), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_15 (.CI(n50482), .I0(n3222), 
            .I1(VCC_net), .CO(n50483));
    SB_LUT4 encoder0_position_30__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n50481), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_30 (.CI(n49538), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n49539));
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n49537), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_14 (.CI(n50481), .I0(n3223), 
            .I1(VCC_net), .CO(n50482));
    SB_LUT4 encoder0_position_30__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n50480), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_13 (.CI(n50480), .I0(n3224), 
            .I1(VCC_net), .CO(n50481));
    SB_LUT4 encoder0_position_30__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n50479), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_12 (.CI(n50479), .I0(n3225), 
            .I1(VCC_net), .CO(n50480));
    SB_LUT4 encoder0_position_30__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n50478), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_11 (.CI(n50478), .I0(n3226), 
            .I1(VCC_net), .CO(n50479));
    SB_LUT4 encoder0_position_30__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n50477), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_10 (.CI(n50477), .I0(n3227), 
            .I1(VCC_net), .CO(n50478));
    SB_LUT4 encoder0_position_30__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n50476), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_9 (.CI(n50476), .I0(n3228), 
            .I1(VCC_net), .CO(n50477));
    SB_LUT4 encoder0_position_30__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n50475), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_8 (.CI(n50475), .I0(n3229), 
            .I1(GND_net), .CO(n50476));
    SB_LUT4 encoder0_position_30__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n50474), .O(n65588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_7 (.CI(n50474), .I0(n3230), 
            .I1(GND_net), .CO(n50475));
    SB_LUT4 encoder0_position_30__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n50473), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_6 (.CI(n50473), .I0(n3231), 
            .I1(VCC_net), .CO(n50474));
    SB_LUT4 i15623_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n22792), .I3(GND_net), .O(n29699));   // verilog/coms.v(130[12] 305[6])
    defparam i15623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_2173_5_lut (.I0(n6_adj_5852), .I1(n3232), 
            .I2(GND_net), .I3(n50472), .O(n65579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_30__I_0_add_2173_5 (.CI(n50472), .I0(n3232), 
            .I1(GND_net), .CO(n50473));
    SB_LUT4 encoder0_position_30__I_0_add_2173_4_lut (.I0(n3301), .I1(n3233), 
            .I2(VCC_net), .I3(n50471), .O(n6_adj_5852)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_4 (.CI(n50471), .I0(n3233), 
            .I1(VCC_net), .CO(n50472));
    SB_LUT4 encoder0_position_30__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n50470), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_3 (.CI(n50470), .I0(n957), 
            .I1(GND_net), .CO(n50471));
    SB_CARRY encoder0_position_30__I_0_add_2173_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n50470));
    SB_LUT4 encoder0_position_30__I_0_add_2106_31_lut (.I0(n68813), .I1(n3105), 
            .I2(VCC_net), .I3(n50469), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n50468), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_30 (.CI(n50468), .I0(n3106), 
            .I1(VCC_net), .CO(n50469));
    SB_LUT4 i15624_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n22792), .I3(GND_net), .O(n29700));   // verilog/coms.v(130[12] 305[6])
    defparam i15624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n50467), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_29 (.CI(n50467), .I0(n3107), 
            .I1(VCC_net), .CO(n50468));
    SB_LUT4 encoder0_position_30__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n50466), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_28 (.CI(n50466), .I0(n3108), 
            .I1(VCC_net), .CO(n50467));
    SB_LUT4 encoder0_position_30__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n50465), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_27 (.CI(n50465), .I0(n3109), 
            .I1(VCC_net), .CO(n50466));
    SB_LUT4 encoder0_position_30__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n50464), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_26 (.CI(n50464), .I0(n3110), 
            .I1(VCC_net), .CO(n50465));
    SB_LUT4 encoder0_position_30__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n50463), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_25 (.CI(n50463), .I0(n3111), 
            .I1(VCC_net), .CO(n50464));
    SB_LUT4 encoder0_position_30__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n50462), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_24 (.CI(n50462), .I0(n3112), 
            .I1(VCC_net), .CO(n50463));
    SB_LUT4 encoder0_position_30__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n50461), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_23 (.CI(n50461), .I0(n3113), 
            .I1(VCC_net), .CO(n50462));
    SB_LUT4 encoder0_position_30__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n50460), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_22 (.CI(n50460), .I0(n3114), 
            .I1(VCC_net), .CO(n50461));
    SB_LUT4 encoder0_position_30__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n50459), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_21 (.CI(n50459), .I0(n3115), 
            .I1(VCC_net), .CO(n50460));
    SB_LUT4 encoder0_position_30__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n50458), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_20 (.CI(n50458), .I0(n3116), 
            .I1(VCC_net), .CO(n50459));
    SB_LUT4 encoder0_position_30__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n50457), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_29 (.CI(n49537), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n49538));
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n49536), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_19 (.CI(n50457), .I0(n3117), 
            .I1(VCC_net), .CO(n50458));
    SB_LUT4 add_1097_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n49650), .O(n4905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n50456), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_18 (.CI(n50456), .I0(n3118), 
            .I1(VCC_net), .CO(n50457));
    SB_CARRY add_151_28 (.CI(n49536), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n49537));
    SB_LUT4 encoder0_position_30__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n50455), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_24_lut (.I0(GND_net), .I1(GND_net), .I2(n12185), 
            .I3(n49649), .O(n4906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_17_lut (.I0(n69206), .I1(n1719), 
            .I2(VCC_net), .I3(n50072), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1097_24 (.CI(n49649), .I0(GND_net), .I1(n12185), .CO(n49650));
    SB_CARRY encoder0_position_30__I_0_add_2106_17 (.CI(n50455), .I0(n3119), 
            .I1(VCC_net), .CO(n50456));
    SB_LUT4 encoder0_position_30__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n50454), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n49535), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n49853), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n50071), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_16 (.CI(n50071), .I0(n1720), 
            .I1(VCC_net), .CO(n50072));
    SB_LUT4 encoder0_position_30__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n49852), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_16 (.CI(n50454), .I0(n3120), 
            .I1(VCC_net), .CO(n50455));
    SB_LUT4 encoder0_position_30__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n50453), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n50070), .O(n1788_adj_5813)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_15 (.CI(n50070), .I0(n1721), 
            .I1(VCC_net), .CO(n50071));
    SB_CARRY encoder0_position_30__I_0_add_699_9 (.CI(n49852), .I0(n1027), 
            .I1(VCC_net), .CO(n49853));
    SB_LUT4 add_1097_23_lut (.I0(GND_net), .I1(GND_net), .I2(n12187), 
            .I3(n49648), .O(n4907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n49851), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n50069), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_14 (.CI(n50069), .I0(n1722), 
            .I1(VCC_net), .CO(n50070));
    SB_CARRY encoder0_position_30__I_0_add_699_8 (.CI(n49851), .I0(n1028), 
            .I1(VCC_net), .CO(n49852));
    SB_CARRY encoder0_position_30__I_0_add_2106_15 (.CI(n50453), .I0(n3121), 
            .I1(VCC_net), .CO(n50454));
    SB_LUT4 encoder0_position_30__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n50068), .O(n1790_adj_5814)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n49850), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n50452), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_14 (.CI(n50452), .I0(n3122), 
            .I1(VCC_net), .CO(n50453));
    SB_CARRY encoder0_position_30__I_0_add_1168_13 (.CI(n50068), .I0(n1723), 
            .I1(VCC_net), .CO(n50069));
    SB_CARRY encoder0_position_30__I_0_add_699_7 (.CI(n49850), .I0(n1029), 
            .I1(GND_net), .CO(n49851));
    SB_CARRY add_1097_23 (.CI(n49648), .I0(GND_net), .I1(n12187), .CO(n49649));
    SB_LUT4 encoder0_position_30__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n50067), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n50451), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n49849), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_12 (.CI(n50067), .I0(n1724), 
            .I1(VCC_net), .CO(n50068));
    SB_LUT4 encoder0_position_30__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n50066), .O(n1792_adj_5815)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_22_lut (.I0(GND_net), .I1(GND_net), .I2(n12189), 
            .I3(n49647), .O(n4908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_22 (.CI(n49647), .I0(GND_net), .I1(n12189), .CO(n49648));
    SB_LUT4 add_1097_21_lut (.I0(GND_net), .I1(GND_net), .I2(n12191), 
            .I3(n49646), .O(n4909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_6 (.CI(n49849), .I0(n1030), 
            .I1(GND_net), .CO(n49850));
    SB_LUT4 encoder0_position_30__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n49848), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_11 (.CI(n50066), .I0(n1725), 
            .I1(VCC_net), .CO(n50067));
    SB_CARRY encoder0_position_30__I_0_add_2106_13 (.CI(n50451), .I0(n3123), 
            .I1(VCC_net), .CO(n50452));
    SB_LUT4 encoder0_position_30__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n50450), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_27 (.CI(n49535), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n49536));
    SB_CARRY add_1097_21 (.CI(n49646), .I0(GND_net), .I1(n12191), .CO(n49647));
    SB_LUT4 encoder0_position_30__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n50065), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_5 (.CI(n49848), .I0(n1031), 
            .I1(VCC_net), .CO(n49849));
    SB_CARRY encoder0_position_30__I_0_add_1168_10 (.CI(n50065), .I0(n1726), 
            .I1(VCC_net), .CO(n50066));
    SB_LUT4 encoder0_position_30__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n49847), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_4 (.CI(n49847), .I0(n1032), 
            .I1(GND_net), .CO(n49848));
    SB_LUT4 encoder0_position_30__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n49846), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_12 (.CI(n50450), .I0(n3124), 
            .I1(VCC_net), .CO(n50451));
    SB_LUT4 encoder0_position_30__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n50449), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n49534), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_20_lut (.I0(GND_net), .I1(GND_net), .I2(n12193), 
            .I3(n49645), .O(n4910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_11 (.CI(n50449), .I0(n3125), 
            .I1(VCC_net), .CO(n50450));
    SB_CARRY encoder0_position_30__I_0_add_699_3 (.CI(n49846), .I0(n1033), 
            .I1(VCC_net), .CO(n49847));
    SB_LUT4 encoder0_position_30__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n50448), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n50064), .O(n1794_adj_5816)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_10 (.CI(n50448), .I0(n3126), 
            .I1(VCC_net), .CO(n50449));
    SB_LUT4 encoder0_position_30__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n50447), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_26 (.CI(n49534), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n49535));
    SB_CARRY encoder0_position_30__I_0_add_699_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n49846));
    SB_CARRY encoder0_position_30__I_0_add_1168_9 (.CI(n50064), .I0(n1727), 
            .I1(VCC_net), .CO(n50065));
    SB_LUT4 encoder0_position_30__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n50063), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_9 (.CI(n50447), .I0(n3127), 
            .I1(VCC_net), .CO(n50448));
    SB_LUT4 encoder0_position_30__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n50446), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_8 (.CI(n50446), .I0(n3128), 
            .I1(VCC_net), .CO(n50447));
    SB_CARRY encoder0_position_30__I_0_add_1168_8 (.CI(n50063), .I0(n1728), 
            .I1(VCC_net), .CO(n50064));
    SB_LUT4 encoder0_position_30__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n50445), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_7 (.CI(n50445), .I0(n3129), 
            .I1(GND_net), .CO(n50446));
    SB_LUT4 encoder0_position_30__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n50444), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_6 (.CI(n50444), .I0(n3130), 
            .I1(GND_net), .CO(n50445));
    SB_LUT4 encoder0_position_30__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n50062), .O(n1796_adj_5817)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n50443), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_7 (.CI(n50062), .I0(n1729), 
            .I1(GND_net), .CO(n50063));
    SB_CARRY add_1097_20 (.CI(n49645), .I0(GND_net), .I1(n12193), .CO(n49646));
    SB_CARRY encoder0_position_30__I_0_add_2106_5 (.CI(n50443), .I0(n3131), 
            .I1(VCC_net), .CO(n50444));
    SB_LUT4 mux_4310_i25_3_lut (.I0(encoder0_position[24]), .I1(n8_adj_5721), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1097_19_lut (.I0(GND_net), .I1(GND_net), .I2(n12195), 
            .I3(n49644), .O(n4911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n50442), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n50061), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_6 (.CI(n50061), .I0(n1730), 
            .I1(GND_net), .CO(n50062));
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n49518), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_4 (.CI(n50442), .I0(n3132), 
            .I1(GND_net), .CO(n50443));
    SB_LUT4 encoder0_position_30__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n50060), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15631_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n29707));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15631_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n50441), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_5 (.CI(n50060), .I0(n1731), 
            .I1(VCC_net), .CO(n50061));
    SB_LUT4 encoder0_position_30__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n50059), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_4 (.CI(n50059), .I0(n1732), 
            .I1(GND_net), .CO(n50060));
    SB_CARRY encoder0_position_30__I_0_add_2106_3 (.CI(n50441), .I0(n3133), 
            .I1(VCC_net), .CO(n50442));
    SB_LUT4 encoder0_position_30__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n50058), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_3 (.CI(n50058), .I0(n1733), 
            .I1(VCC_net), .CO(n50059));
    SB_LUT4 encoder0_position_30__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_19 (.CI(n49644), .I0(GND_net), .I1(n12195), .CO(n49645));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n49533), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n50058));
    SB_CARRY encoder0_position_30__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n50441));
    SB_LUT4 add_1097_18_lut (.I0(GND_net), .I1(GND_net), .I2(n12197), 
            .I3(n49643), .O(n4912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_30_lut (.I0(n68809), .I1(n3006), 
            .I2(VCC_net), .I3(n50440), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n50439), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_29 (.CI(n50439), .I0(n3007), 
            .I1(VCC_net), .CO(n50440));
    SB_CARRY add_1097_18 (.CI(n49643), .I0(GND_net), .I1(n12197), .CO(n49644));
    SB_CARRY add_151_4 (.CI(n49512), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n49513));
    SB_LUT4 encoder0_position_30__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n50438), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_28 (.CI(n50438), .I0(n3008), 
            .I1(VCC_net), .CO(n50439));
    SB_LUT4 encoder0_position_30__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n50437), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_27 (.CI(n50437), .I0(n3009), 
            .I1(VCC_net), .CO(n50438));
    SB_LUT4 add_1097_17_lut (.I0(GND_net), .I1(GND_net), .I2(n12199), 
            .I3(n49642), .O(n4913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n50436), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_26 (.CI(n50436), .I0(n3010), 
            .I1(VCC_net), .CO(n50437));
    SB_CARRY add_151_25 (.CI(n49533), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n49534));
    SB_LUT4 encoder0_position_30__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n50435), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_17 (.CI(n49642), .I0(GND_net), .I1(n12199), .CO(n49643));
    SB_CARRY encoder0_position_30__I_0_add_2039_25 (.CI(n50435), .I0(n3011), 
            .I1(VCC_net), .CO(n50436));
    SB_LUT4 encoder0_position_30__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n50434), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_24 (.CI(n50434), .I0(n3012), 
            .I1(VCC_net), .CO(n50435));
    SB_CARRY add_151_10 (.CI(n49518), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n49519));
    SB_LUT4 encoder0_position_30__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n50433), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_16_lut (.I0(GND_net), .I1(GND_net), .I2(n12201), 
            .I3(n49641), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7479_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n20965));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i7479_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n49532), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_23 (.CI(n50433), .I0(n3013), 
            .I1(VCC_net), .CO(n50434));
    SB_LUT4 encoder0_position_30__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n50432), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_22 (.CI(n50432), .I0(n3014), 
            .I1(VCC_net), .CO(n50433));
    SB_LUT4 encoder0_position_30__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n50431), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_21 (.CI(n50431), .I0(n3015), 
            .I1(VCC_net), .CO(n50432));
    SB_LUT4 encoder0_position_30__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n50430), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_20 (.CI(n50430), .I0(n3016), 
            .I1(VCC_net), .CO(n50431));
    SB_LUT4 encoder0_position_30__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n50429), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_19 (.CI(n50429), .I0(n3017), 
            .I1(VCC_net), .CO(n50430));
    SB_LUT4 encoder0_position_30__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n50428), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_18 (.CI(n50428), .I0(n3018), 
            .I1(VCC_net), .CO(n50429));
    SB_LUT4 encoder0_position_30__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n50427), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_17 (.CI(n50427), .I0(n3019), 
            .I1(VCC_net), .CO(n50428));
    SB_LUT4 encoder0_position_30__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n50426), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_16 (.CI(n50426), .I0(n3020), 
            .I1(VCC_net), .CO(n50427));
    SB_LUT4 encoder0_position_30__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n50425), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n49532), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n49533));
    SB_CARRY encoder0_position_30__I_0_add_2039_15 (.CI(n50425), .I0(n3021), 
            .I1(VCC_net), .CO(n50426));
    SB_LUT4 encoder0_position_30__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n50424), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_14 (.CI(n50424), .I0(n3022), 
            .I1(VCC_net), .CO(n50425));
    SB_LUT4 encoder0_position_30__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n50423), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_13 (.CI(n50423), .I0(n3023), 
            .I1(VCC_net), .CO(n50424));
    SB_LUT4 encoder0_position_30__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n50422), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n49531), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_12 (.CI(n50422), .I0(n3024), 
            .I1(VCC_net), .CO(n50423));
    SB_LUT4 encoder0_position_30__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n50421), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_11 (.CI(n50421), .I0(n3025), 
            .I1(VCC_net), .CO(n50422));
    SB_LUT4 encoder0_position_30__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n50420), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_10 (.CI(n50420), .I0(n3026), 
            .I1(VCC_net), .CO(n50421));
    SB_LUT4 encoder0_position_30__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n50419), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_9 (.CI(n50419), .I0(n3027), 
            .I1(VCC_net), .CO(n50420));
    SB_LUT4 encoder0_position_30__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n50418), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8783_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i8783_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY encoder0_position_30__I_0_add_2039_8 (.CI(n50418), .I0(n3028), 
            .I1(VCC_net), .CO(n50419));
    SB_LUT4 encoder0_position_30__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n50417), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_7 (.CI(n50417), .I0(n3029), 
            .I1(GND_net), .CO(n50418));
    SB_LUT4 encoder0_position_30__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n50416), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_6 (.CI(n50416), .I0(n3030), 
            .I1(GND_net), .CO(n50417));
    SB_LUT4 encoder0_position_30__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n50415), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_5 (.CI(n50415), .I0(n3031), 
            .I1(VCC_net), .CO(n50416));
    SB_LUT4 encoder0_position_30__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n50414), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_16 (.CI(n49641), .I0(GND_net), .I1(n12201), .CO(n49642));
    SB_CARRY encoder0_position_30__I_0_add_2039_4 (.CI(n50414), .I0(n3032), 
            .I1(GND_net), .CO(n50415));
    SB_LUT4 encoder0_position_30__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n50413), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_3 (.CI(n50413), .I0(n3033), 
            .I1(VCC_net), .CO(n50414));
    SB_LUT4 encoder0_position_30__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n50413));
    SB_LUT4 add_1097_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12203), 
            .I3(n49640), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_29_lut (.I0(n68881), .I1(n2907), 
            .I2(VCC_net), .I3(n50412), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n50411), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_28 (.CI(n50411), .I0(n2908), 
            .I1(VCC_net), .CO(n50412));
    SB_LUT4 encoder0_position_30__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n50410), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_27 (.CI(n50410), .I0(n2909), 
            .I1(VCC_net), .CO(n50411));
    SB_LUT4 encoder0_position_30__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n50409), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_26 (.CI(n50409), .I0(n2910), 
            .I1(VCC_net), .CO(n50410));
    SB_CARRY add_1097_15 (.CI(n49640), .I0(GND_net), .I1(n12203), .CO(n49641));
    SB_LUT4 encoder0_position_30__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n50408), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n49517), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_25 (.CI(n50408), .I0(n2911), 
            .I1(VCC_net), .CO(n50409));
    SB_LUT4 encoder0_position_30__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n50407), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_14_lut (.I0(GND_net), .I1(GND_net), .I2(n12205), 
            .I3(n49639), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_24 (.CI(n50407), .I0(n2912), 
            .I1(VCC_net), .CO(n50408));
    SB_CARRY add_1097_14 (.CI(n49639), .I0(GND_net), .I1(n12205), .CO(n49640));
    SB_LUT4 encoder0_position_30__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n50406), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_23 (.CI(n50406), .I0(n2913), 
            .I1(VCC_net), .CO(n50407));
    SB_LUT4 encoder0_position_30__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n50405), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_22 (.CI(n50405), .I0(n2914), 
            .I1(VCC_net), .CO(n50406));
    SB_LUT4 add_1097_13_lut (.I0(GND_net), .I1(GND_net), .I2(n12207), 
            .I3(n49638), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n49531), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n49532));
    SB_LUT4 encoder0_position_30__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n50404), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_21 (.CI(n50404), .I0(n2915), 
            .I1(VCC_net), .CO(n50405));
    SB_LUT4 encoder0_position_30__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n50403), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_20 (.CI(n50403), .I0(n2916), 
            .I1(VCC_net), .CO(n50404));
    SB_CARRY add_1097_13 (.CI(n49638), .I0(GND_net), .I1(n12207), .CO(n49639));
    SB_LUT4 encoder0_position_30__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n50402), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_19 (.CI(n50402), .I0(n2917), 
            .I1(VCC_net), .CO(n50403));
    SB_LUT4 encoder0_position_30__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n50401), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_18 (.CI(n50401), .I0(n2918), 
            .I1(VCC_net), .CO(n50402));
    SB_LUT4 encoder0_position_30__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n50400), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_17 (.CI(n50400), .I0(n2919), 
            .I1(VCC_net), .CO(n50401));
    SB_LUT4 encoder0_position_30__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n50399), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_16 (.CI(n50399), .I0(n2920), 
            .I1(VCC_net), .CO(n50400));
    SB_LUT4 encoder0_position_30__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n50398), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_15 (.CI(n50398), .I0(n2921), 
            .I1(VCC_net), .CO(n50399));
    SB_LUT4 encoder0_position_30__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n50397), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_14 (.CI(n50397), .I0(n2922), 
            .I1(VCC_net), .CO(n50398));
    SB_LUT4 encoder0_position_30__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n50396), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_12_lut (.I0(GND_net), .I1(GND_net), .I2(n12209), 
            .I3(n49637), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_13 (.CI(n50396), .I0(n2923), 
            .I1(VCC_net), .CO(n50397));
    SB_LUT4 encoder0_position_30__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n50395), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_12 (.CI(n50395), .I0(n2924), 
            .I1(VCC_net), .CO(n50396));
    SB_LUT4 encoder0_position_30__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n50394), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_12 (.CI(n49637), .I0(GND_net), .I1(n12209), .CO(n49638));
    SB_LUT4 encoder0_position_30__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n49834), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1972_11 (.CI(n50394), .I0(n2925), 
            .I1(VCC_net), .CO(n50395));
    SB_LUT4 encoder0_position_30__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n50393), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n49833), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_10 (.CI(n50393), .I0(n2926), 
            .I1(VCC_net), .CO(n50394));
    SB_LUT4 encoder0_position_30__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n50392), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_11_lut (.I0(GND_net), .I1(GND_net), .I2(n12211), 
            .I3(n49636), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_9 (.CI(n50392), .I0(n2927), 
            .I1(VCC_net), .CO(n50393));
    SB_LUT4 encoder0_position_30__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n50391), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_8 (.CI(n50391), .I0(n2928), 
            .I1(VCC_net), .CO(n50392));
    SB_CARRY encoder0_position_30__I_0_add_632_8 (.CI(n49833), .I0(n928), 
            .I1(VCC_net), .CO(n49834));
    SB_LUT4 encoder0_position_30__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n50390), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_7 (.CI(n50390), .I0(n2929), 
            .I1(GND_net), .CO(n50391));
    SB_LUT4 encoder0_position_30__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n50389), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_6 (.CI(n50389), .I0(n2930), 
            .I1(GND_net), .CO(n50390));
    SB_LUT4 encoder0_position_30__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n49832), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n50388), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_5 (.CI(n50388), .I0(n2931), 
            .I1(VCC_net), .CO(n50389));
    SB_CARRY encoder0_position_30__I_0_add_632_7 (.CI(n49832), .I0(n929), 
            .I1(GND_net), .CO(n49833));
    SB_LUT4 encoder0_position_30__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n50387), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_4 (.CI(n50387), .I0(n2932), 
            .I1(GND_net), .CO(n50388));
    SB_CARRY add_1097_11 (.CI(n49636), .I0(GND_net), .I1(n12211), .CO(n49637));
    SB_LUT4 encoder0_position_30__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n50386), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_3 (.CI(n50386), .I0(n2933), 
            .I1(VCC_net), .CO(n50387));
    SB_LUT4 encoder0_position_30__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n50386));
    SB_LUT4 encoder0_position_30__I_0_add_1905_28_lut (.I0(n68915), .I1(n2808), 
            .I2(VCC_net), .I3(n50385), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n49831), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_10_lut (.I0(GND_net), .I1(GND_net), .I2(n12213), 
            .I3(n49635), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n50384), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_27 (.CI(n50384), .I0(n2809), 
            .I1(VCC_net), .CO(n50385));
    SB_CARRY encoder0_position_30__I_0_add_632_6 (.CI(n49831), .I0(n930), 
            .I1(GND_net), .CO(n49832));
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n49530), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n50383), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_26 (.CI(n50383), .I0(n2810), 
            .I1(VCC_net), .CO(n50384));
    SB_CARRY add_151_22 (.CI(n49530), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n49531));
    SB_LUT4 encoder0_position_30__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n49830), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_5 (.CI(n49830), .I0(n931), 
            .I1(VCC_net), .CO(n49831));
    SB_LUT4 encoder0_position_30__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n49829), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_10 (.CI(n49635), .I0(GND_net), .I1(n12213), .CO(n49636));
    SB_CARRY encoder0_position_30__I_0_add_632_4 (.CI(n49829), .I0(n932), 
            .I1(GND_net), .CO(n49830));
    SB_LUT4 i42492_3_lut (.I0(n4_adj_5913), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n58169));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i42492_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 encoder0_position_30__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n49828), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_9_lut (.I0(GND_net), .I1(GND_net), .I2(n12215), .I3(n49634), 
            .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_3 (.CI(n49828), .I0(n933), 
            .I1(VCC_net), .CO(n49829));
    SB_CARRY add_1097_9 (.CI(n49634), .I0(GND_net), .I1(n12215), .CO(n49635));
    SB_LUT4 add_1097_8_lut (.I0(GND_net), .I1(GND_net), .I2(n12217), .I3(n49633), 
            .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22496_3_lut (.I0(n219), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [12]));
    defparam i22496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1101_16_lut (.I0(GND_net), .I1(n1620), 
            .I2(VCC_net), .I3(n50030), .O(n1687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n50029), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n50382), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_25 (.CI(n50382), .I0(n2811), 
            .I1(VCC_net), .CO(n50383));
    SB_CARRY encoder0_position_30__I_0_add_1101_15 (.CI(n50029), .I0(n1621), 
            .I1(VCC_net), .CO(n50030));
    SB_LUT4 encoder0_position_30__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n50381), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_24 (.CI(n50381), .I0(n2812), 
            .I1(VCC_net), .CO(n50382));
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n49529), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_2_lut (.I0(GND_net), .I1(n520), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_21 (.CI(n49529), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n49530));
    SB_LUT4 encoder0_position_30__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n50380), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_23 (.CI(n50380), .I0(n2813), 
            .I1(VCC_net), .CO(n50381));
    SB_LUT4 encoder0_position_30__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n50379), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_2 (.CI(VCC_net), .I0(n520), 
            .I1(GND_net), .CO(n49828));
    SB_CARRY encoder0_position_30__I_0_add_1905_22 (.CI(n50379), .I0(n2814), 
            .I1(VCC_net), .CO(n50380));
    SB_LUT4 encoder0_position_30__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n50028), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_14 (.CI(n50028), .I0(n1622), 
            .I1(VCC_net), .CO(n50029));
    SB_LUT4 encoder0_position_30__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n50378), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_21 (.CI(n50378), .I0(n2815), 
            .I1(VCC_net), .CO(n50379));
    SB_LUT4 encoder0_position_30__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n50377), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n50027), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_2108 (.I0(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I1(Ki[0]), .I2(GND_net), .I3(GND_net), .O(n38));
    defparam i1_2_lut_adj_2108.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_1101_13 (.CI(n50027), .I0(n1623), 
            .I1(VCC_net), .CO(n50028));
    SB_CARRY encoder0_position_30__I_0_add_1905_20 (.CI(n50377), .I0(n2816), 
            .I1(VCC_net), .CO(n50378));
    SB_LUT4 encoder0_position_30__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n50376), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_8 (.CI(n49633), .I0(GND_net), .I1(n12217), .CO(n49634));
    SB_CARRY encoder0_position_30__I_0_add_1905_19 (.CI(n50376), .I0(n2817), 
            .I1(VCC_net), .CO(n50377));
    SB_LUT4 encoder0_position_30__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n50375), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_18 (.CI(n50375), .I0(n2818), 
            .I1(VCC_net), .CO(n50376));
    SB_CARRY add_151_9 (.CI(n49517), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n49518));
    SB_LUT4 encoder0_position_30__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n50374), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n50026), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n49528), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_17 (.CI(n50374), .I0(n2819), 
            .I1(VCC_net), .CO(n50375));
    SB_LUT4 encoder0_position_30__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820_adj_5823), 
            .I2(VCC_net), .I3(n50373), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_16 (.CI(n50373), .I0(n2820_adj_5823), 
            .I1(VCC_net), .CO(n50374));
    SB_LUT4 encoder0_position_30__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n50372), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_15 (.CI(n50372), .I0(n2821), 
            .I1(VCC_net), .CO(n50373));
    SB_LUT4 encoder0_position_30__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n50371), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_14 (.CI(n50371), .I0(n2822), 
            .I1(VCC_net), .CO(n50372));
    SB_LUT4 add_1097_7_lut (.I0(GND_net), .I1(GND_net), .I2(n12219), .I3(n49632), 
            .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n50370), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_13 (.CI(n50370), .I0(n2823), 
            .I1(VCC_net), .CO(n50371));
    SB_LUT4 encoder0_position_30__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n50369), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_12 (.CI(n50369), .I0(n2824), 
            .I1(VCC_net), .CO(n50370));
    SB_LUT4 encoder0_position_30__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n50368), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_11 (.CI(n50368), .I0(n2825), 
            .I1(VCC_net), .CO(n50369));
    SB_LUT4 encoder0_position_30__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n50367), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_12 (.CI(n50026), .I0(n1624), 
            .I1(VCC_net), .CO(n50027));
    SB_CARRY add_1097_7 (.CI(n49632), .I0(GND_net), .I1(n12219), .CO(n49633));
    SB_CARRY encoder0_position_30__I_0_add_1905_10 (.CI(n50367), .I0(n2826), 
            .I1(VCC_net), .CO(n50368));
    SB_LUT4 encoder0_position_30__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n50366), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_9 (.CI(n50366), .I0(n2827), 
            .I1(VCC_net), .CO(n50367));
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n49516), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n50365), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_8 (.CI(n50365), .I0(n2828), 
            .I1(VCC_net), .CO(n50366));
    SB_LUT4 encoder0_position_30__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n50364), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_7 (.CI(n50364), .I0(n2829), 
            .I1(GND_net), .CO(n50365));
    SB_LUT4 add_1097_6_lut (.I0(GND_net), .I1(GND_net), .I2(n12221), .I3(n49631), 
            .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_20 (.CI(n49528), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n49529));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n49527), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n50363), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_6 (.CI(n50363), .I0(n2830), 
            .I1(GND_net), .CO(n50364));
    SB_LUT4 encoder0_position_30__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n50362), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n49511), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_5 (.CI(n50362), .I0(n2831), 
            .I1(VCC_net), .CO(n50363));
    SB_CARRY add_1097_6 (.CI(n49631), .I0(GND_net), .I1(n12221), .CO(n49632));
    SB_LUT4 encoder0_position_30__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n50361), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n50025), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_5_lut (.I0(GND_net), .I1(GND_net), .I2(n12223), .I3(n49630), 
            .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15642_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n22792), .I3(GND_net), .O(n29718));   // verilog/coms.v(130[12] 305[6])
    defparam i15642_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1905_4 (.CI(n50361), .I0(n2832), 
            .I1(GND_net), .CO(n50362));
    SB_LUT4 encoder0_position_30__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n50360), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_3 (.CI(n50360), .I0(n2833), 
            .I1(VCC_net), .CO(n50361));
    SB_CARRY add_1097_5 (.CI(n49630), .I0(GND_net), .I1(n12223), .CO(n49631));
    SB_CARRY encoder0_position_30__I_0_add_1101_11 (.CI(n50025), .I0(n1625), 
            .I1(VCC_net), .CO(n50026));
    SB_LUT4 encoder0_position_30__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n50360));
    SB_LUT4 encoder0_position_30__I_0_add_1838_27_lut (.I0(GND_net), .I1(n2709), 
            .I2(VCC_net), .I3(n50359), .O(n2776)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n50024), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_10 (.CI(n50024), .I0(n1626), 
            .I1(VCC_net), .CO(n50025));
    SB_LUT4 add_1097_4_lut (.I0(GND_net), .I1(GND_net), .I2(n12225), .I3(n49629), 
            .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n50358), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_26 (.CI(n50358), .I0(n2710), 
            .I1(VCC_net), .CO(n50359));
    SB_LUT4 encoder0_position_30__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n50357), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n50023), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_9 (.CI(n50023), .I0(n1627), 
            .I1(VCC_net), .CO(n50024));
    SB_CARRY add_151_8 (.CI(n49516), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n49517));
    SB_LUT4 encoder0_position_30__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n50022), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_8 (.CI(n50022), .I0(n1628), 
            .I1(VCC_net), .CO(n50023));
    SB_CARRY add_151_19 (.CI(n49527), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n49528));
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n49526), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_25 (.CI(n50357), .I0(n2711), 
            .I1(VCC_net), .CO(n50358));
    SB_LUT4 encoder0_position_30__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n50021), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n49822), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_151_3 (.CI(n49511), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n49512));
    SB_CARRY encoder0_position_30__I_0_add_1101_7 (.CI(n50021), .I0(n1629), 
            .I1(GND_net), .CO(n50022));
    SB_CARRY add_151_18 (.CI(n49526), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n49527));
    SB_LUT4 encoder0_position_30__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n50020), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n50356), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n49821), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_6 (.CI(n50020), .I0(n1630), 
            .I1(GND_net), .CO(n50021));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n49515), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n49525), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_7 (.CI(n49821), .I0(n829), 
            .I1(GND_net), .CO(n49822));
    SB_CARRY encoder0_position_30__I_0_add_1838_24 (.CI(n50356), .I0(n2712), 
            .I1(VCC_net), .CO(n50357));
    SB_LUT4 encoder0_position_30__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n50355), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n50019), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_7 (.CI(n49515), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n49516));
    SB_CARRY encoder0_position_30__I_0_add_1838_23 (.CI(n50355), .I0(n2713), 
            .I1(VCC_net), .CO(n50356));
    SB_CARRY add_1097_4 (.CI(n49629), .I0(GND_net), .I1(n12225), .CO(n49630));
    SB_LUT4 encoder0_position_30__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n49820), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_5 (.CI(n50019), .I0(n1631), 
            .I1(VCC_net), .CO(n50020));
    SB_CARRY add_151_17 (.CI(n49525), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n49526));
    SB_CARRY encoder0_position_30__I_0_add_565_6 (.CI(n49820), .I0(n830), 
            .I1(GND_net), .CO(n49821));
    SB_LUT4 encoder0_position_30__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n50354), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_3_lut (.I0(GND_net), .I1(GND_net), .I2(n12227), .I3(n49628), 
            .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_3 (.CI(n49628), .I0(GND_net), .I1(n12227), .CO(n49629));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n49524), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_2_lut (.I0(GND_net), .I1(GND_net), .I2(n11642), .I3(VCC_net), 
            .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_22 (.CI(n50354), .I0(n2714), 
            .I1(VCC_net), .CO(n50355));
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n50353), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_16 (.CI(n49524), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n49525));
    SB_LUT4 encoder0_position_30__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n50018), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_21 (.CI(n50353), .I0(n2715), 
            .I1(VCC_net), .CO(n50354));
    SB_LUT4 encoder0_position_30__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n49819), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n50352), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_5 (.CI(n49819), .I0(n831), 
            .I1(VCC_net), .CO(n49820));
    SB_CARRY encoder0_position_30__I_0_add_1838_20 (.CI(n50352), .I0(n2716), 
            .I1(VCC_net), .CO(n50353));
    SB_CARRY encoder0_position_30__I_0_add_1101_4 (.CI(n50018), .I0(n1632), 
            .I1(GND_net), .CO(n50019));
    SB_CARRY add_1097_2 (.CI(VCC_net), .I0(GND_net), .I1(n11642), .CO(n49628));
    SB_LUT4 encoder0_position_30__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n50351), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_19 (.CI(n50351), .I0(n2717), 
            .I1(VCC_net), .CO(n50352));
    SB_LUT4 encoder0_position_30__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n50350), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_18 (.CI(n50350), .I0(n2718), 
            .I1(VCC_net), .CO(n50351));
    SB_LUT4 encoder0_position_30__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n50017), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n50349), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_17 (.CI(n50349), .I0(n2719), 
            .I1(VCC_net), .CO(n50350));
    SB_LUT4 encoder0_position_30__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n50348), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_3 (.CI(n50017), .I0(n1633), 
            .I1(VCC_net), .CO(n50018));
    SB_CARRY encoder0_position_30__I_0_add_1838_16 (.CI(n50348), .I0(n2720), 
            .I1(VCC_net), .CO(n50349));
    SB_LUT4 encoder0_position_30__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n50347), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_15 (.CI(n50347), .I0(n2721), 
            .I1(VCC_net), .CO(n50348));
    SB_LUT4 encoder0_position_30__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n50346), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_14 (.CI(n50346), .I0(n2722), 
            .I1(VCC_net), .CO(n50347));
    SB_LUT4 encoder0_position_30__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n50345), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n50017));
    SB_CARRY encoder0_position_30__I_0_add_1838_13 (.CI(n50345), .I0(n2723), 
            .I1(VCC_net), .CO(n50346));
    SB_LUT4 encoder0_position_30__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n50344), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_12 (.CI(n50344), .I0(n2724), 
            .I1(VCC_net), .CO(n50345));
    SB_LUT4 encoder0_position_30__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n50343), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_11 (.CI(n50343), .I0(n2725), 
            .I1(VCC_net), .CO(n50344));
    SB_LUT4 encoder0_position_30__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n50342), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_10 (.CI(n50342), .I0(n2726), 
            .I1(VCC_net), .CO(n50343));
    SB_LUT4 encoder0_position_30__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n50341), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n49818), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_9 (.CI(n50341), .I0(n2727), 
            .I1(VCC_net), .CO(n50342));
    SB_LUT4 encoder0_position_30__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n50340), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_8 (.CI(n50340), .I0(n2728), 
            .I1(VCC_net), .CO(n50341));
    SB_CARRY encoder0_position_30__I_0_add_565_4 (.CI(n49818), .I0(n832), 
            .I1(GND_net), .CO(n49819));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n49523), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n50339), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_7 (.CI(n50339), .I0(n2729), 
            .I1(GND_net), .CO(n50340));
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n49514), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_15 (.CI(n49523), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n49524));
    SB_LUT4 encoder0_position_30__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n50338), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n49522), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_6 (.CI(n50338), .I0(n2730), 
            .I1(GND_net), .CO(n50339));
    SB_LUT4 encoder0_position_30__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n50337), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_5 (.CI(n50337), .I0(n2731), 
            .I1(VCC_net), .CO(n50338));
    SB_LUT4 encoder0_position_30__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n50336), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n49817), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_4 (.CI(n50336), .I0(n2732), 
            .I1(GND_net), .CO(n50337));
    SB_CARRY add_151_14 (.CI(n49522), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n49523));
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n49511));
    SB_CARRY encoder0_position_30__I_0_add_565_3 (.CI(n49817), .I0(n833), 
            .I1(VCC_net), .CO(n49818));
    SB_LUT4 encoder0_position_30__I_0_add_565_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n49817));
    SB_LUT4 encoder0_position_30__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n50335), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_3 (.CI(n50335), .I0(n2733), 
            .I1(VCC_net), .CO(n50336));
    SB_LUT4 encoder0_position_30__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n50335));
    SB_LUT4 encoder0_position_30__I_0_add_1771_26_lut (.I0(n69063), .I1(n2610), 
            .I2(VCC_net), .I3(n50334), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n50333), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_25 (.CI(n50333), .I0(n2611), 
            .I1(VCC_net), .CO(n50334));
    SB_CARRY add_151_6 (.CI(n49514), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n49515));
    SB_LUT4 encoder0_position_30__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n50332), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_24 (.CI(n50332), .I0(n2612), 
            .I1(VCC_net), .CO(n50333));
    SB_LUT4 encoder0_position_30__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n50331), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_23 (.CI(n50331), .I0(n2613), 
            .I1(VCC_net), .CO(n50332));
    SB_LUT4 encoder0_position_30__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n50330), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_22 (.CI(n50330), .I0(n2614), 
            .I1(VCC_net), .CO(n50331));
    SB_LUT4 encoder0_position_30__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n50329), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47201_3_lut (.I0(n4908), .I1(duty[20]), .I2(n11579), .I3(GND_net), 
            .O(n62929));
    defparam i47201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47203_3_lut (.I0(n62929), .I1(n62927), .I2(n11577), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i47203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47198_3_lut (.I0(n4907), .I1(duty[21]), .I2(n11579), .I3(GND_net), 
            .O(n62926));
    defparam i47198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47200_3_lut (.I0(n62926), .I1(n62927), .I2(n11577), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i47200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2109 (.I0(n2120), .I1(n2121), .I2(n2123), .I3(n2124), 
            .O(n61590));
    defparam i1_4_lut_adj_2109.LUT_INIT = 16'hfffe;
    SB_LUT4 i47199_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n11579), 
            .I3(GND_net), .O(n62927));
    defparam i47199_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1771_21 (.CI(n50329), .I0(n2615), 
            .I1(VCC_net), .CO(n50330));
    SB_LUT4 i47195_3_lut (.I0(n4906), .I1(duty[22]), .I2(n11579), .I3(GND_net), 
            .O(n62923));
    defparam i47195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47197_3_lut (.I0(n62923), .I1(n62927), .I2(n11577), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i47197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n50328), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7219_3_lut (.I0(n4905), .I1(current[15]), .I2(n11577), .I3(GND_net), 
            .O(n20969));
    defparam i7219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7220_3_lut (.I0(n20969), .I1(duty[23]), .I2(n11579), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i7220_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1771_20 (.CI(n50328), .I0(n2616), 
            .I1(VCC_net), .CO(n50329));
    SB_LUT4 encoder0_position_30__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n50327), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2110 (.I0(n2129), .I1(n61580), .I2(n43685), .I3(n2130), 
            .O(n61582));
    defparam i1_4_lut_adj_2110.LUT_INIT = 16'heccc;
    SB_CARRY encoder0_position_30__I_0_add_1771_19 (.CI(n50327), .I0(n2617), 
            .I1(VCC_net), .CO(n50328));
    SB_LUT4 encoder0_position_30__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n50326), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_18 (.CI(n50326), .I0(n2618), 
            .I1(VCC_net), .CO(n50327));
    SB_LUT4 encoder0_position_30__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n50325), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_17 (.CI(n50325), .I0(n2619), 
            .I1(VCC_net), .CO(n50326));
    SB_LUT4 i15742_3_lut_4_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29818));   // verilog/coms.v(130[12] 305[6])
    defparam i15742_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15741_3_lut_4_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29817));   // verilog/coms.v(130[12] 305[6])
    defparam i15741_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i573_3_lut (.I0(n519), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n50324), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15740_3_lut_4_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29816));   // verilog/coms.v(130[12] 305[6])
    defparam i15740_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15739_3_lut_4_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29815));   // verilog/coms.v(130[12] 305[6])
    defparam i15739_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15645_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n22792), .I3(GND_net), .O(n29721));   // verilog/coms.v(130[12] 305[6])
    defparam i15645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15649_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n22792), .I3(GND_net), .O(n29725));   // verilog/coms.v(130[12] 305[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23915_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n22792), .I3(GND_net), .O(n29729));
    defparam i23915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15654_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n22792), .I3(GND_net), .O(n29730));   // verilog/coms.v(130[12] 305[6])
    defparam i15654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15738_3_lut_4_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29814));   // verilog/coms.v(130[12] 305[6])
    defparam i15738_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_1771_16 (.CI(n50324), .I0(n2620), 
            .I1(VCC_net), .CO(n50325));
    SB_LUT4 i15737_3_lut_4_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29813));   // verilog/coms.v(130[12] 305[6])
    defparam i15737_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15736_3_lut_4_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29812));   // verilog/coms.v(130[12] 305[6])
    defparam i15736_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15735_3_lut_4_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29811));   // verilog/coms.v(130[12] 305[6])
    defparam i15735_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n50323), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15734_3_lut_4_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29810));   // verilog/coms.v(130[12] 305[6])
    defparam i15734_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_1771_15 (.CI(n50323), .I0(n2621), 
            .I1(VCC_net), .CO(n50324));
    SB_LUT4 encoder0_position_30__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n50322), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5768));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1771_14 (.CI(n50322), .I0(n2622), 
            .I1(VCC_net), .CO(n50323));
    SB_LUT4 encoder0_position_30__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n50321), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_13 (.CI(n50321), .I0(n2623), 
            .I1(VCC_net), .CO(n50322));
    SB_LUT4 encoder0_position_30__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n50320), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_12 (.CI(n50320), .I0(n2624), 
            .I1(VCC_net), .CO(n50321));
    SB_LUT4 encoder0_position_30__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n50319), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2460_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n49816), 
            .O(n7450)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_11 (.CI(n50319), .I0(n2625), 
            .I1(VCC_net), .CO(n50320));
    SB_LUT4 encoder0_position_30__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n50318), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_10 (.CI(n50318), .I0(n2626), 
            .I1(VCC_net), .CO(n50319));
    SB_LUT4 i1_4_lut_adj_2111 (.I0(n2116), .I1(n2117), .I2(n2119), .I3(n61590), 
            .O(n61596));
    defparam i1_4_lut_adj_2111.LUT_INIT = 16'hfffe;
    SB_LUT4 i15733_3_lut_4_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29809));   // verilog/coms.v(130[12] 305[6])
    defparam i15733_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5769));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n50317), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_9 (.CI(n50317), .I0(n2627), 
            .I1(VCC_net), .CO(n50318));
    SB_LUT4 i15732_3_lut_4_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29808));   // verilog/coms.v(130[12] 305[6])
    defparam i15732_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n50316), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_8 (.CI(n50316), .I0(n2628), 
            .I1(VCC_net), .CO(n50317));
    SB_LUT4 i15731_3_lut_4_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29807));   // verilog/coms.v(130[12] 305[6])
    defparam i15731_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n50315), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_7 (.CI(n50315), .I0(n2629), 
            .I1(GND_net), .CO(n50316));
    SB_LUT4 encoder0_position_30__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n50314), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_6 (.CI(n50314), .I0(n2630), 
            .I1(GND_net), .CO(n50315));
    SB_LUT4 i15729_3_lut_4_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29805));   // verilog/coms.v(130[12] 305[6])
    defparam i15729_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n50313), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_5 (.CI(n50313), .I0(n2631), 
            .I1(VCC_net), .CO(n50314));
    SB_LUT4 add_2460_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n49815), 
            .O(n7451)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2460_6 (.CI(n49815), .I0(n622), .I1(GND_net), .CO(n49816));
    SB_LUT4 encoder0_position_30__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n50312), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_4 (.CI(n50312), .I0(n2632), 
            .I1(GND_net), .CO(n50313));
    SB_LUT4 encoder0_position_30__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n50311), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_3 (.CI(n50311), .I0(n2633), 
            .I1(VCC_net), .CO(n50312));
    SB_LUT4 encoder0_position_30__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2460_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n49814), 
            .O(n7452)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n50311));
    SB_LUT4 encoder0_position_30__I_0_add_1704_25_lut (.I0(n69034), .I1(n2511), 
            .I2(VCC_net), .I3(n50310), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n50309), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_24 (.CI(n50309), .I0(n2512), 
            .I1(VCC_net), .CO(n50310));
    SB_LUT4 encoder0_position_30__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n50308), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_23 (.CI(n50308), .I0(n2513), 
            .I1(VCC_net), .CO(n50309));
    SB_CARRY add_2460_5 (.CI(n49814), .I0(n623), .I1(VCC_net), .CO(n49815));
    SB_LUT4 encoder0_position_30__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n50307), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_22 (.CI(n50307), .I0(n2514), 
            .I1(VCC_net), .CO(n50308));
    SB_LUT4 encoder0_position_30__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n50306), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2460_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n49813), 
            .O(n7453)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_21 (.CI(n50306), .I0(n2515), 
            .I1(VCC_net), .CO(n50307));
    SB_LUT4 encoder0_position_30__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n50305), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2460_4 (.CI(n49813), .I0(n516), .I1(GND_net), .CO(n49814));
    SB_CARRY encoder0_position_30__I_0_add_1704_20 (.CI(n50305), .I0(n2516), 
            .I1(VCC_net), .CO(n50306));
    SB_LUT4 encoder0_position_30__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n50304), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_19 (.CI(n50304), .I0(n2517), 
            .I1(VCC_net), .CO(n50305));
    SB_LUT4 encoder0_position_30__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n50303), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_18 (.CI(n50303), .I0(n2518), 
            .I1(VCC_net), .CO(n50304));
    SB_LUT4 encoder0_position_30__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n50302), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_17 (.CI(n50302), .I0(n2519), 
            .I1(VCC_net), .CO(n50303));
    SB_LUT4 add_2460_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n49812), 
            .O(n7454)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n50301), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_16 (.CI(n50301), .I0(n2520), 
            .I1(VCC_net), .CO(n50302));
    SB_LUT4 encoder0_position_30__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n50300), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53410_4_lut (.I0(n2118), .I1(n61596), .I2(n61582), .I3(n2115), 
            .O(n2148));
    defparam i53410_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_30__I_0_add_1704_15 (.CI(n50300), .I0(n2521), 
            .I1(VCC_net), .CO(n50301));
    SB_LUT4 encoder0_position_30__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n50299), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_14 (.CI(n50299), .I0(n2522), 
            .I1(VCC_net), .CO(n50300));
    SB_LUT4 encoder0_position_30__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n50298), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_13 (.CI(n50298), .I0(n2523), 
            .I1(VCC_net), .CO(n50299));
    SB_LUT4 encoder0_position_30__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n50297), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_12 (.CI(n50297), .I0(n2524), 
            .I1(VCC_net), .CO(n50298));
    SB_CARRY add_2460_3 (.CI(n49812), .I0(n625), .I1(VCC_net), .CO(n49813));
    SB_LUT4 encoder0_position_30__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n50296), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_11 (.CI(n50296), .I0(n2525), 
            .I1(VCC_net), .CO(n50297));
    SB_LUT4 encoder0_position_30__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n50295), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_10 (.CI(n50295), .I0(n2526), 
            .I1(VCC_net), .CO(n50296));
    SB_LUT4 encoder0_position_30__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n50294), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2460_2_lut (.I0(GND_net), .I1(n518), .I2(GND_net), .I3(VCC_net), 
            .O(n7455)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_9 (.CI(n50294), .I0(n2527), 
            .I1(VCC_net), .CO(n50295));
    SB_CARRY add_2460_2 (.CI(VCC_net), .I0(n518), .I1(GND_net), .CO(n49812));
    SB_LUT4 encoder0_position_30__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n50293), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_8 (.CI(n50293), .I0(n2528), 
            .I1(VCC_net), .CO(n50294));
    SB_LUT4 encoder0_position_30__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n50292), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_7 (.CI(n50292), .I0(n2529), 
            .I1(GND_net), .CO(n50293));
    SB_LUT4 encoder0_position_30__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n50291), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28745_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i28745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28868_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i28868_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_1704_6 (.CI(n50291), .I0(n2530), 
            .I1(GND_net), .CO(n50292));
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n60507));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i15662_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n22792), .I3(GND_net), .O(n29738));   // verilog/coms.v(130[12] 305[6])
    defparam i15662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29640_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n43615));
    defparam i29640_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n50290), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50242_2_lut (.I0(n69808), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65564));
    defparam i50242_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY encoder0_position_30__I_0_add_1704_5 (.CI(n50290), .I0(n2531), 
            .I1(VCC_net), .CO(n50291));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5770));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15432_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n22792), .I3(GND_net), .O(n29508));   // verilog/coms.v(130[12] 305[6])
    defparam i15432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53727_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5924));
    defparam i53727_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 i15669_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n22792), .I3(GND_net), .O(n29745));   // verilog/coms.v(130[12] 305[6])
    defparam i15669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15670_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n22792), .I3(GND_net), .O(n29746));   // verilog/coms.v(130[12] 305[6])
    defparam i15670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15434_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n22792), .I3(GND_net), .O(n29510));   // verilog/coms.v(130[12] 305[6])
    defparam i15434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15671_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n22792), .I3(GND_net), .O(n29747));   // verilog/coms.v(130[12] 305[6])
    defparam i15671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15672_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n22792), .I3(GND_net), .O(n29748));   // verilog/coms.v(130[12] 305[6])
    defparam i15672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15673_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n22792), .I3(GND_net), .O(n29749));   // verilog/coms.v(130[12] 305[6])
    defparam i15673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15674_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n22792), .I3(GND_net), .O(n29750));   // verilog/coms.v(130[12] 305[6])
    defparam i15674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15676_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n22792), .I3(GND_net), .O(n29752));   // verilog/coms.v(130[12] 305[6])
    defparam i15676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15677_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n22792), .I3(GND_net), .O(n29753));   // verilog/coms.v(130[12] 305[6])
    defparam i15677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15678_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n22792), .I3(GND_net), .O(n29754));   // verilog/coms.v(130[12] 305[6])
    defparam i15678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15121_2_lut_3_lut (.I0(n22917), .I1(dti), .I2(n15_adj_5743), 
            .I3(GND_net), .O(n29192));
    defparam i15121_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_2_lut_3_lut_adj_2112 (.I0(n22917), .I1(dti), .I2(n15_adj_5743), 
            .I3(GND_net), .O(n27810));
    defparam i1_2_lut_3_lut_adj_2112.LUT_INIT = 16'hf8f8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5775));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15684_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n22792), .I3(GND_net), .O(n29760));   // verilog/coms.v(130[12] 305[6])
    defparam i15684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29430_2_lut_3_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57410), .I3(n8_adj_5757), .O(n43400));
    defparam i29430_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5777));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29428_2_lut_3_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57410), .I3(n8_adj_5774), .O(n43398));
    defparam i29428_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29426_2_lut_3_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57410), .I3(n8_adj_5801), .O(n43396));
    defparam i29426_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15691_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29767));   // verilog/coms.v(130[12] 305[6])
    defparam i15691_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_3_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n33801), .I3(GND_net), .O(n22792));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5778));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47426_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63154));
    defparam i47426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47427_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63155));
    defparam i47427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230_adj_5808));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47280_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63008));
    defparam i47280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47279_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n63007));
    defparam i47279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15675_3_lut_4_lut (.I0(n1742), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3827), .O(n29751));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15675_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_4_lut_4_lut_adj_2113 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n42725), .O(n55740));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_4_lut_4_lut_adj_2113.LUT_INIT = 16'hb1f1;
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5779));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15655_3_lut_4_lut (.I0(n1784), .I1(b_prev_adj_5753), .I2(a_new_adj_5965[1]), 
            .I3(position_31__N_3827_adj_5754), .O(n29731));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15655_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_2_lut_adj_2114 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n57317));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_2114.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_2115 (.I0(n2222), .I1(n2224), .I2(n2225), .I3(n2228), 
            .O(n61822));
    defparam i1_4_lut_adj_2115.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2116 (.I0(n2227), .I1(n61822), .I2(n2226), .I3(n2223), 
            .O(n61824));
    defparam i1_4_lut_adj_2116.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i841_3_lut (.I0(n1230_adj_5808), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2117 (.I0(n2229), .I1(n43615), .I2(n2230), .I3(n2231), 
            .O(n59100));
    defparam i1_4_lut_adj_2117.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2118 (.I0(n2219), .I1(n2220), .I2(n2221), .I3(n61824), 
            .O(n61830));
    defparam i1_4_lut_adj_2118.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i27_3_lut (.I0(encoder0_position[26]), .I1(n6_adj_5723), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15720_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n61170), 
            .I3(n27_adj_5825), .O(n29796));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15720_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_4310_i28_3_lut (.I0(encoder0_position[27]), .I1(n5_adj_5725), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2119 (.I0(n2217), .I1(n2218), .I2(n61830), .I3(n59100), 
            .O(n61836));
    defparam i1_4_lut_adj_2119.LUT_INIT = 16'hfffe;
    SB_LUT4 i15721_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n61154), 
            .I3(n27_adj_5825), .O(n29797));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15721_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_4310_i29_3_lut (.I0(encoder0_position[28]), .I1(n4_adj_5730), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53435_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n61836), 
            .O(n2247));
    defparam i53435_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_4310_i30_3_lut (.I0(encoder0_position[29]), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15722_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n61090), 
            .I3(n27_adj_5825), .O(n29798));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15722_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6055_2_lut (.I0(n2_adj_5731), .I1(encoder0_position[30]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i6055_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_245_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1086_i15_2_lut (.I0(r_Clock_Count_adj_5997[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5843));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1086_i9_2_lut (.I0(r_Clock_Count_adj_5997[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5840));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1086_i13_2_lut (.I0(r_Clock_Count_adj_5997[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5842));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_1086_i11_2_lut (.I0(r_Clock_Count_adj_5997[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5841));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15614_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5996[1]), 
            .I2(r_SM_Main_adj_5996[2]), .I3(n6_adj_5893), .O(n29690));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i15614_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i28746_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i28746_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15460_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n22792), .I3(GND_net), .O(n29536));   // verilog/coms.v(130[12] 305[6])
    defparam i15460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15597_3_lut_4_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29673));   // verilog/coms.v(130[12] 305[6])
    defparam i15597_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_1584_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n11642));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1584_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n12227));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_3_lut_adj_2120 (.I0(n5_adj_5895), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n61788));
    defparam i1_3_lut_adj_2120.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_30__I_0_i500_4_lut (.I0(n2_adj_5731), .I1(n7450), 
            .I2(n61788), .I3(encoder0_position[30]), .O(n828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 mux_1584_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n12225));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_2121 (.I0(n36888), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n125));
    defparam i1_2_lut_adj_2121.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_2122 (.I0(n36852), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_2122.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1584_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n12223));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_2123 (.I0(n36888), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n198));
    defparam i1_2_lut_adj_2123.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_2124 (.I0(n36888), .I1(Ki[3]), .I2(GND_net), 
            .I3(GND_net), .O(n271));
    defparam i1_2_lut_adj_2124.LUT_INIT = 16'h8888;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15585_3_lut_4_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29661));   // verilog/coms.v(130[12] 305[6])
    defparam i15585_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15584_3_lut_4_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29660));   // verilog/coms.v(130[12] 305[6])
    defparam i15584_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 LessThan_1086_i4_4_lut (.I0(r_Clock_Count_adj_5997[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5997[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5837));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i1_3_lut_adj_2125 (.I0(n2326), .I1(n2324), .I2(n2325), .I3(GND_net), 
            .O(n61614));
    defparam i1_3_lut_adj_2125.LUT_INIT = 16'hfefe;
    SB_LUT4 i52218_3_lut (.I0(n4_adj_5837), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5841), 
            .I3(GND_net), .O(n67946));   // verilog/uart_tx.v(117[17:57])
    defparam i52218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52219_3_lut (.I0(n67946), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5842), 
            .I3(GND_net), .O(n67947));   // verilog/uart_tx.v(117[17:57])
    defparam i52219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51630_4_lut (.I0(n13_adj_5842), .I1(n11_adj_5841), .I2(n9_adj_5840), 
            .I3(n66470), .O(n67358));
    defparam i51630_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1086_i8_3_lut (.I0(n6_adj_5838), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5840), .I3(GND_net), .O(n8_adj_5839));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51209_3_lut (.I0(n67947), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5843), 
            .I3(GND_net), .O(n66937));   // verilog/uart_tx.v(117[17:57])
    defparam i51209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52206_4_lut (.I0(n66937), .I1(n8_adj_5839), .I2(n15_adj_5843), 
            .I3(n67358), .O(n67934));   // verilog/uart_tx.v(117[17:57])
    defparam i52206_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52207_3_lut (.I0(n67934), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5997[8]), 
            .I3(GND_net), .O(n4940));   // verilog/uart_tx.v(117[17:57])
    defparam i52207_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_1584_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n12221));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_2126 (.I0(n36888), .I1(Ki[4]), .I2(GND_net), 
            .I3(GND_net), .O(n344));
    defparam i1_2_lut_adj_2126.LUT_INIT = 16'h8888;
    SB_LUT4 i42620_2_lut (.I0(r_SM_Main_adj_5996[2]), .I1(r_SM_Main_adj_5996[0]), 
            .I2(GND_net), .I3(GND_net), .O(n58304));
    defparam i42620_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15568_3_lut_4_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29644));   // verilog/coms.v(130[12] 305[6])
    defparam i15568_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_1584_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n12219));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5780));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5791));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_2127 (.I0(n36888), .I1(Ki[5]), .I2(GND_net), 
            .I3(GND_net), .O(n417));
    defparam i1_2_lut_adj_2127.LUT_INIT = 16'h8888;
    SB_LUT4 i16154_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n61074), 
            .I3(n27_adj_5825), .O(n30230));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16154_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16155_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n61122), 
            .I3(n27_adj_5825), .O(n30231));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16155_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1237_3_lut (.I0(n1818), .I1(n1885), 
            .I2(n1851), .I3(GND_net), .O(n1917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_2128 (.I0(\data_in_frame[19] [6]), .I1(n28409), 
            .I2(n28464), .I3(rx_data[6]), .O(n56534));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2128.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_2129 (.I0(\data_in_frame[19] [5]), .I1(n31_adj_5822), 
            .I2(n28464), .I3(n57340), .O(n56536));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2129.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2130 (.I0(\data_in_frame[19] [4]), .I1(n28409), 
            .I2(n28464), .I3(rx_data[4]), .O(n56538));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2130.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15518_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n28464), .I3(GND_net), .O(n29594));   // verilog/coms.v(130[12] 305[6])
    defparam i15518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1083_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5836));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_2131 (.I0(rx_data[5]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57410), .I3(GND_net), .O(n57340));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_2131.LUT_INIT = 16'h0202;
    SB_LUT4 i12_4_lut_adj_2132 (.I0(\data_in_frame[19] [2]), .I1(n28409), 
            .I2(n28464), .I3(rx_data[2]), .O(n56540));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2132.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_1083_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5833));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i16164_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[1]), 
            .I2(n10_adj_5892), .I3(n25595), .O(n30240));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16164_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16165_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[2]), 
            .I2(n4_adj_5745), .I3(n25600), .O(n30241));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16165_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_adj_2133 (.I0(n2323), .I1(n2327), .I2(n2328), .I3(GND_net), 
            .O(n61616));
    defparam i1_3_lut_adj_2133.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_1083_i8_3_lut (.I0(n6_adj_5834), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5836), .I3(GND_net), .O(n8_adj_5835));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16166_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[3]), 
            .I2(n4_adj_5745), .I3(n25595), .O(n30242));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16166_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16167_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[4]), 
            .I2(n4_adj_5746), .I3(n25600), .O(n30243));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16167_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52631_4_lut (.I0(n8_adj_5835), .I1(n4_adj_5833), .I2(n9_adj_5836), 
            .I3(n66483), .O(n68359));   // verilog/uart_rx.v(119[17:57])
    defparam i52631_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_2134 (.I0(n36888), .I1(Ki[6]), .I2(GND_net), 
            .I3(GND_net), .O(n490));
    defparam i1_2_lut_adj_2134.LUT_INIT = 16'h8888;
    SB_LUT4 i16168_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[5]), 
            .I2(n4_adj_5746), .I3(n25595), .O(n30244));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16168_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52632_3_lut (.I0(n68359), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n68360));   // verilog/uart_rx.v(119[17:57])
    defparam i52632_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16169_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[6]), 
            .I2(n42890), .I3(n25600), .O(n30245));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16169_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i52512_3_lut (.I0(n68360), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n68240));   // verilog/uart_rx.v(119[17:57])
    defparam i52512_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51207_3_lut (.I0(n68240), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4937));   // verilog/uart_rx.v(119[17:57])
    defparam i51207_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16170_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5978[7]), 
            .I2(n42890), .I3(n25595), .O(n30246));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16170_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5792));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2135 (.I0(state[0]), .I1(n23_adj_5922), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5832));
    defparam i1_2_lut_adj_2135.LUT_INIT = 16'h2222;
    SB_LUT4 i13_4_lut_adj_2136 (.I0(n111), .I1(n43567), .I2(state[1]), 
            .I3(n4_adj_5832), .O(n5_adj_5902));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13_4_lut_adj_2136.LUT_INIT = 16'hcafa;
    SB_LUT4 i12_4_lut_adj_2137 (.I0(\data_in_frame[19] [1]), .I1(n28409), 
            .I2(n28464), .I3(rx_data[1]), .O(n56542));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2137.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_4_lut_adj_2138 (.I0(control_mode[3]), .I1(control_mode[4]), 
            .I2(control_mode[2]), .I3(control_mode[6]), .O(n62220));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_4_lut_adj_2138.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2139 (.I0(n62220), .I1(control_mode[7]), .I2(control_mode[5]), 
            .I3(GND_net), .O(n25564));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_3_lut_adj_2139.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_2140 (.I0(n25465), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_adj_2140.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_adj_2141 (.I0(control_mode[0]), .I1(n25564), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5701));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut_adj_2141.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_4_lut_adj_2142 (.I0(\data_in_frame[19] [0]), .I1(n28409), 
            .I2(n28464), .I3(rx_data[0]), .O(n56546));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2142.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13_4_lut_adj_2143 (.I0(\data_in_frame[18] [7]), .I1(n8_adj_5757), 
            .I2(n43400), .I3(n57336), .O(n56430));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2143.LUT_INIT = 16'ha3a0;
    SB_LUT4 i13_4_lut_adj_2144 (.I0(\data_in_frame[18] [6]), .I1(n58292), 
            .I2(n43400), .I3(rx_data[6]), .O(n56434));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2144.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5793));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15500_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n43400), .I3(GND_net), .O(n29576));   // verilog/coms.v(130[12] 305[6])
    defparam i15500_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5794));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15497_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n43400), .I3(GND_net), .O(n29573));   // verilog/coms.v(130[12] 305[6])
    defparam i15497_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15494_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n43400), .I3(GND_net), .O(n29570));   // verilog/coms.v(130[12] 305[6])
    defparam i15494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_2145 (.I0(\data_in_frame[18] [2]), .I1(n58292), 
            .I2(n43400), .I3(rx_data[2]), .O(n56438));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2145.LUT_INIT = 16'ha3a0;
    SB_LUT4 i13_4_lut_adj_2146 (.I0(\data_in_frame[18] [1]), .I1(n58292), 
            .I2(n43400), .I3(rx_data[1]), .O(n56442));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2146.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5795));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47071_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n62790));
    defparam i47071_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53667_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6617), .I2(n62790), 
            .I3(n25_adj_5898), .O(n17_adj_5897));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i53667_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 mux_4310_i8_3_lut (.I0(encoder0_position[7]), .I1(n25_adj_5706), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_1584_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n12217));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_1584_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n12215));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5796));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29638_3_lut (.I0(n948), .I1(n2332), .I2(n2333), .I3(GND_net), 
            .O(n43613));
    defparam i29638_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_i1176_3_lut (.I0(n1725), .I1(n1792_adj_5815), 
            .I2(n1752), .I3(GND_net), .O(n1824_adj_5819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2147 (.I0(n2321), .I1(n2322), .I2(n61616), .I3(n61614), 
            .O(n61622));
    defparam i1_4_lut_adj_2147.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1243_3_lut (.I0(n1824_adj_5819), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2148 (.I0(n2329), .I1(n43613), .I2(n2330), .I3(n2331), 
            .O(n59080));
    defparam i1_4_lut_adj_2148.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16127_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n58278), .I3(GND_net), .O(n30203));   // verilog/coms.v(130[12] 305[6])
    defparam i16127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16123_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n58278), .I3(GND_net), .O(n30199));   // verilog/coms.v(130[12] 305[6])
    defparam i16123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_2149 (.I0(\data_in_frame[22] [3]), .I1(n58294), 
            .I2(n43396), .I3(rx_data[3]), .O(n56410));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2149.LUT_INIT = 16'ha3a0;
    SB_LUT4 i16120_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n58278), .I3(GND_net), .O(n30196));   // verilog/coms.v(130[12] 305[6])
    defparam i16120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52889_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[12] [4]), 
            .I2(n58278), .I3(GND_net), .O(n56690));   // verilog/coms.v(94[13:20])
    defparam i52889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1584_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n12213));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i52886_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[12] [3]), 
            .I2(n58278), .I3(GND_net), .O(n56636));   // verilog/coms.v(94[13:20])
    defparam i52886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16110_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n58278), .I3(GND_net), .O(n30186));   // verilog/coms.v(130[12] 305[6])
    defparam i16110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15625_3_lut (.I0(\data_in_frame[0] [1]), .I1(rx_data[1]), .I2(n7_adj_5921), 
            .I3(GND_net), .O(n29701));   // verilog/coms.v(130[12] 305[6])
    defparam i15625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16473_3_lut_4_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30549));   // verilog/coms.v(130[12] 305[6])
    defparam i16473_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16107_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n58278), .I3(GND_net), .O(n30183));   // verilog/coms.v(130[12] 305[6])
    defparam i16107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16472_3_lut_4_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30548));   // verilog/coms.v(130[12] 305[6])
    defparam i16472_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16471_3_lut_4_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30547));   // verilog/coms.v(130[12] 305[6])
    defparam i16471_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16470_3_lut_4_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30546));   // verilog/coms.v(130[12] 305[6])
    defparam i16470_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16104_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n58278), .I3(GND_net), .O(n30180));   // verilog/coms.v(130[12] 305[6])
    defparam i16104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16101_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n30177));   // verilog/coms.v(130[12] 305[6])
    defparam i16101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16469_3_lut_4_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30545));   // verilog/coms.v(130[12] 305[6])
    defparam i16469_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16468_3_lut_4_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30544));   // verilog/coms.v(130[12] 305[6])
    defparam i16468_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16097_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n30173));   // verilog/coms.v(130[12] 305[6])
    defparam i16097_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16094_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n30170));   // verilog/coms.v(130[12] 305[6])
    defparam i16094_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16091_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n30167));   // verilog/coms.v(130[12] 305[6])
    defparam i16091_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52885_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[11] [3]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n56604));   // verilog/coms.v(94[13:20])
    defparam i52885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52888_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[11] [2]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n56678));   // verilog/coms.v(94[13:20])
    defparam i52888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52887_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[11] [1]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n56662));   // verilog/coms.v(94[13:20])
    defparam i52887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16078_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n7_adj_5920), .I3(GND_net), .O(n30154));   // verilog/coms.v(130[12] 305[6])
    defparam i16078_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5727));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1584_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n12211));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16075_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n57424), .I3(GND_net), .O(n30151));   // verilog/coms.v(130[12] 305[6])
    defparam i16075_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16072_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n57424), .I3(GND_net), .O(n30148));   // verilog/coms.v(130[12] 305[6])
    defparam i16072_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16068_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n57424), .I3(GND_net), .O(n30144));   // verilog/coms.v(130[12] 305[6])
    defparam i16068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1584_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n12209));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16065_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n57424), .I3(GND_net), .O(n30141));   // verilog/coms.v(130[12] 305[6])
    defparam i16065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16062_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n57424), .I3(GND_net), .O(n30138));   // verilog/coms.v(130[12] 305[6])
    defparam i16062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16058_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n57424), .I3(GND_net), .O(n30134));   // verilog/coms.v(130[12] 305[6])
    defparam i16058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16055_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n57424), .I3(GND_net), .O(n30131));   // verilog/coms.v(130[12] 305[6])
    defparam i16055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16467_3_lut_4_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30543));   // verilog/coms.v(130[12] 305[6])
    defparam i16467_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5677));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16049_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n57426), 
            .I3(GND_net), .O(n30125));   // verilog/coms.v(130[12] 305[6])
    defparam i16049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16046_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n57426), 
            .I3(GND_net), .O(n30122));   // verilog/coms.v(130[12] 305[6])
    defparam i16046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5678));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16042_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n57426), 
            .I3(GND_net), .O(n30118));   // verilog/coms.v(130[12] 305[6])
    defparam i16042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5799));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1584_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n12207));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16039_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n57426), 
            .I3(GND_net), .O(n30115));   // verilog/coms.v(130[12] 305[6])
    defparam i16039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5680));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50792_4_lut (.I0(n11), .I1(n9), .I2(n7_adj_5678), .I3(n5_adj_5680), 
            .O(n66520));
    defparam i50792_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16036_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n57426), 
            .I3(GND_net), .O(n30112));   // verilog/coms.v(130[12] 305[6])
    defparam i16036_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16032_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n57426), 
            .I3(GND_net), .O(n30108));   // verilog/coms.v(130[12] 305[6])
    defparam i16032_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16029_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n57426), 
            .I3(GND_net), .O(n30105));   // verilog/coms.v(130[12] 305[6])
    defparam i16029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8), .I1(current_limit[9]), .I2(n19), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5681));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i16026_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n57426), 
            .I3(GND_net), .O(n30102));   // verilog/coms.v(130[12] 305[6])
    defparam i16026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52126_3_lut (.I0(n4_adj_5681), .I1(current_limit[5]), .I2(n11), 
            .I3(GND_net), .O(n67854));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52127_3_lut (.I0(n67854), .I1(current_limit[6]), .I2(n13), 
            .I3(GND_net), .O(n67855));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2150 (.I0(n2319), .I1(n59080), .I2(n2320), .I3(n61622), 
            .O(n61628));
    defparam i1_4_lut_adj_2150.LUT_INIT = 16'hfffe;
    SB_LUT4 i50782_4_lut (.I0(n17), .I1(n15_adj_5677), .I2(n13), .I3(n66520), 
            .O(n66510));
    defparam i50782_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52658_4_lut (.I0(n16), .I1(n6_adj_5679), .I2(n19), .I3(n66508), 
            .O(n68386));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52658_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_1584_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n12205));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16023_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n58317), 
            .I3(GND_net), .O(n30099));   // verilog/coms.v(130[12] 305[6])
    defparam i16023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16020_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n58317), 
            .I3(GND_net), .O(n30096));   // verilog/coms.v(130[12] 305[6])
    defparam i16020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16017_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n58317), 
            .I3(GND_net), .O(n30093));   // verilog/coms.v(130[12] 305[6])
    defparam i16017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut_adj_2151 (.I0(data_ready), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5912));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i2_3_lut_4_lut_adj_2151.LUT_INIT = 16'h080c;
    SB_LUT4 i1855_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42725), .O(n6617));   // verilog/TinyFPGA_B.v(361[5] 387[12])
    defparam i1855_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5701), .I3(n15), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_2152 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42725), .O(n24_adj_5896));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_adj_2152.LUT_INIT = 16'hffbf;
    SB_LUT4 i51036_3_lut (.I0(n67855), .I1(current_limit[7]), .I2(n15_adj_5677), 
            .I3(GND_net), .O(n66764));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52819_4_lut (.I0(n66764), .I1(n68386), .I2(n19), .I3(n66510), 
            .O(n68547));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52819_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i23914_3_lut (.I0(n58317), .I1(rx_data[4]), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n30314));   // verilog/coms.v(94[13:20])
    defparam i23914_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i52820_3_lut (.I0(n68547), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n68548));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52820_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52745_3_lut (.I0(n68548), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n68473));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52745_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_14_i26_3_lut (.I0(n68473), .I1(current_limit[12]), 
            .I2(current[15]), .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16011_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n58317), 
            .I3(GND_net), .O(n30087));   // verilog/coms.v(130[12] 305[6])
    defparam i16011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2153 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n61628), 
            .O(n61634));
    defparam i1_4_lut_adj_2153.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53249_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n61634), 
            .O(n2346));
    defparam i53249_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i50926_2_lut_3_lut (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(state_adj_5979[1]), .I3(GND_net), .O(n65782));   // verilog/eeprom.v(35[8] 81[4])
    defparam i50926_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5740));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1584_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n12203));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15923_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29999));
    defparam i15923_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15900_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29976));
    defparam i15900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16007_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n58317), 
            .I3(GND_net), .O(n30083));   // verilog/coms.v(130[12] 305[6])
    defparam i16007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15903_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29979));
    defparam i15903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15907_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29983));
    defparam i15907_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16004_3_lut (.I0(\data_in_frame[8] [1]), .I1(rx_data[1]), .I2(n58317), 
            .I3(GND_net), .O(n30080));   // verilog/coms.v(130[12] 305[6])
    defparam i16004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42633_3_lut (.I0(reset), .I1(n8_adj_5776), .I2(n57437), .I3(GND_net), 
            .O(n58317));
    defparam i42633_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5738));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16001_3_lut (.I0(\data_in_frame[8] [0]), .I1(rx_data[0]), .I2(n58317), 
            .I3(GND_net), .O(n30077));   // verilog/coms.v(130[12] 305[6])
    defparam i16001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5732));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_2154 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5899));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_2154.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5729));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15910_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29986));
    defparam i15910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15913_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29989));
    defparam i15913_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut (.I0(commutation_state[0]), .I1(n4_adj_5899), .I2(commutation_state_prev[0]), 
            .I3(GND_net), .O(n15_adj_5743));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i2_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i15992_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n7_adj_5917), 
            .I3(GND_net), .O(n30068));   // verilog/coms.v(130[12] 305[6])
    defparam i15992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15989_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n7_adj_5917), 
            .I3(GND_net), .O(n30065));   // verilog/coms.v(130[12] 305[6])
    defparam i15989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5728));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15986_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n7_adj_5917), 
            .I3(GND_net), .O(n30062));   // verilog/coms.v(130[12] 305[6])
    defparam i15986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i24_3_lut (.I0(encoder0_position[23]), .I1(n9_adj_5720), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5736));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15983_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n7_adj_5917), 
            .I3(GND_net), .O(n30059));   // verilog/coms.v(130[12] 305[6])
    defparam i15983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5735));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i641_3_lut (.I0(n520), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15979_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n7_adj_5917), 
            .I3(GND_net), .O(n30055));   // verilog/coms.v(130[12] 305[6])
    defparam i15979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5734));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27754), .O(n53222));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 encoder0_position_30__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5698));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5685));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231_adj_5809));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5682));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5686));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i842_3_lut (.I0(n1231_adj_5809), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5703));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_6010[0]), .I1(n65775), .I2(n6428), 
            .I3(n10_adj_5747), .O(n8_adj_5918));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 mux_1584_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n12201));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16428_3_lut_4_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30504));   // verilog/coms.v(130[12] 305[6])
    defparam i16428_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i2_2_lut_adj_2155 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5905));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut_adj_2155.LUT_INIT = 16'heeee;
    SB_LUT4 i16427_3_lut_4_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30503));   // verilog/coms.v(130[12] 305[6])
    defparam i16427_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16424_3_lut_4_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30500));   // verilog/coms.v(130[12] 305[6])
    defparam i16424_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1584_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n12199));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5771));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_4_lut_adj_2156 (.I0(\data_in_frame[18] [0]), .I1(n58292), 
            .I2(n43400), .I3(rx_data[0]), .O(n56446));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2156.LUT_INIT = 16'ha3a0;
    SB_LUT4 i13_4_lut_adj_2157 (.I0(\data_in_frame[17] [7]), .I1(n8_adj_5774), 
            .I2(n43398), .I3(n57336), .O(n56450));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2157.LUT_INIT = 16'ha3a0;
    SB_LUT4 i13_4_lut_adj_2158 (.I0(\data_in_frame[17] [6]), .I1(n58290), 
            .I2(n43398), .I3(rx_data[6]), .O(n56454));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2158.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_30__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5702));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n65589), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16266_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30342));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16267_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n57425), .I3(GND_net), .O(n30343));   // verilog/coms.v(130[12] 305[6])
    defparam i16267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_2159 (.I0(\data_in_frame[17] [5]), .I1(n8_adj_5774), 
            .I2(n43398), .I3(n57340), .O(n56458));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2159.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5772));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52339_3_lut (.I0(n4), .I1(n305), .I2(n11_adj_5702), .I3(GND_net), 
            .O(n68067));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52340_3_lut (.I0(n68067), .I1(n304), .I2(n13_adj_5703), .I3(GND_net), 
            .O(n68068));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16423_3_lut_4_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30499));   // verilog/coms.v(130[12] 305[6])
    defparam i16423_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_1584_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n12197));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16271_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30347));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16272_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30348));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16273_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30349));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16274_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30350));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1584_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n12195));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16275_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30351));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5773));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16276_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30352));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16277_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30353));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16278_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30354));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16279_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30355));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16279_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16422_3_lut_4_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30498));   // verilog/coms.v(130[12] 305[6])
    defparam i16422_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_1584_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n12193));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1584_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n12191));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16414_3_lut_4_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30490));   // verilog/coms.v(130[12] 305[6])
    defparam i16414_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_1584_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n12189));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1584_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n12187));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1103_3_lut (.I0(n1620), .I1(n1687), 
            .I2(n1653), .I3(GND_net), .O(n1719));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17_adj_5686), 
            .I3(GND_net), .O(n8_adj_5683));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_2160 (.I0(\data_in_frame[17] [3]), .I1(n58290), 
            .I2(n43398), .I3(rx_data[3]), .O(n56466));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2160.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_30__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_2161 (.I0(\data_in_frame[17] [2]), .I1(n58290), 
            .I2(n43398), .I3(rx_data[2]), .O(n56470));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2161.LUT_INIT = 16'ha3a0;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5697));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7), .I3(GND_net), 
            .O(n6_adj_5676));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5683), .I1(n301), .I2(n19_adj_5685), 
            .I3(GND_net), .O(n16_adj_5687));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_2162 (.I0(\data_in_frame[17] [1]), .I1(n58290), 
            .I2(n43398), .I3(rx_data[1]), .O(n56474));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2162.LUT_INIT = 16'ha3a0;
    SB_LUT4 i50879_4_lut (.I0(n11_adj_5702), .I1(n9_adj_5682), .I2(n7), 
            .I3(n5), .O(n66607));
    defparam i50879_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13_4_lut_adj_2163 (.I0(\data_in_frame[17] [0]), .I1(n58290), 
            .I2(n43398), .I3(rx_data[0]), .O(n56478));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2163.LUT_INIT = 16'ha3a0;
    SB_LUT4 mux_1584_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n12185));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i50824_4_lut (.I0(n17_adj_5686), .I1(n15_adj_5698), .I2(n13_adj_5703), 
            .I3(n66607), .O(n66552));
    defparam i50824_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_30__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52660_4_lut (.I0(n16_adj_5687), .I1(n6_adj_5676), .I2(n19_adj_5685), 
            .I3(n66548), .O(n68388));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52660_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51020_3_lut (.I0(n68068), .I1(n303), .I2(n15_adj_5698), .I3(GND_net), 
            .O(n66748));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_2164 (.I0(n59370), .I1(\data_in_frame[16] [2]), 
            .I2(n106), .I3(rx_data[2]), .O(n56566));   // verilog/coms.v(130[12] 305[6])
    defparam i14_4_lut_adj_2164.LUT_INIT = 16'hc5c0;
    SB_LUT4 i52825_4_lut (.I0(n66748), .I1(n68388), .I2(n19_adj_5685), 
            .I3(n66552), .O(n68553));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52825_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_3_lut_adj_2165 (.I0(rx_data[7]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57410), .I3(GND_net), .O(n57336));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_2165.LUT_INIT = 16'h0202;
    SB_LUT4 i16296_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n57425), .I3(GND_net), .O(n30372));   // verilog/coms.v(130[12] 305[6])
    defparam i16296_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52826_3_lut (.I0(n68553), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n68554));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52826_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_2166 (.I0(reset), .I1(n105), .I2(GND_net), .I3(GND_net), 
            .O(n106));
    defparam i1_2_lut_adj_2166.LUT_INIT = 16'heeee;
    SB_LUT4 i52743_3_lut (.I0(n68554), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n68471));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52743_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i14_4_lut_adj_2167 (.I0(n59370), .I1(\data_in_frame[16] [0]), 
            .I2(n106), .I3(rx_data[0]), .O(n56568));   // verilog/coms.v(130[12] 305[6])
    defparam i14_4_lut_adj_2167.LUT_INIT = 16'hc5c0;
    SB_LUT4 i46861_3_lut (.I0(duty[22]), .I1(duty[17]), .I2(n294), .I3(GND_net), 
            .O(n62578));
    defparam i46861_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 LessThan_17_i26_3_lut (.I0(n68471), .I1(n298), .I2(duty[12]), 
            .I3(GND_net), .O(n26_adj_5684));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_30__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16363_3_lut_4_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30439));   // verilog/coms.v(130[12] 305[6])
    defparam i16363_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i46865_3_lut (.I0(duty[13]), .I1(duty[21]), .I2(n294), .I3(GND_net), 
            .O(n62582));
    defparam i46865_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i47075_4_lut (.I0(duty[15]), .I1(n62578), .I2(duty[20]), .I3(n294), 
            .O(n62794));
    defparam i47075_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i46857_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n294), .I3(GND_net), 
            .O(n62574));
    defparam i46857_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i10_4_lut (.I0(n294), .I1(n62794), .I2(n62582), .I3(n26_adj_5684), 
            .O(n22_adj_5911));
    defparam i10_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i47073_4_lut (.I0(duty[19]), .I1(n62574), .I2(duty[16]), .I3(n294), 
            .O(n62792));
    defparam i47073_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i16355_3_lut_4_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30431));   // verilog/coms.v(130[12] 305[6])
    defparam i16355_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i51596_3_lut (.I0(n15_adj_5734), .I1(n13_adj_5735), .I2(n11_adj_5736), 
            .I3(GND_net), .O(n67324));
    defparam i51596_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i51536_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n67324), .O(n67264));
    defparam i51536_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i50674_4_lut (.I0(n21_adj_5728), .I1(n19_adj_5729), .I2(n17_adj_5732), 
            .I3(n9_adj_5738), .O(n66402));
    defparam i50674_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51646_4_lut (.I0(n9_adj_5738), .I1(n7_adj_5740), .I2(current[2]), 
            .I3(duty[2]), .O(n67374));
    defparam i51646_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i16353_3_lut_4_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30429));   // verilog/coms.v(130[12] 305[6])
    defparam i16353_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16352_3_lut_4_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30428));   // verilog/coms.v(130[12] 305[6])
    defparam i16352_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_243_i12_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i52046_4_lut (.I0(n15_adj_5734), .I1(n13_adj_5735), .I2(n11_adj_5736), 
            .I3(n67374), .O(n67774));
    defparam i52046_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52038_4_lut (.I0(n21_adj_5728), .I1(n19_adj_5729), .I2(n17_adj_5732), 
            .I3(n67774), .O(n67766));
    defparam i52038_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mux_243_i13_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i14_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i15_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i16_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i52585_4_lut (.I0(current[15]), .I1(n23_adj_5727), .I2(duty[12]), 
            .I3(n67766), .O(n68313));
    defparam i52585_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i51552_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n68313), .O(n67280));
    defparam i51552_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5742));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i21_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(n19_adj_5820), 
            .I3(encoder0_position_scaled[16]), .O(n20_adj_5821));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i6575_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6575_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_30__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6573_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6573_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 mux_243_i18_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i52333_3_lut (.I0(n4_adj_5742), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n68061));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52333_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51482_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5734), .O(n67210));
    defparam i51482_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5726));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i50606_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n67264), .O(n66334));
    defparam i50606_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 encoder0_position_30__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i35_rep_151_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n69974));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_151_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52656_3_lut (.I0(n30_adj_5726), .I1(n10_adj_5737), .I2(n67210), 
            .I3(GND_net), .O(n68384));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51044_4_lut (.I0(n68061), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n66772));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51044_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i52331_3_lut (.I0(n6_adj_5741), .I1(duty[10]), .I2(n21_adj_5728), 
            .I3(GND_net), .O(n68059));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2168 (.I0(n2421), .I1(n2425), .I2(n2428), .I3(n2423), 
            .O(n61852));
    defparam i1_4_lut_adj_2168.LUT_INIT = 16'hfffe;
    SB_LUT4 i52332_3_lut (.I0(n68059), .I1(duty[11]), .I2(n23_adj_5727), 
            .I3(GND_net), .O(n68060));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52030_4_lut (.I0(current[15]), .I1(n23_adj_5727), .I2(duty[12]), 
            .I3(n66402), .O(n67758));
    defparam i52030_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5739), .I1(duty[9]), .I2(n19_adj_5729), 
            .I3(GND_net), .O(n16_adj_5733));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51046_3_lut (.I0(n68060), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n66774));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51046_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52353_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n67280), .O(n68081));
    defparam i52353_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 mux_243_i19_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52793_4_lut (.I0(n66772), .I1(n68384), .I2(n69974), .I3(n66334), 
            .O(n68521));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52793_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_243_i20_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i52130_3_lut (.I0(n66774), .I1(n16_adj_5733), .I2(n67758), 
            .I3(GND_net), .O(n67858));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52864_4_lut (.I0(n67858), .I1(n68521), .I2(n69974), .I3(n68081), 
            .O(n68592));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52864_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29636_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n43611));
    defparam i29636_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i52865_3_lut (.I0(n68592), .I1(duty[18]), .I2(current[15]), 
            .I3(GND_net), .O(n68593));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52865_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_243_i21_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i22_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i52439_4_lut (.I0(n68593), .I1(duty[20]), .I2(current[15]), 
            .I3(duty[19]), .O(n68167));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52439_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i2_4_lut (.I0(n21_adj_5853), .I1(n68167), .I2(duty[21]), .I3(current[15]), 
            .O(n6_adj_5923));
    defparam i2_4_lut.LUT_INIT = 16'heafe;
    SB_LUT4 i7_4_lut_adj_2169 (.I0(duty[22]), .I1(duty[23]), .I2(n6_adj_5923), 
            .I3(current[15]), .O(n11579));
    defparam i7_4_lut_adj_2169.LUT_INIT = 16'h3332;
    SB_LUT4 mux_243_i23_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i24_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i1_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i2_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i27766_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(n41755), 
            .I3(encoder0_position_scaled[6]), .O(n41756));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i27766_3_lut_4_lut.LUT_INIT = 16'he0f1;
    SB_LUT4 mux_243_i6_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i9_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i10_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_2170 (.I0(n61852), .I1(n2427), .I2(n2426), .I3(n2424), 
            .O(n61854));
    defparam i1_4_lut_adj_2170.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i8_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i3_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i11_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i28324_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(n42304), 
            .I3(encoder0_position_scaled[3]), .O(n42305));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i28324_3_lut_4_lut.LUT_INIT = 16'he0f1;
    SB_LUT4 mux_243_i5_3_lut_4_lut (.I0(n25465), .I1(control_mode[1]), .I2(motor_state_23__N_91[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_2171 (.I0(n2429), .I1(n43611), .I2(n2430), .I3(n2431), 
            .O(n59115));
    defparam i1_4_lut_adj_2171.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i26_3_lut (.I0(encoder0_position[25]), .I1(n7_adj_5722), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2172 (.I0(n2417), .I1(n59115), .I2(n61854), .I3(n2420), 
            .O(n61860));
    defparam i1_4_lut_adj_2172.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_2173 (.I0(\data_in_frame[22] [2]), .I1(n58294), 
            .I2(n43396), .I3(rx_data[2]), .O(n56414));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2173.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_4_lut_adj_2174 (.I0(n4_adj_5730), .I1(n5_adj_5725), .I2(n518), 
            .I3(n6_adj_5723), .O(n5_adj_5895));
    defparam i1_4_lut_adj_2174.LUT_INIT = 16'heeea;
    \quadrature_decoder(1)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1779(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .\a_new[1] (a_new_adj_5965[1]), 
            .n29731(n29731), .n1784(n1784), .position_31__N_3827(position_31__N_3827_adj_5754), 
            .n1824(n1824), .n1786(n1786), .n1788(n1788), .n1790(n1790), 
            .n1792(n1792), .n1794(n1794), .n1796(n1796), .\encoder1_position[25] (encoder1_position[25]), 
            .\encoder1_position[24] (encoder1_position[24]), .\encoder1_position[23] (encoder1_position[23]), 
            .\encoder1_position[22] (encoder1_position[22]), .\encoder1_position[21] (encoder1_position[21]), 
            .\encoder1_position[20] (encoder1_position[20]), .\encoder1_position[19] (encoder1_position[19]), 
            .\encoder1_position[18] (encoder1_position[18]), .\encoder1_position[17] (encoder1_position[17]), 
            .\encoder1_position[16] (encoder1_position[16]), .\encoder1_position[15] (encoder1_position[15]), 
            .\encoder1_position[14] (encoder1_position[14]), .\encoder1_position[13] (encoder1_position[13]), 
            .\encoder1_position[12] (encoder1_position[12]), .\encoder1_position[11] (encoder1_position[11]), 
            .\encoder1_position[10] (encoder1_position[10]), .\encoder1_position[9] (encoder1_position[9]), 
            .\encoder1_position[8] (encoder1_position[8]), .\encoder1_position[7] (encoder1_position[7]), 
            .\encoder1_position[6] (encoder1_position[6]), .\encoder1_position[5] (encoder1_position[5]), 
            .\encoder1_position[4] (encoder1_position[4]), .\encoder1_position[3] (encoder1_position[3]), 
            .\encoder1_position[2] (encoder1_position[2]), .n1822(n1822), 
            .GND_net(GND_net), .VCC_net(VCC_net), .b_prev(b_prev_adj_5753)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[49] 318[6])
    SB_LUT4 i1_3_lut_adj_2175 (.I0(n2418), .I1(n2419), .I2(n2422), .I3(GND_net), 
            .O(n61902));
    defparam i1_3_lut_adj_2175.LUT_INIT = 16'hfefe;
    SB_LUT4 i35544_3_lut_4_lut (.I0(n36852), .I1(Ki[3]), .I2(n4_adj_5700), 
            .I3(n20252), .O(n6_adj_5699));
    defparam i35544_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut (.I0(n36852), .I1(Ki[3]), .I2(n4_adj_5700), 
            .I3(n20252), .O(n20203));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i35490_3_lut_4_lut (.I0(n36823), .I1(Ki[2]), .I2(n49420), 
            .I3(n20283), .O(n4_adj_5851));
    defparam i35490_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_2176 (.I0(n36823), .I1(Ki[2]), .I2(n49420), 
            .I3(n20283), .O(n20252));
    defparam i1_3_lut_4_lut_adj_2176.LUT_INIT = 16'h8778;
    SB_LUT4 i13_4_lut_adj_2177 (.I0(\data_in_frame[22] [1]), .I1(n58294), 
            .I2(n43396), .I3(rx_data[1]), .O(n56418));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2177.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_3_lut_adj_2178 (.I0(n3), .I1(n2_adj_5731), .I2(n5_adj_5895), 
            .I3(GND_net), .O(n58170));
    defparam i1_3_lut_adj_2178.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_2179 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5901));
    defparam i1_2_lut_adj_2179.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_2180 (.I0(delay_counter[9]), .I1(n4_adj_5901), 
            .I2(delay_counter[10]), .I3(n25505), .O(n60225));
    defparam i2_4_lut_adj_2180.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_2181 (.I0(n60225), .I1(n25477), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n60151));
    defparam i2_4_lut_adj_2181.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5914));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_2182 (.I0(delay_counter[22]), .I1(n60151), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5915));
    defparam i2_4_lut_adj_2182.LUT_INIT = 16'ha8a0;
    SB_LUT4 i28945_4_lut (.I0(n7_adj_5915), .I1(delay_counter[31]), .I2(n25480), 
            .I3(n8_adj_5914), .O(n1319));   // verilog/TinyFPGA_B.v(379[14:38])
    defparam i28945_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_4_lut_adj_2183 (.I0(n61902), .I1(n2415), .I2(n61860), .I3(n2416), 
            .O(n61864));
    defparam i1_4_lut_adj_2183.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5900));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i42502_3_lut (.I0(n7_adj_5722), .I1(n7455), .I2(n58170), .I3(GND_net), 
            .O(n58179));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_5900), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n25480));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_2184 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25477));
    defparam i2_3_lut_adj_2184.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5908));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_2185 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5907));
    defparam i6_4_lut_adj_2185.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5907), .I1(delay_counter[2]), .I2(n14_adj_5908), 
            .I3(delay_counter[6]), .O(n25505));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4891_4_lut (.I0(n25505), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5824));
    defparam i4891_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_2186 (.I0(n24_adj_5824), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n60298));
    defparam i2_4_lut_adj_2186.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_2187 (.I0(n60298), .I1(delay_counter[18]), .I2(n25477), 
            .I3(GND_net), .O(n60224));
    defparam i2_3_lut_adj_2187.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_2188 (.I0(delay_counter[23]), .I1(n60224), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5744));
    defparam i2_4_lut_adj_2188.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_2189 (.I0(n7_adj_5744), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n25480), .O(n62));
    defparam i4_4_lut_adj_2189.LUT_INIT = 16'hfffe;
    SB_LUT4 i28942_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(365[12:35])
    defparam i28942_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 LessThan_1083_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5834));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i42503_3_lut (.I0(encoder0_position[25]), .I1(n58179), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50755_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n66483));   // verilog/uart_rx.v(119[17:57])
    defparam i50755_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i6_4_lut_adj_2190 (.I0(ID[4]), .I1(ID[7]), .I2(ID[6]), .I3(ID[5]), 
            .O(n14_adj_5909));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i6_4_lut_adj_2190.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_2191 (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5910));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i5_4_lut_adj_2191.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28757_4_lut (.I0(n13_adj_5910), .I1(baudrate[0]), .I2(n14_adj_5909), 
            .I3(n25593), .O(n42725));
    defparam i28757_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 i14839_4_lut (.I0(n27728), .I1(n1319), .I2(n65611), .I3(n42845), 
            .O(n28915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i14839_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 mux_4310_i9_3_lut (.I0(encoder0_position[8]), .I1(n24_adj_5707), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut_adj_2192 (.I0(n36852), .I1(Ki[2]), .I2(n49470), 
            .I3(n20253), .O(n20204));
    defparam i1_3_lut_4_lut_adj_2192.LUT_INIT = 16'h8778;
    SB_LUT4 i35536_3_lut_4_lut (.I0(n36852), .I1(Ki[2]), .I2(n49470), 
            .I3(n20253), .O(n4_adj_5700));
    defparam i35536_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i15556_3_lut_4_lut (.I0(reset), .I1(n28413), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29632));
    defparam i15556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21719_3_lut_4_lut (.I0(reset), .I1(n28413), .I2(\data_in_frame[20] [6]), 
            .I3(rx_data[6]), .O(n30176));
    defparam i21719_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i15548_3_lut_4_lut (.I0(reset), .I1(n28413), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29624));
    defparam i15548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15545_3_lut_4_lut (.I0(reset), .I1(n28413), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29621));
    defparam i15545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15542_3_lut_4_lut (.I0(reset), .I1(n28413), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29618));
    defparam i15542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15533_3_lut_4_lut (.I0(reset), .I1(n28413), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29609));
    defparam i15533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35523_2_lut_3_lut_4_lut (.I0(n36823), .I1(Ki[0]), .I2(Ki[1]), 
            .I3(n36852), .O(n20205));
    defparam i35523_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i35525_2_lut_3_lut_4_lut (.I0(n36823), .I1(Ki[0]), .I2(Ki[1]), 
            .I3(n36852), .O(n49470));
    defparam i35525_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 encoder0_position_30__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_2193 (.I0(n15_adj_5743), .I1(n22917), .I2(dti), 
            .I3(GND_net), .O(n27652));
    defparam i1_2_lut_3_lut_adj_2193.LUT_INIT = 16'hbaba;
    SB_LUT4 encoder0_position_30__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53281_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n61864), 
            .O(n2445));
    defparam i53281_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50742_3_lut_4_lut (.I0(r_Clock_Count_adj_5997[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5997[2]), .O(n66470));   // verilog/uart_tx.v(117[17:57])
    defparam i50742_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_30__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229_adj_5807));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i840_3_lut (.I0(n1229_adj_5807), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1086_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5997[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5838));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 encoder0_position_30__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(1)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1779(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .\a_new[1] (a_new[1]), 
            .b_prev(b_prev), .n29751(n29751), .n1742(n1742), .position_31__N_3827(position_31__N_3827), 
            .n1744(n1744), .\encoder0_position[30] (encoder0_position[30]), 
            .\encoder0_position[29] (encoder0_position[29]), .\encoder0_position[28] (encoder0_position[28]), 
            .\encoder0_position[27] (encoder0_position[27]), .\encoder0_position[26] (encoder0_position[26]), 
            .\encoder0_position[25] (encoder0_position[25]), .\encoder0_position[24] (encoder0_position[24]), 
            .\encoder0_position[23] (encoder0_position[23]), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(304[49] 310[6])
    SB_LUT4 i13_3_lut_4_lut (.I0(rx_data[4]), .I1(n41114), .I2(n43396), 
            .I3(\data_in_frame[22] [4]), .O(n56406));   // verilog/coms.v(130[12] 305[6])
    defparam i13_3_lut_4_lut.LUT_INIT = 16'hf202;
    SB_LUT4 i13_3_lut_4_lut_adj_2194 (.I0(rx_data[4]), .I1(n41114), .I2(n43398), 
            .I3(\data_in_frame[17] [4]), .O(n56462));   // verilog/coms.v(130[12] 305[6])
    defparam i13_3_lut_4_lut_adj_2194.LUT_INIT = 16'hf202;
    SB_LUT4 encoder0_position_30__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    TLI4970 tli (.\state[1] (state_adj_5987[1]), .clk16MHz(clk16MHz), .clk_out(clk_out), 
            .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), .GND_net(GND_net), .n15(n15_adj_5750), 
            .\state[0] (state_adj_5987[0]), .n11(n11_adj_5751), .n29691(n29691), 
            .\data[15] (data_adj_5985[15]), .n9(n9_adj_5916), .n29677(n29677), 
            .n29675(n29675), .\current[0] (current[0]), .n29672(n29672), 
            .\data[12] (data_adj_5985[12]), .n29671(n29671), .\data[11] (data_adj_5985[11]), 
            .n29656(n29656), .\data[10] (data_adj_5985[10]), .n29655(n29655), 
            .\data[9] (data_adj_5985[9]), .n29654(n29654), .\data[8] (data_adj_5985[8]), 
            .n29653(n29653), .\data[7] (data_adj_5985[7]), .n29652(n29652), 
            .\data[6] (data_adj_5985[6]), .n29645(n29645), .\data[5] (data_adj_5985[5]), 
            .n29637(n29637), .\data[4] (data_adj_5985[4]), .n29636(n29636), 
            .\data[3] (data_adj_5985[3]), .n29635(n29635), .\data[2] (data_adj_5985[2]), 
            .n29628(n29628), .\data[1] (data_adj_5985[1]), .VCC_net(VCC_net), 
            .n30538(n30538), .\data[0] (data_adj_5985[0]), .n30427(n30427), 
            .\current[1] (current[1]), .n30426(n30426), .\current[2] (current[2]), 
            .n30425(n30425), .\current[3] (current[3]), .n30424(n30424), 
            .\current[4] (current[4]), .n30423(n30423), .\current[5] (current[5]), 
            .n30422(n30422), .\current[6] (current[6]), .n30421(n30421), 
            .\current[7] (current[7]), .n30420(n30420), .\current[8] (current[8]), 
            .n30419(n30419), .\current[9] (current[9]), .n30418(n30418), 
            .\current[10] (current[10]), .n30417(n30417), .\current[11] (current[11]), 
            .n6(n6_adj_5749), .n27736(n27736), .\current[15] (current[15]), 
            .n5(n5_adj_5798), .n6_adj_31(n6_adj_5748), .state_7__N_4317(state_7__N_4317), 
            .n42880(n42880), .n25615(n25615), .n25587(n25587), .n25590(n25590), 
            .n25578(n25578), .n25583(n25583), .n6_adj_32(n6), .n5_adj_33(n5_adj_5724)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(404[11] 410[4])
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i15667_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [1]), 
            .I3(current_limit[9]), .O(n29743));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15666_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [2]), 
            .I3(current_limit[10]), .O(n29742));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15659_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [3]), 
            .I3(current_limit[11]), .O(n29735));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15658_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [4]), 
            .I3(current_limit[12]), .O(n29734));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15668_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [0]), 
            .I3(current_limit[8]), .O(n29744));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16295_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [1]), 
            .I3(current_limit[1]), .O(n30371));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16295_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i21724_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [6]), 
            .I3(current_limit[14]), .O(n29732));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i21724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15681_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n29757));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15681_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15682_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n29758));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16305_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n30381));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16305_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16240_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [4]), 
            .I3(current_limit[4]), .O(n30316));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16240_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21728_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [7]), 
            .I3(current_limit[15]), .O(n29692));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i21728_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15587_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n29663));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15587_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i21729_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[20] [5]), 
            .I3(current_limit[13]), .O(n29733));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i21729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16241_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [3]), 
            .I3(current_limit[3]), .O(n30317));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16241_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16339_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n30415));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16339_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16211_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [5]), 
            .I3(current_limit[5]), .O(n30287));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16211_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16425_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n30501));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_4310_i23_3_lut (.I0(encoder0_position[22]), .I1(n10), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15680_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n29756));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15680_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15683_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [7]), 
            .I3(current_limit[7]), .O(n29759));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15683_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i709_3_lut (.I0(n521), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16260_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [2]), 
            .I3(current_limit[2]), .O(n30336));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16260_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15588_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [0]), 
            .I3(current_limit[0]), .O(n29664));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15588_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16189_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[21] [6]), 
            .I3(current_limit[6]), .O(n30265));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16189_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15679_3_lut_4_lut (.I0(n2873), .I1(n27726), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n29755));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15679_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232_adj_5810));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i843_3_lut (.I0(n1232_adj_5810), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1178_3_lut (.I0(n1727), .I1(n1794_adj_5816), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15803_3_lut_4_lut (.I0(deadband[2]), .I1(\data_in_frame[16] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29879));   // verilog/coms.v(130[12] 305[6])
    defparam i15803_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    coms neopxl_color_23__I_0 (.n56422(n56422), .\data_in_frame[22] ({\data_in_frame[22] }), 
         .clk16MHz(clk16MHz), .VCC_net(VCC_net), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .GND_net(GND_net), .n2873(n2873), .rx_data({rx_data}), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_in_frame[3] ({Open_3, Open_4, \data_in_frame[3] [5], Open_5, 
         Open_6, Open_7, Open_8, Open_9}), .n7(n7_adj_5921), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n29989(n29989), .n29986(n29986), .n29983(n29983), .n56418(n56418), 
         .n29979(n29979), .n29976(n29976), .n56414(n56414), .\data_in_frame[3][6] (\data_in_frame[3] [6]), 
         .\data_in_frame[3][4] (\data_in_frame[3] [4]), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .\data_in_frame[3][2] (\data_in_frame[3] [2]), .n29701(n29701), 
         .\data_in_frame[0][1] (\data_in_frame[0] [1]), .\data_in_frame[3][1] (\data_in_frame[3] [1]), 
         .\data_in_frame[3][0] (\data_in_frame[3] [0]), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .n56410(n56410), .\data_in_frame[10] ({Open_10, \data_in_frame[10] [6], 
         Open_11, \data_in_frame[10] [4], Open_12, Open_13, Open_14, 
         Open_15}), .n58117(n58117), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[0][7] (\data_in_frame[0] [7]), .Kp_23__N_1748(Kp_23__N_1748), 
         .reset(reset), .n56406(n56406), .setpoint({setpoint}), .n56402(n56402), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .n57657(n57657), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .\byte_transmit_counter[2] (byte_transmit_counter[2]), .\byte_transmit_counter[1] (byte_transmit_counter[1]), 
         .\data_in_frame[14] ({\data_in_frame[14] }), .n6(n6_adj_5704), 
         .n69640(n69640), .n43(n43_adj_5831), .n379(n379), .n405(n405), 
         .n4(n4_adj_5826), .pwm_setpoint({pwm_setpoint}), .n29714(n29714), 
         .encoder0_position_scaled({encoder0_position_scaled}), .n459(n459), 
         .n11610(n11610), .n37308(n37308), .n57425(n57425), .n56398(n56398), 
         .\FRAME_MATCHER.i[4] (\FRAME_MATCHER.i [4]), .\FRAME_MATCHER.i[5] (\FRAME_MATCHER.i [5]), 
         .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), .DE_c(DE_c), .n29739(n29739), 
         .\data_in_frame[0][2] (\data_in_frame[0] [2]), .LED_c(LED_c), .n33801(n33801), 
         .\FRAME_MATCHER.i_31__N_2513 (\FRAME_MATCHER.i_31__N_2513 ), .n27726(n27726), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .n29764(n29764), .\data_in_frame[0][3] (\data_in_frame[0] [3]), 
         .\data_out_frame[20] ({\data_out_frame[20] [7:6], Open_16, Open_17, 
         Open_18, Open_19, Open_20, Open_21}), .n29802(n29802), .deadband({deadband}), 
         .n29879(n29879), .n29878(n29878), .n29877(n29877), .n29876(n29876), 
         .n29875(n29875), .n29874(n29874), .n29873(n29873), .n29872(n29872), 
         .n29871(n29871), .n29870(n29870), .n29869(n29869), .n29868(n29868), 
         .n29867(n29867), .n29866(n29866), .n29865(n29865), .n29864(n29864), 
         .n29863(n29863), .n29862(n29862), .n29861(n29861), .n29860(n29860), 
         .n29859(n29859), .n29858(n29858), .n29857(n29857), .IntegralLimit({IntegralLimit}), 
         .n29856(n29856), .n29855(n29855), .n29854(n29854), .n29853(n29853), 
         .n53095(n53095), .n52011(n52011), .n29852(n29852), .n29851(n29851), 
         .n57836(n57836), .\data_out_frame[18][3] (\data_out_frame[18] [3]), 
         .n3470(n3470), .rx_data_ready(rx_data_ready), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .\data_out_frame[23][3] (\data_out_frame[23] [3]), .\data_out_frame[16][3] (\data_out_frame[16] [3]), 
         .n29850(n29850), .n29849(n29849), .n29848(n29848), .n29847(n29847), 
         .\data_out_frame[25][2] (\data_out_frame[25] [2]), .n29846(n29846), 
         .n29845(n29845), .n29844(n29844), .n29843(n29843), .\data_in_frame[0][0] (\data_in_frame[0] [0]), 
         .n29842(n29842), .n29841(n29841), .n29840(n29840), .n29839(n29839), 
         .n29838(n29838), .n29837(n29837), .n29836(n29836), .n29835(n29835), 
         .n29834(n29834), .\Kp[1] (Kp[1]), .\data_out_frame[24][2] (\data_out_frame[24] [2]), 
         .n29833(n29833), .\Kp[2] (Kp[2]), .n29832(n29832), .\Kp[3] (Kp[3]), 
         .n29831(n29831), .\Kp[4] (Kp[4]), .n29830(n29830), .\Kp[5] (Kp[5]), 
         .n29829(n29829), .\Kp[6] (Kp[6]), .n57437(n57437), .\Kp[7] (Kp[7]), 
         .n29827(n29827), .\Kp[8] (Kp[8]), .n29826(n29826), .\Kp[9] (Kp[9]), 
         .n29825(n29825), .\Kp[10] (Kp[10]), .n29824(n29824), .\Kp[11] (Kp[11]), 
         .n172(n172), .\data_out_frame[20][3] (\data_out_frame[20] [3]), 
         .n29823(n29823), .\Kp[12] (Kp[12]), .n29822(n29822), .\Kp[13] (Kp[13]), 
         .n28413(n28413), .n29821(n29821), .\Kp[14] (Kp[14]), .n29820(n29820), 
         .\Kp[15] (Kp[15]), .n29819(n29819), .\Ki[1] (Ki[1]), .n29818(n29818), 
         .\Ki[2] (Ki[2]), .n29817(n29817), .\Ki[3] (Ki[3]), .n29816(n29816), 
         .\Ki[4] (Ki[4]), .n29815(n29815), .\Ki[5] (Ki[5]), .n29814(n29814), 
         .\Ki[6] (Ki[6]), .n29813(n29813), .\Ki[7] (Ki[7]), .n29812(n29812), 
         .\Ki[8] (Ki[8]), .n29811(n29811), .\Ki[9] (Ki[9]), .n29810(n29810), 
         .\Ki[10] (Ki[10]), .n29809(n29809), .\Ki[11] (Ki[11]), .n29808(n29808), 
         .\Ki[12] (Ki[12]), .n29807(n29807), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
         .n29805(n29805), .\Ki[15] (Ki[15]), .\data_in_frame[16] ({\data_in_frame[16] }), 
         .n105(n105), .\data_out_frame[18][4] (\data_out_frame[18] [4]), 
         .\data_out_frame[17][3] (\data_out_frame[17] [3]), .n25848(n25848), 
         .n29767(n29767), .n26517(n26517), .n29760(n29760), .neopxl_color({neopxl_color}), 
         .n29759(n29759), .current_limit({current_limit}), .n29758(n29758), 
         .control_mode({control_mode}), .n29757(n29757), .n29756(n29756), 
         .n29755(n29755), .n29754(n29754), .n29753(n29753), .n29752(n29752), 
         .n29750(n29750), .n29749(n29749), .n29748(n29748), .n29747(n29747), 
         .n29746(n29746), .n29745(n29745), .n29744(n29744), .n29743(n29743), 
         .n29742(n29742), .n161(n161), .n31(n31_adj_5822), .\data_out_frame[19][3] (\data_out_frame[19] [3]), 
         .n29738(n29738), .n7_adj_10(n7_adj_5917), .n29735(n29735), .encoder1_position_scaled({encoder1_position_scaled}), 
         .n29734(n29734), .n29733(n29733), .n29732(n29732), .n25(n25_adj_5812), 
         .n29730(n29730), .n29729(n29729), .n29725(n29725), .n29721(n29721), 
         .n29718(n29718), .\data_out_frame[22][3] (\data_out_frame[22] [3]), 
         .n57879(n57879), .n59684(n59684), .n57499(n57499), .n29700(n29700), 
         .n29699(n29699), .n29692(n29692), .n29673(n29673), .PWMLimit({PWMLimit}), 
         .n29664(n29664), .n29663(n29663), .n29662(n29662), .n29661(n29661), 
         .\Ki[0] (Ki[0]), .n29660(n29660), .\Kp[0] (Kp[0]), .n29644(n29644), 
         .\data_in_frame[18] ({\data_in_frame[18] }), .\pwm_counter[22] (pwm_counter[22]), 
         .n45(n45), .\pwm_counter[21] (pwm_counter[21]), .n43_adj_11(n43), 
         .\data_out_frame[21][0] (\data_out_frame[21] [0]), .\data_out_frame[21][3] (\data_out_frame[21] [3]), 
         .\data_in_frame[19] ({Open_22, \data_in_frame[19] [6:0]}), .n53127(n53127), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .\current[7] (current[7]), 
         .\current[6] (current[6]), .n29471(n29471), .n30549(n30549), 
         .n30548(n30548), .n30547(n30547), .n30546(n30546), .n30545(n30545), 
         .n30544(n30544), .n30543(n30543), .n29474(n29474), .n30534(n30534), 
         .n29477(n29477), .n30512(n30512), .n30506(n30506), .n30504(n30504), 
         .n30503(n30503), .n30501(n30501), .n30500(n30500), .n30499(n30499), 
         .n30498(n30498), .n30490(n30490), .n30439(n30439), .n30431(n30431), 
         .n30429(n30429), .n30428(n30428), .n30415(n30415), .tx_active(tx_active), 
         .n30383(n30383), .n30382(n30382), .n30381(n30381), .n30380(n30380), 
         .n30378(n30378), .n56568(n56568), .n30372(n30372), .n30371(n30371), 
         .n56566(n56566), .n29520(n29520), .n29523(n29523), .n29526(n29526), 
         .n29530(n29530), .n56478(n56478), .n56474(n56474), .n56470(n56470), 
         .n56466(n56466), .n56462(n56462), .n56458(n56458), .n30343(n30343), 
         .n56454(n56454), .n56450(n56450), .n56446(n56446), .\data_in_frame[6] ({Open_23, 
         Open_24, \data_in_frame[6] [5:0]}), .n30336(n30336), .n30055(n30055), 
         .\data_in_frame[7][1] (\data_in_frame[7] [1]), .n30059(n30059), 
         .\data_in_frame[7][2] (\data_in_frame[7] [2]), .n30062(n30062), 
         .\data_in_frame[7][3] (\data_in_frame[7] [3]), .n30065(n30065), 
         .\data_in_frame[7][4] (\data_in_frame[7] [4]), .n30068(n30068), 
         .\data_in_frame[7][5] (\data_in_frame[7] [5]), .n30077(n30077), 
         .n30080(n30080), .n30083(n30083), .n30317(n30317), .n30316(n30316), 
         .n30087(n30087), .n30314(n30314), .n30093(n30093), .n30096(n30096), 
         .n30099(n30099), .n30102(n30102), .n30105(n30105), .n30108(n30108), 
         .n30112(n30112), .n30115(n30115), .n30118(n30118), .n30122(n30122), 
         .n30125(n30125), .n30131(n30131), .\data_in_frame[10][1] (\data_in_frame[10] [1]), 
         .n30134(n30134), .\data_in_frame[10][2] (\data_in_frame[10] [2]), 
         .n30138(n30138), .\data_in_frame[10][3] (\data_in_frame[10] [3]), 
         .n30141(n30141), .n30144(n30144), .\data_in_frame[10][5] (\data_in_frame[10] [5]), 
         .n30148(n30148), .n30151(n30151), .\data_in_frame[10][7] (\data_in_frame[10] [7]), 
         .n30154(n30154), .\data_in_frame[11] ({\data_in_frame[11] }), .n56662(n56662), 
         .n56678(n56678), .n56604(n56604), .n30167(n30167), .n30170(n30170), 
         .n30173(n30173), .n30287(n30287), .n30177(n30177), .n30180(n30180), 
         .n30183(n30183), .n30186(n30186), .n56636(n56636), .n56690(n56690), 
         .n30196(n30196), .n30199(n30199), .n30203(n30203), .n56442(n56442), 
         .n56438(n56438), .\current[5] (current[5]), .n30265(n30265), 
         .n29570(n29570), .n29573(n29573), .n29576(n29576), .n56434(n56434), 
         .n56430(n56430), .n56546(n56546), .n56542(n56542), .\current[4] (current[4]), 
         .\current[3] (current[3]), .n56540(n56540), .n29594(n29594), 
         .n56538(n56538), .n56536(n56536), .n56534(n56534), .n29609(n29609), 
         .\data_in_frame[20] ({\data_in_frame[20] }), .n29618(n29618), .n29621(n29621), 
         .\current[2] (current[2]), .\current[1] (current[1]), .n29624(n29624), 
         .\current[0] (current[0]), .n30176(n30176), .\current[15] (current[15]), 
         .n29632(n29632), .n8(n8_adj_5801), .\current[11] (current[11]), 
         .\current[10] (current[10]), .\current[9] (current[9]), .\current[8] (current[8]), 
         .displacement({displacement}), .n8_adj_12(n8_adj_5774), .n57426(n57426), 
         .n29536(n29536), .n57956(n57956), .n8_adj_13(n8_adj_5757), .n57424(n57424), 
         .n380(n380), .n460(n460), .n27722(n27722), .n29510(n29510), 
         .n33(n33), .n38(n38_adj_5847), .n34(n34), .n57990(n57990), 
         .n57737(n57737), .n33793(n33793), .n29508(n29508), .n52054(n52054), 
         .n58132(n58132), .n53024(n53024), .n57862(n57862), .n52186(n52186), 
         .n57625(n57625), .n57410(n57410), .n28409(n28409), .n53215(n53215), 
         .\data_out_frame[26][2] (\data_out_frame[26] [2]), .\data_out_frame[27][2] (\data_out_frame[27] [2]), 
         .n29999(n29999), .n22792(n22792), .n35(n35), .n4_adj_14(n4_adj_5827), 
         .Kp_23__N_1389(Kp_23__N_1389), .n57685(n57685), .n8_adj_15(n8_adj_5776), 
         .n4_adj_16(n4_adj_5830), .ID({ID}), .n15(n15_adj_5701), .n15_adj_17(n15), 
         .n19(n19_adj_5820), .n28464(n28464), .n91(n91), .n58278(n58278), 
         .n7_adj_18(n7_adj_5920), .n26(n26), .n21(n21_adj_5853), .n260(n260), 
         .n41114(n41114), .n59370(n59370), .n69808(n69808), .n63007(n63007), 
         .n63008(n63008), .n63155(n63155), .n63154(n63154), .n30(n30_adj_5828), 
         .n365(n365), .n32(n32_adj_5829), .n65564(n65564), .tx_o(tx_o), 
         .r_SM_Main({r_SM_Main_adj_5996}), .n29690(n29690), .n58304(n58304), 
         .r_Clock_Count({r_Clock_Count_adj_5997}), .n6_adj_19(n6_adj_5893), 
         .n4940(n4940), .n27(n27_adj_5825), .tx_enable(tx_enable), .baudrate({baudrate}), 
         .\r_SM_Main[2]_adj_20 (r_SM_Main[2]), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
         .n4937(n4937), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), .n61106(n61106), 
         .n29912(n29912), .n61058(n61058), .n57317(n57317), .\r_SM_Main[1]_adj_21 (r_SM_Main[1]), 
         .n27754(n27754), .n61138(n61138), .n29900(n29900), .n25593(n25593), 
         .n29798(n29798), .n29797(n29797), .n29796(n29796), .\r_Bit_Index[0] (r_Bit_Index[0]), 
         .r_Clock_Count_adj_30({r_Clock_Count}), .n27996(n27996), .n58373(n58373), 
         .n30533(n30533), .n53222(n53222), .n30529(n30529), .n30231(n30231), 
         .n30230(n30230), .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), 
         .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), 
         .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), 
         .n61170(n61170), .n61154(n61154), .n61090(n61090), .n61074(n61074), 
         .n61122(n61122)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 encoder0_position_30__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15802_3_lut_4_lut (.I0(deadband[3]), .I1(\data_in_frame[16] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29878));   // verilog/coms.v(130[12] 305[6])
    defparam i15802_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13_4_lut_adj_2195 (.I0(\data_in_frame[22] [0]), .I1(n58294), 
            .I2(n43396), .I3(rx_data[0]), .O(n56422));   // verilog/coms.v(130[12] 305[6])
    defparam i13_4_lut_adj_2195.LUT_INIT = 16'ha3a0;
    SB_LUT4 encoder0_position_30__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_2196 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5904));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_2196.LUT_INIT = 16'hfffe;
    SB_LUT4 i15801_3_lut_4_lut (.I0(deadband[4]), .I1(\data_in_frame[16] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29877));   // verilog/coms.v(130[12] 305[6])
    defparam i15801_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i29680_4_lut (.I0(n519), .I1(n831), .I2(n832), .I3(n833), 
            .O(n43655));
    defparam i29680_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15800_3_lut_4_lut (.I0(deadband[5]), .I1(\data_in_frame[16] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29876));   // verilog/coms.v(130[12] 305[6])
    defparam i15800_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i29790_4_lut (.I0(n829), .I1(n828), .I2(n43655), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i29790_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    motorControl control (.\Ki[10] (Ki[10]), .\PID_CONTROLLER.integral_23__N_3715[0] (\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .GND_net(GND_net), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
            .\Kp[0] (Kp[0]), .\Kp[1] (Kp[1]), .\Ki[14] (Ki[14]), .n365(n365), 
            .control_update(control_update), .duty({duty}), .clk16MHz(clk16MHz), 
            .reset(reset), .IntegralLimit({IntegralLimit}), .n155(n155), 
            .\Kp[5] (Kp[5]), .PWMLimit({PWMLimit}), .\Kp[6] (Kp[6]), .\Kp[9] (Kp[9]), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[7] (Kp[7]), .\Kp[12] (Kp[12]), 
            .\Kp[8] (Kp[8]), .\Kp[13] (Kp[13]), .\Ki[1] (Ki[1]), .\PID_CONTROLLER.integral_23__N_3715[16] (\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .\Ki[15] (Ki[15]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Kp[14] (Kp[14]), 
            .\Ki[4] (Ki[4]), .\Kp[15] (Kp[15]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Kp[3] (Kp[3]), .deadband({deadband}), .n380(n380), 
            .n379(n379), .setpoint({setpoint}), .\motor_state[10] (motor_state[10]), 
            .\motor_state[9] (motor_state[9]), .\motor_state[8] (motor_state[8]), 
            .\motor_state[7] (motor_state[7]), .n41756(n41756), .\PID_CONTROLLER.integral_23__N_3715[23] (\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .\motor_state[5] (motor_state[5]), .\Kp[2] (Kp[2]), .\Kp[4] (Kp[4]), 
            .\motor_state[4] (motor_state[4]), .n42305(n42305), .\motor_state[2] (motor_state[2]), 
            .\PID_CONTROLLER.integral_23__N_3715[22] (\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .\PID_CONTROLLER.integral_23__N_3715[21] (\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .\PID_CONTROLLER.integral_23__N_3715[20] (\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .n212(n212), .n213(n213), .n214(n214), .\motor_state[1] (motor_state[1]), 
            .n4(n4_adj_5826), .n37308(n37308), .n11610(n11610), .\PID_CONTROLLER.integral_23__N_3715[15] (\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .\PID_CONTROLLER.integral_23__N_3715[14] (\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .\Ki[0] (Ki[0]), .\motor_state[0] (motor_state[0]), .VCC_net(VCC_net), 
            .\Ki[8] (Ki[8]), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .\Ki[9] (Ki[9]), .n38(n38), .n29669(n29669), .n110(n110), 
            .n30497(n30497), .n30496(n30496), .n30495(n30495), .n30494(n30494), 
            .n30493(n30493), .n30491(n30491), .n30489(n30489), .n30488(n30488), 
            .n30487(n30487), .n30486(n30486), .n30485(n30485), .n30484(n30484), 
            .n30483(n30483), .n30482(n30482), .n30481(n30481), .n30480(n30480), 
            .n30479(n30479), .n30478(n30478), .n30477(n30477), .n30476(n30476), 
            .n30475(n30475), .n30474(n30474), .n30473(n30473), .\PID_CONTROLLER.integral_23__N_3715[13] (\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .\PID_CONTROLLER.integral_23__N_3715[12] (\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .n27722(n27722), .n53(n53), .n459(n459), .n460(n460), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .n219(n219), .\motor_state[20] (motor_state[20]), .\PID_CONTROLLER.integral_23__N_3715[11] (\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .\motor_state[19] (motor_state[19]), .n490(n490), .n417(n417), 
            .\motor_state[18] (motor_state[18]), .n20203(n20203), .n344(n344), 
            .\motor_state[17] (motor_state[17]), .n20204(n20204), .n271(n271), 
            .n20205(n20205), .n198(n198), .n56(n56), .n125(n125), .n20(n20_adj_5821), 
            .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .n405(n405), .\motor_state[13] (motor_state[13]), .\motor_state[12] (motor_state[12]), 
            .n43(n43_adj_5831), .\motor_state[11] (motor_state[11]), .\PID_CONTROLLER.integral_23__N_3715[10] (\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .n4_adj_7(n4_adj_5827), .n30(n30_adj_5828), .\PID_CONTROLLER.integral_23__N_3715[9] (\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .\PID_CONTROLLER.integral_23__N_3715[8] (\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .\PID_CONTROLLER.integral_23__N_3715[7] (\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .\PID_CONTROLLER.integral_23__N_3715[6] (\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .n6(n6_adj_5699), .n36852(n36852), .n4_adj_8(n4_adj_5851), 
            .n36823(n36823), .\PID_CONTROLLER.integral_23__N_3715[5] (\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .\PID_CONTROLLER.integral_23__N_3715[4] (\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .\PID_CONTROLLER.integral_23__N_3715[3] (\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .\PID_CONTROLLER.integral_23__N_3715[2] (\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .\PID_CONTROLLER.integral_23__N_3715[1] (\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .n43450(n43450), .n20253(n20253), .n49420(n49420), .n20283(n20283), 
            .n35(n35), .n4_adj_9(n4_adj_5830), .n32(n32_adj_5829)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 302[4])
    SB_LUT4 i42498_3_lut (.I0(n5_adj_5725), .I1(n7453), .I2(n58170), .I3(GND_net), 
            .O(n58175));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42498_3_lut.LUT_INIT = 16'hcaca;
    pwm PWM (.n2873(n2873), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .\pwm_counter[21] (pwm_counter[21]), .\pwm_counter[22] (pwm_counter[22]), 
        .pwm_setpoint({pwm_setpoint}), .reset(reset), .n45(n45), .n43(n43), 
        .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    EEPROM eeprom (.enable_slow_N_4211(enable_slow_N_4211), .ready_prev(ready_prev), 
           .clk16MHz(clk16MHz), .n5773({n5774}), .\state[2] (state_adj_5979[2]), 
           .\state[0] (state_adj_6010[0]), .n57392(n57392), .GND_net(GND_net), 
           .n3(n3_adj_5800), .\state[1] (state_adj_5979[1]), .\state[0]_adj_4 (state_adj_5979[0]), 
           .data({data_adj_5978}), .ID({ID}), .n25471(n25471), .n28027(n28027), 
           .n29676(n29676), .rw(rw), .n56774(n56774), .data_ready(data_ready), 
           .n56368(n56368), .n56570(n56570), .baudrate({baudrate}), .n30440(n30440), 
           .n30438(n30438), .n30437(n30437), .n30436(n30436), .n30435(n30435), 
           .n30434(n30434), .n30433(n30433), .n30432(n30432), .n42792(n42792), 
           .n25612(n25612), .\state_7__N_3916[0] (state_7__N_3916[0]), .scl_enable(scl_enable), 
           .VCC_net(VCC_net), .\state_7__N_4108[0] (state_7__N_4108[0]), 
           .\saved_addr[0] (saved_addr[0]), .\state_7__N_4124[3] (state_7__N_4124[3]), 
           .n10(n10_adj_5747), .n6428(n6428), .n10_adj_5(n10_adj_5892), 
           .n29683(n29683), .n30523(n30523), .n8(n8_adj_5918), .n30246(n30246), 
           .n30245(n30245), .n30244(n30244), .n30243(n30243), .n30242(n30242), 
           .n30241(n30241), .n30240(n30240), .scl(scl), .sda_enable(sda_enable), 
           .n65775(n65775), .n25595(n25595), .n25600(n25600), .sda_out(sda_out), 
           .n4(n4_adj_5745), .n4_adj_6(n4_adj_5746), .n42890(n42890)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(390[10] 402[6])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, \neo_pixel_transmitter.t0 , 
            GND_net, state, bit_ctr, timer, neopxl_color, n23, n43567, 
            n27950, n29707, n111, VCC_net, n30355, n30354, n30353, 
            n30352, n30351, n30350, n30349, n30348, n30347, n30342, 
            n30251, n5, NEOPXL_c, n25, LED_c) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output [10:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    output [1:0]state;
    output [4:0]bit_ctr;
    output [10:0]timer;
    input [23:0]neopxl_color;
    output n23;
    output n43567;
    output n27950;
    input n29707;
    output n111;
    input VCC_net;
    input n30355;
    input n30354;
    input n30353;
    input n30352;
    input n30351;
    input n30350;
    input n30349;
    input n30348;
    input n30347;
    input n30342;
    input n30251;
    input n5;
    output NEOPXL_c;
    output n25;
    input LED_c;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n60559, \neo_pixel_transmitter.done , 
        start_N_507, n7, start;
    wire [10:0]n13;
    
    wire n75, n58397, n58415, n41, n48, n112, \neo_pixel_transmitter.done_N_524 , 
        n54, n27707, n65742, n58298, n51632, n29203, n69508, n69496;
    wire [5:0]color_bit_N_502;
    
    wire n63106, n69460, n69814, n67842, n65791, n58165, n67966, 
        n52115;
    wire [1:0]state_1__N_440;
    
    wire n25553, n25554, n1;
    wire [10:0]one_wire_N_479;
    
    wire n49558, n69457, n115, n49557, n69493, n69505, n49556, 
        n49555, n7_adj_5667, n49554, n6_adj_5668, n49553, n8, n49552, 
        n69811, n49551;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(17[11:18])
    
    wire n41_adj_5671, n49550, n6897, n29199;
    wire [10:0]n49;
    
    wire n65744, n63160, n63161, n69625;
    wire [31:0]n137;
    
    wire n43457, n50777, n50776, n50775, n50774, n50773, n50772, 
        n50771, n50770, n50769, n50768, n49549, n4_adj_5674, n58296, 
        n40890, n63149, n63148, n69628, n27940, n28911, n27954, 
        n60566, n59_adj_5675, n33, n62744;
    
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n60559), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i42730_2_lut (.I0(n75), .I1(n58397), .I2(GND_net), .I3(GND_net), 
            .O(n58415));
    defparam i42730_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i71_4_lut (.I0(n41), .I1(n58415), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[1]), .O(n48));
    defparam i71_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut (.I0(n112), .I1(\neo_pixel_transmitter.done_N_524 ), 
            .I2(n75), .I3(state[0]), .O(n54));
    defparam i1_4_lut.LUT_INIT = 16'h5d55;
    SB_LUT4 i1_4_lut_adj_1969 (.I0(state[0]), .I1(n54), .I2(n48), .I3(n58397), 
            .O(n27707));
    defparam i1_4_lut_adj_1969.LUT_INIT = 16'h50dc;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_524 ));   // verilog/neopixel.v(34[12] 116[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(n65742), .I1(n58298), .I2(\neo_pixel_transmitter.done ), 
            .I3(n51632), .O(n29203));   // verilog/neopixel.v(34[12] 116[6])
    defparam i14_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i47378_3_lut (.I0(n69508), .I1(n69496), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n63106));
    defparam i47378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52114_3_lut (.I0(n69460), .I1(n69814), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n67842));
    defparam i52114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28759_4_lut (.I0(n65791), .I1(n58165), .I2(n67966), .I3(n52115), 
            .O(state_1__N_440[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i28759_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 state_1__I_0_102_Mux_0_i1_4_lut (.I0(n25553), .I1(n25554), .I2(state[0]), 
            .I3(bit_ctr[0]), .O(n1));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_102_Mux_0_i1_4_lut.LUT_INIT = 16'hca35;
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n49558), .O(one_wire_N_479[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut_53759_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n69457));   // verilog/neopixel.v(18[6:15])
    defparam bit_ctr_0__bdd_4_lut_53759_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 sub_67_add_2_11_lut (.I0(one_wire_N_479[8]), .I1(timer[9]), 
            .I2(n13[9]), .I3(n49557), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_53769_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n69493));
    defparam bit_ctr_0__bdd_4_lut_53769_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_54019_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n69505));
    defparam bit_ctr_0__bdd_4_lut_54019_4_lut.LUT_INIT = 16'heea0;
    SB_CARRY sub_67_add_2_11 (.CI(n49557), .I0(timer[9]), .I1(n13[9]), 
            .CO(n49558));
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n49556), .O(one_wire_N_479[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n49556), .I0(timer[8]), .I1(n13[8]), 
            .CO(n49557));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n49555), .O(one_wire_N_479[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n49555), .I0(timer[7]), .I1(n13[7]), 
            .CO(n49556));
    SB_LUT4 sub_67_add_2_8_lut (.I0(one_wire_N_479[10]), .I1(timer[6]), 
            .I2(n13[6]), .I3(n49554), .O(n7_adj_5667)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_8 (.CI(n49554), .I0(timer[6]), .I1(n13[6]), 
            .CO(n49555));
    SB_LUT4 sub_67_add_2_7_lut (.I0(n115), .I1(timer[5]), .I2(n13[5]), 
            .I3(n49553), .O(n6_adj_5668)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_7 (.CI(n49553), .I0(timer[5]), .I1(n13[5]), 
            .CO(n49554));
    SB_LUT4 sub_67_add_2_6_lut (.I0(n6_adj_5668), .I1(timer[4]), .I2(n13[4]), 
            .I3(n49552), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n69811));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_CARRY sub_67_add_2_6 (.CI(n49552), .I0(timer[4]), .I1(n13[4]), 
            .CO(n49553));
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n49551), .O(one_wire_N_479[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_5 (.CI(n49551), .I0(timer[3]), .I1(n13[3]), 
            .CO(n49552));
    SB_LUT4 i52_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr_c[3]), .I2(bit_ctr[1]), 
            .I3(GND_net), .O(n41_adj_5671));
    defparam i52_3_lut.LUT_INIT = 16'h2424;
    SB_LUT4 i3_4_lut (.I0(n52115), .I1(n41_adj_5671), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n23));
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i42488_2_lut (.I0(n23), .I1(n43567), .I2(GND_net), .I3(GND_net), 
            .O(n58165));
    defparam i42488_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n49550), .O(one_wire_N_479[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50624_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(one_wire_N_479[10]), 
            .I3(n115), .O(n65742));   // verilog/neopixel.v(34[12] 116[6])
    defparam i50624_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i2089_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6897));   // verilog/neopixel.v(68[23:32])
    defparam i2089_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15123_2_lut (.I0(n27950), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29199));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15123_2_lut.LUT_INIT = 16'h8888;
    SB_DFF timer_1938__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29707));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i50864_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n51632), 
            .I2(start), .I3(GND_net), .O(n65744));   // verilog/neopixel.v(16[11:16])
    defparam i50864_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(color_bit_N_502[1]), .I1(n63160), 
            .I2(n63161), .I3(color_bit_N_502[2]), .O(n69625));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n51632), 
            .I2(start), .I3(GND_net), .O(n111));   // verilog/neopixel.v(16[11:16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_CARRY sub_67_add_2_4 (.CI(n49550), .I0(timer[2]), .I1(n13[2]), 
            .CO(n49551));
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n27950), 
            .D(n137[2]), .R(n29199));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr_c[3]), .C(clk16MHz), .E(n27950), 
            .D(n137[3]), .R(n29199));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i4 (.Q(bit_ctr_c[4]), .C(clk16MHz), .E(n27950), 
            .D(n137[4]), .R(n29199));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF timer_1938__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i29486_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n43457));
    defparam i29486_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1970 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1970.LUT_INIT = 16'h1e1e;
    SB_LUT4 timer_1938_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n50777), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1938_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n50776), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_11 (.CI(n50776), .I0(GND_net), .I1(timer[9]), 
            .CO(n50777));
    SB_LUT4 timer_1938_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n50775), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_10 (.CI(n50775), .I0(GND_net), .I1(timer[8]), 
            .CO(n50776));
    SB_LUT4 timer_1938_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n50774), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_9 (.CI(n50774), .I0(GND_net), .I1(timer[7]), 
            .CO(n50775));
    SB_LUT4 timer_1938_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n50773), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_8 (.CI(n50773), .I0(GND_net), .I1(timer[6]), 
            .CO(n50774));
    SB_LUT4 timer_1938_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n50772), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_7 (.CI(n50772), .I0(GND_net), .I1(timer[5]), 
            .CO(n50773));
    SB_LUT4 timer_1938_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n50771), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_6 (.CI(n50771), .I0(GND_net), .I1(timer[4]), 
            .CO(n50772));
    SB_LUT4 timer_1938_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n50770), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_5 (.CI(n50770), .I0(GND_net), .I1(timer[3]), 
            .CO(n50771));
    SB_LUT4 timer_1938_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n50769), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_4 (.CI(n50769), .I0(GND_net), .I1(timer[2]), 
            .CO(n50770));
    SB_LUT4 timer_1938_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n50768), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_3 (.CI(n50768), .I0(GND_net), .I1(timer[1]), 
            .CO(n50769));
    SB_LUT4 timer_1938_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n50768));
    SB_LUT4 i47433_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n63161));
    defparam i47433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47432_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n63160));
    defparam i47432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_502[1]));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n30355));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n30354));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n30353));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n30352));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n30351));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n30350));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n30349));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n30348));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n30347));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n30342));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .D(n30251));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n5));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_add_2_3_lut (.I0(n4_adj_5674), .I1(timer[1]), .I2(n13[1]), 
            .I3(n49549), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1971 (.I0(one_wire_N_479[10]), .I1(n115), .I2(GND_net), 
            .I3(GND_net), .O(n41));
    defparam i1_2_lut_adj_1971.LUT_INIT = 16'h8888;
    SB_CARRY sub_67_add_2_3 (.CI(n49549), .I0(timer[1]), .I1(n13[1]), 
            .CO(n49550));
    SB_LUT4 i1_4_lut_adj_1972 (.I0(n75), .I1(n58296), .I2(n112), .I3(state[0]), 
            .O(n51632));   // verilog/neopixel.v(16[11:16])
    defparam i1_4_lut_adj_1972.LUT_INIT = 16'hfcee;
    SB_LUT4 i15_4_lut (.I0(n65744), .I1(n40890), .I2(state[1]), .I3(state[0]), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n49549));
    SB_LUT4 i53461_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 115[11])
    defparam i53461_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 n69625_bdd_4_lut (.I0(n69625), .I1(n63149), .I2(n63148), .I3(color_bit_N_502[2]), 
            .O(n69628));
    defparam n69625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n27940), .D(n1), 
            .R(n28911));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n27954), .D(state_1__N_440[0]), 
            .S(n29203));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n27707), .D(\neo_pixel_transmitter.done_N_524 ), 
            .R(n60566));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i1_4_lut_adj_1973 (.I0(n112), .I1(n59_adj_5675), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n33));
    defparam i1_4_lut_adj_1973.LUT_INIT = 16'hdccd;
    SB_LUT4 i1_4_lut_adj_1974 (.I0(state[1]), .I1(n33), .I2(n58296), .I3(start), 
            .O(n25));
    defparam i1_4_lut_adj_1974.LUT_INIT = 16'haaae;
    SB_LUT4 i1_3_lut (.I0(n75), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n59_adj_5675));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i42586_2_lut (.I0(one_wire_N_479[3]), .I1(one_wire_N_479[2]), 
            .I2(GND_net), .I3(GND_net), .O(n112));
    defparam i42586_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47420_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n63148));
    defparam i47420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47421_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n63149));
    defparam i47421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42614_2_lut (.I0(state[1]), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n58298));
    defparam i42614_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_4_lut (.I0(n111), .I1(state[1]), .I2(n40890), .I3(state[0]), 
            .O(n27954));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'heee2;
    SB_LUT4 i1_2_lut_3_lut_adj_1975 (.I0(n111), .I1(state[1]), .I2(n27940), 
            .I3(GND_net), .O(n27950));
    defparam i1_2_lut_3_lut_adj_1975.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(LED_c), .I2(n58165), .I3(state[1]), 
            .O(n27940));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 sub_67_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14835_2_lut_4_lut (.I0(state[0]), .I1(LED_c), .I2(n58165), 
            .I3(state[1]), .O(n28911));   // verilog/neopixel.v(34[12] 116[6])
    defparam i14835_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29593_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n43457), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n43567));
    defparam i29593_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1976 (.I0(bit_ctr_c[3]), .I1(n43457), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n52115));
    defparam i1_2_lut_3_lut_adj_1976.LUT_INIT = 16'h7878;
    SB_LUT4 i2108_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n6897), .I2(bit_ctr_c[3]), 
            .I3(bit_ctr_c[4]), .O(n137[4]));   // verilog/neopixel.v(68[23:32])
    defparam i2108_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i2101_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(bit_ctr_c[3]), .O(n137[3]));   // verilog/neopixel.v(68[23:32])
    defparam i2101_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53697_4_lut (.I0(n62744), .I1(n112), .I2(one_wire_N_479[7]), 
            .I3(n59_adj_5675), .O(n60559));
    defparam i53697_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i26894_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(16[11:16])
    defparam i26894_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i1_2_lut_adj_1977 (.I0(one_wire_N_479[2]), .I1(one_wire_N_479[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5674));
    defparam i1_2_lut_adj_1977.LUT_INIT = 16'h8888;
    SB_LUT4 sub_67_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1978 (.I0(\neo_pixel_transmitter.done ), .I1(one_wire_N_479[10]), 
            .I2(n115), .I3(GND_net), .O(n40890));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_3_lut_adj_1978.LUT_INIT = 16'h4040;
    SB_LUT4 i2094_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n137[2]));   // verilog/neopixel.v(68[23:32])
    defparam i2094_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n58296), .I3(n112), .O(n25554));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hbbbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1979 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n58296), .I3(n75), .O(n25553));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_3_lut_4_lut_adj_1979.LUT_INIT = 16'hbbbf;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n41), .I3(\neo_pixel_transmitter.done_N_524 ), 
            .O(n60566));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i50961_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n43457), .I2(n69628), 
            .I3(GND_net), .O(n65791));
    defparam i50961_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i52238_3_lut_4_lut (.I0(bit_ctr_c[3]), .I1(n43457), .I2(n63106), 
            .I3(n67842), .O(n67966));
    defparam i52238_3_lut_4_lut.LUT_INIT = 16'hf960;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i42712_2_lut_3_lut (.I0(state[1]), .I1(start), .I2(n58296), 
            .I3(GND_net), .O(n58397));
    defparam i42712_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n69811_bdd_4_lut (.I0(n69811), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_502[1]), .O(n69814));
    defparam n69811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69505_bdd_4_lut (.I0(n69505), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(color_bit_N_502[1]), .O(n69508));
    defparam n69505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69493_bdd_4_lut (.I0(n69493), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(color_bit_N_502[1]), .O(n69496));
    defparam n69493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69457_bdd_4_lut_4_lut (.I0(color_bit_N_502[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n69457), .O(n69460));   // verilog/neopixel.v(18[6:15])
    defparam n69457_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 i47025_2_lut_3_lut (.I0(n7_adj_5667), .I1(n8), .I2(n58298), 
            .I3(GND_net), .O(n62744));   // verilog/neopixel.v(101[14:24])
    defparam i47025_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i42612_2_lut_3_lut (.I0(n7_adj_5667), .I1(n8), .I2(one_wire_N_479[7]), 
            .I3(GND_net), .O(n58296));   // verilog/neopixel.v(101[14:24])
    defparam i42612_2_lut_3_lut.LUT_INIT = 16'hfefe;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (ENCODER1_B_N_keep, n1779, ENCODER1_A_N_keep, 
            \a_new[1] , n29731, n1784, position_31__N_3827, n1824, 
            n1786, n1788, n1790, n1792, n1794, n1796, \encoder1_position[25] , 
            \encoder1_position[24] , \encoder1_position[23] , \encoder1_position[22] , 
            \encoder1_position[21] , \encoder1_position[20] , \encoder1_position[19] , 
            \encoder1_position[18] , \encoder1_position[17] , \encoder1_position[16] , 
            \encoder1_position[15] , \encoder1_position[14] , \encoder1_position[13] , 
            \encoder1_position[12] , \encoder1_position[11] , \encoder1_position[10] , 
            \encoder1_position[9] , \encoder1_position[8] , \encoder1_position[7] , 
            \encoder1_position[6] , \encoder1_position[5] , \encoder1_position[4] , 
            \encoder1_position[3] , \encoder1_position[2] , n1822, GND_net, 
            VCC_net, b_prev) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1779;
    input ENCODER1_A_N_keep;
    output \a_new[1] ;
    input n29731;
    output n1784;
    output position_31__N_3827;
    output n1824;
    output n1786;
    output n1788;
    output n1790;
    output n1792;
    output n1794;
    output n1796;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    output \encoder1_position[3] ;
    output \encoder1_position[2] ;
    output n1822;
    input GND_net;
    input VCC_net;
    output b_prev;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3835, debounce_cnt, n29779, a_prev;
    wire [31:0]n133;
    
    wire direction_N_3832, n50900, n50899, n50898, n50897, n50896, 
        n50895, n50894, n50893, n50892, n50891, n50890, n50889, 
        n50888, n50887, n50886, n50885, n50884, n50883, n50882, 
        n50881, n50880, n50879, n50878, n50877, n50876, n50875, 
        n50874, n50873, n50872, n50871, n50870, n29507, position_31__N_3830;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1779), .D(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1779), .D(n29779));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i52948_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i52948_4_lut.LUT_INIT = 16'h8421;
    SB_DFF direction_40 (.Q(n1784), .C(n1779), .D(n29731));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1944__i0 (.Q(n1824), .C(n1779), .E(position_31__N_3827), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i31 (.Q(n1786), .C(n1779), .E(position_31__N_3827), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i30 (.Q(n1788), .C(n1779), .E(position_31__N_3827), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i29 (.Q(n1790), .C(n1779), .E(position_31__N_3827), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i28 (.Q(n1792), .C(n1779), .E(position_31__N_3827), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i27 (.Q(n1794), .C(n1779), .E(position_31__N_3827), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i26 (.Q(n1796), .C(n1779), .E(position_31__N_3827), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i25 (.Q(\encoder1_position[25] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i24 (.Q(\encoder1_position[24] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i23 (.Q(\encoder1_position[23] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i22 (.Q(\encoder1_position[22] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i21 (.Q(\encoder1_position[21] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i20 (.Q(\encoder1_position[20] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i19 (.Q(\encoder1_position[19] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i18 (.Q(\encoder1_position[18] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i17 (.Q(\encoder1_position[17] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i16 (.Q(\encoder1_position[16] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i15 (.Q(\encoder1_position[15] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i14 (.Q(\encoder1_position[14] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i13 (.Q(\encoder1_position[13] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i12 (.Q(\encoder1_position[12] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i11 (.Q(\encoder1_position[11] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i10 (.Q(\encoder1_position[10] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i9 (.Q(\encoder1_position[9] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i8 (.Q(\encoder1_position[8] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i7 (.Q(\encoder1_position[7] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i6 (.Q(\encoder1_position[6] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i5 (.Q(\encoder1_position[5] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i4 (.Q(\encoder1_position[4] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i3 (.Q(\encoder1_position[3] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i2 (.Q(\encoder1_position[2] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i1 (.Q(n1822), .C(n1779), .E(position_31__N_3827), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_1944_add_4_33_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1786), .I3(n50900), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1944_add_4_32_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1788), .I3(n50899), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_32 (.CI(n50899), .I0(direction_N_3832), 
            .I1(n1788), .CO(n50900));
    SB_LUT4 position_1944_add_4_31_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1790), .I3(n50898), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_31 (.CI(n50898), .I0(direction_N_3832), 
            .I1(n1790), .CO(n50899));
    SB_LUT4 position_1944_add_4_30_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1792), .I3(n50897), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_30 (.CI(n50897), .I0(direction_N_3832), 
            .I1(n1792), .CO(n50898));
    SB_LUT4 position_1944_add_4_29_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1794), .I3(n50896), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_29 (.CI(n50896), .I0(direction_N_3832), 
            .I1(n1794), .CO(n50897));
    SB_LUT4 position_1944_add_4_28_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1796), .I3(n50895), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_28 (.CI(n50895), .I0(direction_N_3832), 
            .I1(n1796), .CO(n50896));
    SB_LUT4 position_1944_add_4_27_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[25] ), .I3(n50894), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_27 (.CI(n50894), .I0(direction_N_3832), 
            .I1(\encoder1_position[25] ), .CO(n50895));
    SB_LUT4 position_1944_add_4_26_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[24] ), .I3(n50893), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_26 (.CI(n50893), .I0(direction_N_3832), 
            .I1(\encoder1_position[24] ), .CO(n50894));
    SB_LUT4 position_1944_add_4_25_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[23] ), .I3(n50892), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_25 (.CI(n50892), .I0(direction_N_3832), 
            .I1(\encoder1_position[23] ), .CO(n50893));
    SB_LUT4 position_1944_add_4_24_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[22] ), .I3(n50891), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_24 (.CI(n50891), .I0(direction_N_3832), 
            .I1(\encoder1_position[22] ), .CO(n50892));
    SB_LUT4 position_1944_add_4_23_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[21] ), .I3(n50890), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_23 (.CI(n50890), .I0(direction_N_3832), 
            .I1(\encoder1_position[21] ), .CO(n50891));
    SB_LUT4 position_1944_add_4_22_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[20] ), .I3(n50889), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_22 (.CI(n50889), .I0(direction_N_3832), 
            .I1(\encoder1_position[20] ), .CO(n50890));
    SB_LUT4 position_1944_add_4_21_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[19] ), .I3(n50888), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_21 (.CI(n50888), .I0(direction_N_3832), 
            .I1(\encoder1_position[19] ), .CO(n50889));
    SB_LUT4 position_1944_add_4_20_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[18] ), .I3(n50887), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_20 (.CI(n50887), .I0(direction_N_3832), 
            .I1(\encoder1_position[18] ), .CO(n50888));
    SB_LUT4 position_1944_add_4_19_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[17] ), .I3(n50886), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_19 (.CI(n50886), .I0(direction_N_3832), 
            .I1(\encoder1_position[17] ), .CO(n50887));
    SB_LUT4 position_1944_add_4_18_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[16] ), .I3(n50885), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_18 (.CI(n50885), .I0(direction_N_3832), 
            .I1(\encoder1_position[16] ), .CO(n50886));
    SB_LUT4 position_1944_add_4_17_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[15] ), .I3(n50884), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_17 (.CI(n50884), .I0(direction_N_3832), 
            .I1(\encoder1_position[15] ), .CO(n50885));
    SB_LUT4 position_1944_add_4_16_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[14] ), .I3(n50883), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_16 (.CI(n50883), .I0(direction_N_3832), 
            .I1(\encoder1_position[14] ), .CO(n50884));
    SB_LUT4 position_1944_add_4_15_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[13] ), .I3(n50882), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_15 (.CI(n50882), .I0(direction_N_3832), 
            .I1(\encoder1_position[13] ), .CO(n50883));
    SB_LUT4 position_1944_add_4_14_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[12] ), .I3(n50881), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_14 (.CI(n50881), .I0(direction_N_3832), 
            .I1(\encoder1_position[12] ), .CO(n50882));
    SB_LUT4 position_1944_add_4_13_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[11] ), .I3(n50880), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_13 (.CI(n50880), .I0(direction_N_3832), 
            .I1(\encoder1_position[11] ), .CO(n50881));
    SB_LUT4 position_1944_add_4_12_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[10] ), .I3(n50879), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_12 (.CI(n50879), .I0(direction_N_3832), 
            .I1(\encoder1_position[10] ), .CO(n50880));
    SB_LUT4 position_1944_add_4_11_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[9] ), .I3(n50878), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_11 (.CI(n50878), .I0(direction_N_3832), 
            .I1(\encoder1_position[9] ), .CO(n50879));
    SB_LUT4 position_1944_add_4_10_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[8] ), .I3(n50877), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_10 (.CI(n50877), .I0(direction_N_3832), 
            .I1(\encoder1_position[8] ), .CO(n50878));
    SB_LUT4 position_1944_add_4_9_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[7] ), .I3(n50876), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_9 (.CI(n50876), .I0(direction_N_3832), 
            .I1(\encoder1_position[7] ), .CO(n50877));
    SB_LUT4 position_1944_add_4_8_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[6] ), .I3(n50875), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_8 (.CI(n50875), .I0(direction_N_3832), 
            .I1(\encoder1_position[6] ), .CO(n50876));
    SB_LUT4 position_1944_add_4_7_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[5] ), .I3(n50874), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_7 (.CI(n50874), .I0(direction_N_3832), 
            .I1(\encoder1_position[5] ), .CO(n50875));
    SB_LUT4 position_1944_add_4_6_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[4] ), .I3(n50873), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_6 (.CI(n50873), .I0(direction_N_3832), 
            .I1(\encoder1_position[4] ), .CO(n50874));
    SB_LUT4 position_1944_add_4_5_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[3] ), .I3(n50872), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_5 (.CI(n50872), .I0(direction_N_3832), 
            .I1(\encoder1_position[3] ), .CO(n50873));
    SB_LUT4 position_1944_add_4_4_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[2] ), .I3(n50871), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_4 (.CI(n50871), .I0(direction_N_3832), 
            .I1(\encoder1_position[2] ), .CO(n50872));
    SB_LUT4 position_1944_add_4_3_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1822), .I3(n50870), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_3 (.CI(n50870), .I0(direction_N_3832), 
            .I1(n1822), .CO(n50871));
    SB_LUT4 position_1944_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1824), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n1824), 
            .CO(n50870));
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1779), .D(n29507));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3830));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3830), 
            .I3(\a_new[1] ), .O(position_31__N_3827));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3832));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i15703_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29779));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15431_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(b_new[1]), 
            .I3(b_prev), .O(n29507));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15431_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (ENCODER0_B_N_keep, n1779, ENCODER0_A_N_keep, 
            \a_new[1] , b_prev, n29751, n1742, position_31__N_3827, 
            n1744, \encoder0_position[30] , \encoder0_position[29] , \encoder0_position[28] , 
            \encoder0_position[27] , \encoder0_position[26] , \encoder0_position[25] , 
            \encoder0_position[24] , \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , GND_net, VCC_net) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1779;
    input ENCODER0_A_N_keep;
    output \a_new[1] ;
    output b_prev;
    input n29751;
    output n1742;
    output position_31__N_3827;
    output n1744;
    output \encoder0_position[30] ;
    output \encoder0_position[29] ;
    output \encoder0_position[28] ;
    output \encoder0_position[27] ;
    output \encoder0_position[26] ;
    output \encoder0_position[25] ;
    output \encoder0_position[24] ;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input GND_net;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3835, debounce_cnt, n29778, a_prev, n29777;
    wire [31:0]n133;
    
    wire direction_N_3832, n50964, n50963, n50962, n50961, n50960, 
        n50959, n50958, n50957, n50956, n50955, n50954, n50953, 
        n50952, n50951, n50950, n50949, n50948, n50947, n50946, 
        n50945, n50944, n50943, n50942, n50941, n50940, n50939, 
        n50938, n50937, n50936, n50935, n50934, position_31__N_3830;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1779), .D(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i52945_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i52945_4_lut.LUT_INIT = 16'h8421;
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1779), .D(n29778));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1779), .D(n29777));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n1742), .C(n1779), .D(n29751));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1956__i31 (.Q(n1744), .C(n1779), .E(position_31__N_3827), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i30 (.Q(\encoder0_position[30] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i29 (.Q(\encoder0_position[29] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i28 (.Q(\encoder0_position[28] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i27 (.Q(\encoder0_position[27] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i26 (.Q(\encoder0_position[26] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i25 (.Q(\encoder0_position[25] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i24 (.Q(\encoder0_position[24] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i23 (.Q(\encoder0_position[23] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i22 (.Q(\encoder0_position[22] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i21 (.Q(\encoder0_position[21] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i20 (.Q(\encoder0_position[20] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i19 (.Q(\encoder0_position[19] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i18 (.Q(\encoder0_position[18] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i17 (.Q(\encoder0_position[17] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i16 (.Q(\encoder0_position[16] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i15 (.Q(\encoder0_position[15] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i14 (.Q(\encoder0_position[14] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i13 (.Q(\encoder0_position[13] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i12 (.Q(\encoder0_position[12] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i11 (.Q(\encoder0_position[11] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i10 (.Q(\encoder0_position[10] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i9 (.Q(\encoder0_position[9] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i8 (.Q(\encoder0_position[8] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i7 (.Q(\encoder0_position[7] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i6 (.Q(\encoder0_position[6] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i5 (.Q(\encoder0_position[5] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i4 (.Q(\encoder0_position[4] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i3 (.Q(\encoder0_position[3] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i2 (.Q(\encoder0_position[2] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i1 (.Q(\encoder0_position[1] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i0 (.Q(\encoder0_position[0] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_1956_add_4_33_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1744), .I3(n50964), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1956_add_4_32_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[30] ), .I3(n50963), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_32 (.CI(n50963), .I0(direction_N_3832), 
            .I1(\encoder0_position[30] ), .CO(n50964));
    SB_LUT4 position_1956_add_4_31_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[29] ), .I3(n50962), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_31 (.CI(n50962), .I0(direction_N_3832), 
            .I1(\encoder0_position[29] ), .CO(n50963));
    SB_LUT4 position_1956_add_4_30_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[28] ), .I3(n50961), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_30 (.CI(n50961), .I0(direction_N_3832), 
            .I1(\encoder0_position[28] ), .CO(n50962));
    SB_LUT4 position_1956_add_4_29_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[27] ), .I3(n50960), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_29 (.CI(n50960), .I0(direction_N_3832), 
            .I1(\encoder0_position[27] ), .CO(n50961));
    SB_LUT4 position_1956_add_4_28_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[26] ), .I3(n50959), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_28 (.CI(n50959), .I0(direction_N_3832), 
            .I1(\encoder0_position[26] ), .CO(n50960));
    SB_LUT4 position_1956_add_4_27_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[25] ), .I3(n50958), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_27 (.CI(n50958), .I0(direction_N_3832), 
            .I1(\encoder0_position[25] ), .CO(n50959));
    SB_LUT4 position_1956_add_4_26_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[24] ), .I3(n50957), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_26 (.CI(n50957), .I0(direction_N_3832), 
            .I1(\encoder0_position[24] ), .CO(n50958));
    SB_LUT4 position_1956_add_4_25_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[23] ), .I3(n50956), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_25 (.CI(n50956), .I0(direction_N_3832), 
            .I1(\encoder0_position[23] ), .CO(n50957));
    SB_LUT4 position_1956_add_4_24_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[22] ), .I3(n50955), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_24 (.CI(n50955), .I0(direction_N_3832), 
            .I1(\encoder0_position[22] ), .CO(n50956));
    SB_LUT4 position_1956_add_4_23_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[21] ), .I3(n50954), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_23 (.CI(n50954), .I0(direction_N_3832), 
            .I1(\encoder0_position[21] ), .CO(n50955));
    SB_LUT4 position_1956_add_4_22_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[20] ), .I3(n50953), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_22 (.CI(n50953), .I0(direction_N_3832), 
            .I1(\encoder0_position[20] ), .CO(n50954));
    SB_LUT4 position_1956_add_4_21_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[19] ), .I3(n50952), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_21 (.CI(n50952), .I0(direction_N_3832), 
            .I1(\encoder0_position[19] ), .CO(n50953));
    SB_LUT4 position_1956_add_4_20_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[18] ), .I3(n50951), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_20 (.CI(n50951), .I0(direction_N_3832), 
            .I1(\encoder0_position[18] ), .CO(n50952));
    SB_LUT4 position_1956_add_4_19_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[17] ), .I3(n50950), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_19 (.CI(n50950), .I0(direction_N_3832), 
            .I1(\encoder0_position[17] ), .CO(n50951));
    SB_LUT4 position_1956_add_4_18_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[16] ), .I3(n50949), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_18 (.CI(n50949), .I0(direction_N_3832), 
            .I1(\encoder0_position[16] ), .CO(n50950));
    SB_LUT4 position_1956_add_4_17_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[15] ), .I3(n50948), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_17 (.CI(n50948), .I0(direction_N_3832), 
            .I1(\encoder0_position[15] ), .CO(n50949));
    SB_LUT4 position_1956_add_4_16_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[14] ), .I3(n50947), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_16 (.CI(n50947), .I0(direction_N_3832), 
            .I1(\encoder0_position[14] ), .CO(n50948));
    SB_LUT4 position_1956_add_4_15_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[13] ), .I3(n50946), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_15 (.CI(n50946), .I0(direction_N_3832), 
            .I1(\encoder0_position[13] ), .CO(n50947));
    SB_LUT4 position_1956_add_4_14_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[12] ), .I3(n50945), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_14 (.CI(n50945), .I0(direction_N_3832), 
            .I1(\encoder0_position[12] ), .CO(n50946));
    SB_LUT4 position_1956_add_4_13_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[11] ), .I3(n50944), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_13 (.CI(n50944), .I0(direction_N_3832), 
            .I1(\encoder0_position[11] ), .CO(n50945));
    SB_LUT4 position_1956_add_4_12_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[10] ), .I3(n50943), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_12 (.CI(n50943), .I0(direction_N_3832), 
            .I1(\encoder0_position[10] ), .CO(n50944));
    SB_LUT4 position_1956_add_4_11_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[9] ), .I3(n50942), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_11 (.CI(n50942), .I0(direction_N_3832), 
            .I1(\encoder0_position[9] ), .CO(n50943));
    SB_LUT4 position_1956_add_4_10_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[8] ), .I3(n50941), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_10 (.CI(n50941), .I0(direction_N_3832), 
            .I1(\encoder0_position[8] ), .CO(n50942));
    SB_LUT4 position_1956_add_4_9_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[7] ), .I3(n50940), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_9 (.CI(n50940), .I0(direction_N_3832), 
            .I1(\encoder0_position[7] ), .CO(n50941));
    SB_LUT4 position_1956_add_4_8_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[6] ), .I3(n50939), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_8 (.CI(n50939), .I0(direction_N_3832), 
            .I1(\encoder0_position[6] ), .CO(n50940));
    SB_LUT4 position_1956_add_4_7_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[5] ), .I3(n50938), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_7 (.CI(n50938), .I0(direction_N_3832), 
            .I1(\encoder0_position[5] ), .CO(n50939));
    SB_LUT4 position_1956_add_4_6_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[4] ), .I3(n50937), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_6 (.CI(n50937), .I0(direction_N_3832), 
            .I1(\encoder0_position[4] ), .CO(n50938));
    SB_LUT4 position_1956_add_4_5_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[3] ), .I3(n50936), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_5 (.CI(n50936), .I0(direction_N_3832), 
            .I1(\encoder0_position[3] ), .CO(n50937));
    SB_LUT4 position_1956_add_4_4_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[2] ), .I3(n50935), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_4 (.CI(n50935), .I0(direction_N_3832), 
            .I1(\encoder0_position[2] ), .CO(n50936));
    SB_LUT4 position_1956_add_4_3_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[1] ), .I3(n50934), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_3 (.CI(n50934), .I0(direction_N_3832), 
            .I1(\encoder0_position[1] ), .CO(n50935));
    SB_LUT4 position_1956_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n50934));
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3830));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3830), 
            .I3(\a_new[1] ), .O(position_31__N_3827));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3832));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i15702_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29778));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15702_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15701_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(b_new[1]), 
            .I3(b_prev), .O(n29777));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15701_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\state[1] , clk16MHz, clk_out, CS_c, CS_CLK_c, GND_net, 
            n15, \state[0] , n11, n29691, \data[15] , n9, n29677, 
            n29675, \current[0] , n29672, \data[12] , n29671, \data[11] , 
            n29656, \data[10] , n29655, \data[9] , n29654, \data[8] , 
            n29653, \data[7] , n29652, \data[6] , n29645, \data[5] , 
            n29637, \data[4] , n29636, \data[3] , n29635, \data[2] , 
            n29628, \data[1] , VCC_net, n30538, \data[0] , n30427, 
            \current[1] , n30426, \current[2] , n30425, \current[3] , 
            n30424, \current[4] , n30423, \current[5] , n30422, \current[6] , 
            n30421, \current[7] , n30420, \current[8] , n30419, \current[9] , 
            n30418, \current[10] , n30417, \current[11] , n6, n27736, 
            \current[15] , n5, n6_adj_31, state_7__N_4317, n42880, 
            n25615, n25587, n25590, n25578, n25583, n6_adj_32, n5_adj_33) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[1] ;
    input clk16MHz;
    output clk_out;
    output CS_c;
    output CS_CLK_c;
    input GND_net;
    output n15;
    output \state[0] ;
    output n11;
    input n29691;
    output \data[15] ;
    input n9;
    input n29677;
    input n29675;
    output \current[0] ;
    input n29672;
    output \data[12] ;
    input n29671;
    output \data[11] ;
    input n29656;
    output \data[10] ;
    input n29655;
    output \data[9] ;
    input n29654;
    output \data[8] ;
    input n29653;
    output \data[7] ;
    input n29652;
    output \data[6] ;
    input n29645;
    output \data[5] ;
    input n29637;
    output \data[4] ;
    input n29636;
    output \data[3] ;
    input n29635;
    output \data[2] ;
    input n29628;
    output \data[1] ;
    input VCC_net;
    input n30538;
    output \data[0] ;
    input n30427;
    output \current[1] ;
    input n30426;
    output \current[2] ;
    input n30425;
    output \current[3] ;
    input n30424;
    output \current[4] ;
    input n30423;
    output \current[5] ;
    input n30422;
    output \current[6] ;
    input n30421;
    output \current[7] ;
    input n30420;
    output \current[8] ;
    input n30419;
    output \current[9] ;
    input n30418;
    output \current[10] ;
    input n30417;
    output \current[11] ;
    output n6;
    output n27736;
    output \current[15] ;
    output n5;
    output n6_adj_31;
    output state_7__N_4317;
    output n42880;
    output n25615;
    output n25587;
    output n25590;
    output n25578;
    output n25583;
    output n6_adj_32;
    output n5_adj_33;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n12183, n28019, n28917, clk_slow_N_4230, n42933, n2;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n65610, n22642, n65659, n22640, n65671, n22638, n22636, 
        n27792;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire delay_counter_15__N_4312;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4231;
    wire [7:0]n37;
    
    wire n29189, n50913, n50912, n50911, n50910, n50909, n50908, 
        n50907, n50906, n50905, n50904, n50903, n50902, n50901, 
        n65672, n50807, n50806, n50805, n50804, n50803, n50802, 
        n50801;
    wire [1:0]n1859;
    
    wire n8, n12, n10, n6_adj_5666;
    
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n28019), .D(n12183), 
            .R(n28917));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4230));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i52957_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n42933));
    defparam i52957_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2397_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));
    defparam i2397_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 equal_264_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_264_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8832_3_lut (.I0(\state[0] ), .I1(n65610), .I2(\state[1] ), 
            .I3(GND_net), .O(n22642));   // verilog/tli4970.v(55[24:39])
    defparam i8832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8830_3_lut (.I0(\state[0] ), .I1(n65659), .I2(\state[1] ), 
            .I3(GND_net), .O(n22640));   // verilog/tli4970.v(55[24:39])
    defparam i8830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8828_3_lut (.I0(\state[0] ), .I1(n65671), .I2(\state[1] ), 
            .I3(GND_net), .O(n22638));   // verilog/tli4970.v(55[24:39])
    defparam i8828_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29691));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29677));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29675));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29672));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29671));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29656));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29655));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29654));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29653));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29652));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29645));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29637));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29636));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29635));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29628));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_1940__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27792), 
            .D(n22636));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_1946_1947__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1948_1949__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1948_1949__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1948_1949__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_1946_1947__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNESR bit_counter_1940__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27792), 
            .D(n37[4]), .R(n29189));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1940__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27792), 
            .D(n37[5]), .R(n29189));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1940__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27792), 
            .D(n37[6]), .R(n29189));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1940__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27792), 
            .D(n37[7]), .R(n29189));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1940__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27792), 
            .D(n22638));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1940__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27792), 
            .D(n22640));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1940__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27792), 
            .D(n22642));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 counter_1948_1949_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n50913), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1948_1949_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1948_1949_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n50912), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1948_1949_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1948_1949_add_4_3 (.CI(n50912), .I0(GND_net), .I1(counter[1]), 
            .CO(n50913));
    SB_LUT4 counter_1948_1949_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1948_1949_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1948_1949_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n50912));
    SB_LUT4 delay_counter_1946_1947_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n50911), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1946_1947_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n50910), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_12 (.CI(n50910), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n50911));
    SB_LUT4 delay_counter_1946_1947_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n50909), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_11 (.CI(n50909), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n50910));
    SB_LUT4 delay_counter_1946_1947_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n50908), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_10 (.CI(n50908), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n50909));
    SB_LUT4 delay_counter_1946_1947_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n50907), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_9 (.CI(n50907), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n50908));
    SB_LUT4 delay_counter_1946_1947_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n50906), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_8 (.CI(n50906), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n50907));
    SB_LUT4 delay_counter_1946_1947_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n50905), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_7 (.CI(n50905), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n50906));
    SB_LUT4 delay_counter_1946_1947_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n50904), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_6 (.CI(n50904), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n50905));
    SB_LUT4 delay_counter_1946_1947_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n50903), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_5 (.CI(n50903), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n50904));
    SB_LUT4 delay_counter_1946_1947_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n50902), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_4 (.CI(n50902), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n50903));
    SB_LUT4 delay_counter_1946_1947_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n50901), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_3 (.CI(n50901), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n50902));
    SB_LUT4 delay_counter_1946_1947_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n50901));
    SB_LUT4 i13985_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27792));
    defparam i13985_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8826_3_lut (.I0(\state[0] ), .I1(n65672), .I2(\state[1] ), 
            .I3(GND_net), .O(n22636));   // verilog/tli4970.v(55[24:39])
    defparam i8826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_counter_1940_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n50807), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_1940_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n50806), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1940_add_4_8 (.CI(n50806), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n50807));
    SB_LUT4 bit_counter_1940_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n50805), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1940_add_4_7 (.CI(n50805), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n50806));
    SB_LUT4 bit_counter_1940_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n50804), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1940_add_4_6 (.CI(n50804), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n50805));
    SB_LUT4 bit_counter_1940_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n50803), .O(n65671)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_5 (.CI(n50803), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n50804));
    SB_LUT4 bit_counter_1940_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n50802), .O(n65659)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_4 (.CI(n50802), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n50803));
    SB_LUT4 bit_counter_1940_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n50801), .O(n65610)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_3 (.CI(n50801), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n50802));
    SB_LUT4 bit_counter_1940_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n65672)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n50801));
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30538));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30427));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30426));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30425));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30424));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30423));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30422));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30421));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30420));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30419));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30418));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30417));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_333_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_333_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27736), 
            .D(n1859[0]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_324_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_324_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_328_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_31));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i52936_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n27736));
    defparam i52936_3_lut.LUT_INIT = 16'h4040;
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n28019), .D(n42933), 
            .S(n28917));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4317));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28912_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n42880));
    defparam i28912_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2121_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1859[0]));
    defparam i2121_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25615));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1964 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25587));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1964.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1965 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25590));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_1965.LUT_INIT = 16'hfbff;
    SB_LUT4 i15114_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29189));   // verilog/tli4970.v(55[24:39])
    defparam i15114_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2065_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4231));
    defparam i2065_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4231), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4230));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1966 (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4312), .O(n28019));
    defparam i1_2_lut_4_lut_adj_1966.LUT_INIT = 16'hffdc;
    SB_LUT4 i14841_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4312), .O(n28917));
    defparam i14841_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25578));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1967 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n25583));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1967.LUT_INIT = 16'hffbf;
    SB_LUT4 equal_335_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_32));   // verilog/tli4970.v(54[9:26])
    defparam equal_335_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_326_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_33));   // verilog/tli4970.v(54[9:26])
    defparam equal_326_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2066_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2066_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(delay_counter[11]), .I1(delay_counter[7]), .I2(delay_counter[8]), 
            .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4312));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5666));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1968 (.I0(bit_counter[6]), .I1(bit_counter[7]), 
            .I2(n11), .I3(n6_adj_5666), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut_adj_1968.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_2033_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n12183));
    defparam mux_2033_i2_3_lut.LUT_INIT = 16'h3535;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n56422, \data_in_frame[22] , clk16MHz, VCC_net, \data_in_frame[4] , 
            GND_net, n2873, rx_data, \data_in_frame[5] , \data_in_frame[3] , 
            n7, \data_in_frame[9] , n29989, n29986, n29983, n56418, 
            n29979, n29976, n56414, \data_in_frame[3][6] , \data_in_frame[3][4] , 
            \data_in_frame[3][3] , \data_in_frame[3][2] , n29701, \data_in_frame[0][1] , 
            \data_in_frame[3][1] , \data_in_frame[3][0] , \data_in_frame[2] , 
            n56410, \data_in_frame[10] , n58117, \data_in_frame[1] , 
            \data_in_frame[0][7] , Kp_23__N_1748, reset, n56406, setpoint, 
            n56402, \data_in_frame[8] , \data_in_frame[12] , n57657, 
            \byte_transmit_counter[0] , \byte_transmit_counter[2] , \byte_transmit_counter[1] , 
            \data_in_frame[14] , n6, n69640, n43, n379, n405, n4, 
            pwm_setpoint, n29714, encoder0_position_scaled, n459, n11610, 
            n37308, n57425, n56398, \FRAME_MATCHER.i[4] , \FRAME_MATCHER.i[5] , 
            \FRAME_MATCHER.i[3] , DE_c, n29739, \data_in_frame[0][2] , 
            LED_c, n33801, \FRAME_MATCHER.i_31__N_2513 , n27726, \data_in_frame[17] , 
            \data_in_frame[15] , \data_in_frame[13] , n29764, \data_in_frame[0][3] , 
            \data_out_frame[20] , n29802, deadband, n29879, n29878, 
            n29877, n29876, n29875, n29874, n29873, n29872, n29871, 
            n29870, n29869, n29868, n29867, n29866, n29865, n29864, 
            n29863, n29862, n29861, n29860, n29859, n29858, n29857, 
            IntegralLimit, n29856, n29855, n29854, n29853, n53095, 
            n52011, n29852, n29851, n57836, \data_out_frame[18][3] , 
            n3470, rx_data_ready, \FRAME_MATCHER.rx_data_ready_prev , 
            \data_out_frame[23][3] , \data_out_frame[16][3] , n29850, 
            n29849, n29848, n29847, \data_out_frame[25][2] , n29846, 
            n29845, n29844, n29843, \data_in_frame[0][0] , n29842, 
            n29841, n29840, n29839, n29838, n29837, n29836, n29835, 
            n29834, \Kp[1] , \data_out_frame[24][2] , n29833, \Kp[2] , 
            n29832, \Kp[3] , n29831, \Kp[4] , n29830, \Kp[5] , n29829, 
            \Kp[6] , n57437, \Kp[7] , n29827, \Kp[8] , n29826, \Kp[9] , 
            n29825, \Kp[10] , n29824, \Kp[11] , n172, \data_out_frame[20][3] , 
            n29823, \Kp[12] , n29822, \Kp[13] , n28413, n29821, 
            \Kp[14] , n29820, \Kp[15] , n29819, \Ki[1] , n29818, 
            \Ki[2] , n29817, \Ki[3] , n29816, \Ki[4] , n29815, \Ki[5] , 
            n29814, \Ki[6] , n29813, \Ki[7] , n29812, \Ki[8] , n29811, 
            \Ki[9] , n29810, \Ki[10] , n29809, \Ki[11] , n29808, 
            \Ki[12] , n29807, \Ki[13] , \Ki[14] , n29805, \Ki[15] , 
            \data_in_frame[16] , n105, \data_out_frame[18][4] , \data_out_frame[17][3] , 
            n25848, n29767, n26517, n29760, neopxl_color, n29759, 
            current_limit, n29758, control_mode, n29757, n29756, n29755, 
            n29754, n29753, n29752, n29750, n29749, n29748, n29747, 
            n29746, n29745, n29744, n29743, n29742, n161, n31, 
            \data_out_frame[19][3] , n29738, n7_adj_10, n29735, encoder1_position_scaled, 
            n29734, n29733, n29732, n25, n29730, n29729, n29725, 
            n29721, n29718, \data_out_frame[22][3] , n57879, n59684, 
            n57499, n29700, n29699, n29692, n29673, PWMLimit, n29664, 
            n29663, n29662, n29661, \Ki[0] , n29660, \Kp[0] , n29644, 
            \data_in_frame[18] , \pwm_counter[22] , n45, \pwm_counter[21] , 
            n43_adj_11, \data_out_frame[21][0] , \data_out_frame[21][3] , 
            \data_in_frame[19] , n53127, \data_in_frame[21] , \current[7] , 
            \current[6] , n29471, n30549, n30548, n30547, n30546, 
            n30545, n30544, n30543, n29474, n30534, n29477, n30512, 
            n30506, n30504, n30503, n30501, n30500, n30499, n30498, 
            n30490, n30439, n30431, n30429, n30428, n30415, tx_active, 
            n30383, n30382, n30381, n30380, n30378, n56568, n30372, 
            n30371, n56566, n29520, n29523, n29526, n29530, n56478, 
            n56474, n56470, n56466, n56462, n56458, n30343, n56454, 
            n56450, n56446, \data_in_frame[6] , n30336, n30055, \data_in_frame[7][1] , 
            n30059, \data_in_frame[7][2] , n30062, \data_in_frame[7][3] , 
            n30065, \data_in_frame[7][4] , n30068, \data_in_frame[7][5] , 
            n30077, n30080, n30083, n30317, n30316, n30087, n30314, 
            n30093, n30096, n30099, n30102, n30105, n30108, n30112, 
            n30115, n30118, n30122, n30125, n30131, \data_in_frame[10][1] , 
            n30134, \data_in_frame[10][2] , n30138, \data_in_frame[10][3] , 
            n30141, n30144, \data_in_frame[10][5] , n30148, n30151, 
            \data_in_frame[10][7] , n30154, \data_in_frame[11] , n56662, 
            n56678, n56604, n30167, n30170, n30173, n30287, n30177, 
            n30180, n30183, n30186, n56636, n56690, n30196, n30199, 
            n30203, n56442, n56438, \current[5] , n30265, n29570, 
            n29573, n29576, n56434, n56430, n56546, n56542, \current[4] , 
            \current[3] , n56540, n29594, n56538, n56536, n56534, 
            n29609, \data_in_frame[20] , n29618, n29621, \current[2] , 
            \current[1] , n29624, \current[0] , n30176, \current[15] , 
            n29632, n8, \current[11] , \current[10] , \current[9] , 
            \current[8] , displacement, n8_adj_12, n57426, n29536, 
            n57956, n8_adj_13, n57424, n380, n460, n27722, n29510, 
            n33, n38, n34, n57990, n57737, n33793, n29508, n52054, 
            n58132, n53024, n57862, n52186, n57625, n57410, n28409, 
            n53215, \data_out_frame[26][2] , \data_out_frame[27][2] , 
            n29999, n22792, n35, n4_adj_14, Kp_23__N_1389, n57685, 
            n8_adj_15, n4_adj_16, ID, n15, n15_adj_17, n19, n28464, 
            n91, n58278, n7_adj_18, n26, n21, n260, n41114, n59370, 
            n69808, n63007, n63008, n63155, n63154, n30, n365, 
            n32, n65564, tx_o, r_SM_Main, n29690, n58304, r_Clock_Count, 
            n6_adj_19, n4940, n27, tx_enable, baudrate, \r_SM_Main[2]_adj_20 , 
            r_Rx_Data, RX_N_2, n4937, \o_Rx_DV_N_3488[8] , n61106, 
            n29912, n61058, n57317, \r_SM_Main[1]_adj_21 , n27754, 
            n61138, n29900, n25593, n29798, n29797, n29796, \r_Bit_Index[0] , 
            r_Clock_Count_adj_30, n27996, n58373, n30533, n53222, 
            n30529, n30231, n30230, \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , 
            n61170, n61154, n61090, n61074, n61122) /* synthesis syn_module_defined=1 */ ;
    input n56422;
    output [7:0]\data_in_frame[22] ;
    input clk16MHz;
    input VCC_net;
    output [7:0]\data_in_frame[4] ;
    input GND_net;
    output n2873;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[3] ;
    output n7;
    output [7:0]\data_in_frame[9] ;
    input n29989;
    input n29986;
    input n29983;
    input n56418;
    input n29979;
    input n29976;
    input n56414;
    output \data_in_frame[3][6] ;
    output \data_in_frame[3][4] ;
    output \data_in_frame[3][3] ;
    output \data_in_frame[3][2] ;
    input n29701;
    output \data_in_frame[0][1] ;
    output \data_in_frame[3][1] ;
    output \data_in_frame[3][0] ;
    output [7:0]\data_in_frame[2] ;
    input n56410;
    output [7:0]\data_in_frame[10] ;
    output n58117;
    output [7:0]\data_in_frame[1] ;
    output \data_in_frame[0][7] ;
    output Kp_23__N_1748;
    input reset;
    input n56406;
    output [23:0]setpoint;
    input n56402;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[12] ;
    output n57657;
    output \byte_transmit_counter[0] ;
    output \byte_transmit_counter[2] ;
    output \byte_transmit_counter[1] ;
    output [7:0]\data_in_frame[14] ;
    output n6;
    input n69640;
    input n43;
    input n379;
    input n405;
    output n4;
    input [23:0]pwm_setpoint;
    input n29714;
    input [23:0]encoder0_position_scaled;
    input n459;
    input n11610;
    output n37308;
    output n57425;
    input n56398;
    output \FRAME_MATCHER.i[4] ;
    output \FRAME_MATCHER.i[5] ;
    output \FRAME_MATCHER.i[3] ;
    output DE_c;
    input n29739;
    output \data_in_frame[0][2] ;
    output LED_c;
    output n33801;
    output \FRAME_MATCHER.i_31__N_2513 ;
    output n27726;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_in_frame[15] ;
    output [7:0]\data_in_frame[13] ;
    input n29764;
    output \data_in_frame[0][3] ;
    output [7:0]\data_out_frame[20] ;
    input n29802;
    output [23:0]deadband;
    input n29879;
    input n29878;
    input n29877;
    input n29876;
    input n29875;
    input n29874;
    input n29873;
    input n29872;
    input n29871;
    input n29870;
    input n29869;
    input n29868;
    input n29867;
    input n29866;
    input n29865;
    input n29864;
    input n29863;
    input n29862;
    input n29861;
    input n29860;
    input n29859;
    input n29858;
    input n29857;
    output [23:0]IntegralLimit;
    input n29856;
    input n29855;
    input n29854;
    input n29853;
    output n53095;
    input n52011;
    input n29852;
    input n29851;
    output n57836;
    output \data_out_frame[18][3] ;
    output n3470;
    output rx_data_ready;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output \data_out_frame[23][3] ;
    output \data_out_frame[16][3] ;
    input n29850;
    input n29849;
    input n29848;
    input n29847;
    output \data_out_frame[25][2] ;
    input n29846;
    input n29845;
    input n29844;
    input n29843;
    output \data_in_frame[0][0] ;
    input n29842;
    input n29841;
    input n29840;
    input n29839;
    input n29838;
    input n29837;
    input n29836;
    input n29835;
    input n29834;
    output \Kp[1] ;
    output \data_out_frame[24][2] ;
    input n29833;
    output \Kp[2] ;
    input n29832;
    output \Kp[3] ;
    input n29831;
    output \Kp[4] ;
    input n29830;
    output \Kp[5] ;
    input n29829;
    output \Kp[6] ;
    output n57437;
    output \Kp[7] ;
    input n29827;
    output \Kp[8] ;
    input n29826;
    output \Kp[9] ;
    input n29825;
    output \Kp[10] ;
    input n29824;
    output \Kp[11] ;
    output n172;
    output \data_out_frame[20][3] ;
    input n29823;
    output \Kp[12] ;
    input n29822;
    output \Kp[13] ;
    output n28413;
    input n29821;
    output \Kp[14] ;
    input n29820;
    output \Kp[15] ;
    input n29819;
    output \Ki[1] ;
    input n29818;
    output \Ki[2] ;
    input n29817;
    output \Ki[3] ;
    input n29816;
    output \Ki[4] ;
    input n29815;
    output \Ki[5] ;
    input n29814;
    output \Ki[6] ;
    input n29813;
    output \Ki[7] ;
    input n29812;
    output \Ki[8] ;
    input n29811;
    output \Ki[9] ;
    input n29810;
    output \Ki[10] ;
    input n29809;
    output \Ki[11] ;
    input n29808;
    output \Ki[12] ;
    input n29807;
    output \Ki[13] ;
    output \Ki[14] ;
    input n29805;
    output \Ki[15] ;
    output [7:0]\data_in_frame[16] ;
    output n105;
    output \data_out_frame[18][4] ;
    output \data_out_frame[17][3] ;
    input n25848;
    input n29767;
    output n26517;
    input n29760;
    output [23:0]neopxl_color;
    input n29759;
    output [15:0]current_limit;
    input n29758;
    output [7:0]control_mode;
    input n29757;
    input n29756;
    input n29755;
    input n29754;
    input n29753;
    input n29752;
    input n29750;
    input n29749;
    input n29748;
    input n29747;
    input n29746;
    input n29745;
    input n29744;
    input n29743;
    input n29742;
    output n161;
    output n31;
    output \data_out_frame[19][3] ;
    input n29738;
    output n7_adj_10;
    input n29735;
    input [23:0]encoder1_position_scaled;
    input n29734;
    input n29733;
    input n29732;
    input n25;
    input n29730;
    input n29729;
    input n29725;
    input n29721;
    input n29718;
    output \data_out_frame[22][3] ;
    output n57879;
    input n59684;
    output n57499;
    input n29700;
    input n29699;
    input n29692;
    input n29673;
    output [23:0]PWMLimit;
    input n29664;
    input n29663;
    input n29662;
    input n29661;
    output \Ki[0] ;
    input n29660;
    output \Kp[0] ;
    input n29644;
    output [7:0]\data_in_frame[18] ;
    input \pwm_counter[22] ;
    output n45;
    input \pwm_counter[21] ;
    output n43_adj_11;
    output \data_out_frame[21][0] ;
    output \data_out_frame[21][3] ;
    output [7:0]\data_in_frame[19] ;
    input n53127;
    output [7:0]\data_in_frame[21] ;
    input \current[7] ;
    input \current[6] ;
    input n29471;
    input n30549;
    input n30548;
    input n30547;
    input n30546;
    input n30545;
    input n30544;
    input n30543;
    input n29474;
    input n30534;
    input n29477;
    input n30512;
    input n30506;
    input n30504;
    input n30503;
    input n30501;
    input n30500;
    input n30499;
    input n30498;
    input n30490;
    input n30439;
    input n30431;
    input n30429;
    input n30428;
    input n30415;
    output tx_active;
    input n30383;
    input n30382;
    input n30381;
    input n30380;
    input n30378;
    input n56568;
    input n30372;
    input n30371;
    input n56566;
    input n29520;
    input n29523;
    input n29526;
    input n29530;
    input n56478;
    input n56474;
    input n56470;
    input n56466;
    input n56462;
    input n56458;
    input n30343;
    input n56454;
    input n56450;
    input n56446;
    output [7:0]\data_in_frame[6] ;
    input n30336;
    input n30055;
    output \data_in_frame[7][1] ;
    input n30059;
    output \data_in_frame[7][2] ;
    input n30062;
    output \data_in_frame[7][3] ;
    input n30065;
    output \data_in_frame[7][4] ;
    input n30068;
    output \data_in_frame[7][5] ;
    input n30077;
    input n30080;
    input n30083;
    input n30317;
    input n30316;
    input n30087;
    input n30314;
    input n30093;
    input n30096;
    input n30099;
    input n30102;
    input n30105;
    input n30108;
    input n30112;
    input n30115;
    input n30118;
    input n30122;
    input n30125;
    input n30131;
    output \data_in_frame[10][1] ;
    input n30134;
    output \data_in_frame[10][2] ;
    input n30138;
    output \data_in_frame[10][3] ;
    input n30141;
    input n30144;
    output \data_in_frame[10][5] ;
    input n30148;
    input n30151;
    output \data_in_frame[10][7] ;
    input n30154;
    output [7:0]\data_in_frame[11] ;
    input n56662;
    input n56678;
    input n56604;
    input n30167;
    input n30170;
    input n30173;
    input n30287;
    input n30177;
    input n30180;
    input n30183;
    input n30186;
    input n56636;
    input n56690;
    input n30196;
    input n30199;
    input n30203;
    input n56442;
    input n56438;
    input \current[5] ;
    input n30265;
    input n29570;
    input n29573;
    input n29576;
    input n56434;
    input n56430;
    input n56546;
    input n56542;
    input \current[4] ;
    input \current[3] ;
    input n56540;
    input n29594;
    input n56538;
    input n56536;
    input n56534;
    input n29609;
    output [7:0]\data_in_frame[20] ;
    input n29618;
    input n29621;
    input \current[2] ;
    input \current[1] ;
    input n29624;
    input \current[0] ;
    input n30176;
    input \current[15] ;
    input n29632;
    output n8;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input [23:0]displacement;
    output n8_adj_12;
    output n57426;
    input n29536;
    output n57956;
    output n8_adj_13;
    output n57424;
    input n380;
    input n460;
    output n27722;
    input n29510;
    input n33;
    input n38;
    input n34;
    output n57990;
    output n57737;
    output n33793;
    input n29508;
    output n52054;
    output n58132;
    output n53024;
    output n57862;
    output n52186;
    output n57625;
    output n57410;
    output n28409;
    output n53215;
    output \data_out_frame[26][2] ;
    output \data_out_frame[27][2] ;
    input n29999;
    input n22792;
    input n35;
    output n4_adj_14;
    output Kp_23__N_1389;
    output n57685;
    output n8_adj_15;
    output n4_adj_16;
    input [7:0]ID;
    input n15;
    input n15_adj_17;
    output n19;
    output n28464;
    input n91;
    output n58278;
    output n7_adj_18;
    input n26;
    output n21;
    output n260;
    output n41114;
    output n59370;
    output n69808;
    input n63007;
    input n63008;
    input n63155;
    input n63154;
    input n30;
    input n365;
    output n32;
    input n65564;
    output tx_o;
    output [2:0]r_SM_Main;
    input n29690;
    input n58304;
    output [8:0]r_Clock_Count;
    output n6_adj_19;
    input n4940;
    output n27;
    output tx_enable;
    input [31:0]baudrate;
    output \r_SM_Main[2]_adj_20 ;
    output r_Rx_Data;
    input RX_N_2;
    input n4937;
    output \o_Rx_DV_N_3488[8] ;
    output n61106;
    input n29912;
    output n61058;
    input n57317;
    output \r_SM_Main[1]_adj_21 ;
    output n27754;
    output n61138;
    input n29900;
    output n25593;
    input n29798;
    input n29797;
    input n29796;
    output \r_Bit_Index[0] ;
    output [7:0]r_Clock_Count_adj_30;
    output n27996;
    output n58373;
    input n30533;
    input n53222;
    input n30529;
    input n30231;
    input n30230;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n61170;
    output n61154;
    output n61090;
    output n61074;
    output n61122;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n29997, n57105;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire n49547, n57097, n2;
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    
    wire n57245, n2_adj_5259, n57244, n29994, n10, n57434, n30022, 
        n57446, n57965, n57551, n25962;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n56712, n52555, n25891, n57593, n6_c, n56700;
    wire [7:0]\data_in_frame[3]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29969, n29966, Kp_23__N_1080, n52308, n29963, n30019, 
        n29960, n29957, n29953, n29950, n29947, n29943, n29940, 
        n29937, n25976, n26324, n57972, n4_c, n3, n58033, n11, 
        n26069, n26336, n26496, Kp_23__N_993, n68623, n57482, n57914, 
        n35692, n57580, n2_adj_5260, n57243, n2_adj_5261, n57242, 
        n49548, n57104, n49546, n2_adj_5262, n57294, n2068, n30015;
    wire [23:0]n4762;
    
    wire n27767, n29933;
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    
    wire n58129, n57933, n25705, n57962, n25698, n1168;
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    
    wire n57918, n29930, n57688, n58024;
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    
    wire n62436, n2_adj_5263, n57241, n2_adj_5264;
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    
    wire n57113, n56714, n56706, n57691, n10_adj_5265, n52028, n52034, 
        n2_adj_5266, n57240, n2_adj_5267, n57239, n2_adj_5268, n57238, 
        n2_adj_5269, n57237, n2_adj_5270, n57236, n2_adj_5271, n57235, 
        n2_adj_5272, n57234, n2_adj_5273, n57233, n2_adj_5274, n57232, 
        n2_adj_5275, n57231, n2_adj_5276, n57230, n2_adj_5277, n57229, 
        n2_adj_5278, n57228, n2_adj_5279, n57227, n2_adj_5280, n57226, 
        n2_adj_5281;
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    
    wire n57225;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    
    wire n65574;
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    
    wire n63068, n63069, n63067, n69520, n69514, n14, n2_adj_5283, 
        n57224, n2_adj_5284, n57223, n2_adj_5285, n57222, n2_adj_5286, 
        n57221, n2_adj_5287, n57220, n2_adj_5288, n57219, n2_adj_5289, 
        n57218, n2_adj_5290;
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    
    wire n57217, n2_adj_5291, n57216, n2_adj_5292, n57215, n2_adj_5293, 
        n57214, n2_adj_5294, n57213, n2_adj_5295, n57212, n29926, 
        n2_adj_5296, n57211, n2_adj_5297, n57210, n65560, n69490, 
        n69562, n67258, n57103, n49545, n2_adj_5298;
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    
    wire n29076, n29923, n2_adj_5299, n57209, n2_adj_5300, n57208, 
        n2_adj_5301, n57207, n2_adj_5302, n57206, n29920, n56993;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n10_adj_5304, n57427;
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    
    wire \FRAME_MATCHER.i_31__N_2509 ;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5305, n2_adj_5306, n2_adj_5307, n29916, n29913;
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    
    wire n2_adj_5308, n2_adj_5309, n57205, n2_adj_5310, n2_adj_5311, 
        n2_adj_5312, n57204, n2_adj_5313, n25709, n62488, n62492, 
        n2_adj_5314, n57203, n2_adj_5315, n57202, n43390, n59293, 
        n2_adj_5316, n2_adj_5317, n57201, n30012, n29480, n2_adj_5318, 
        n2_adj_5319, n57200, n2_adj_5320, n30009, n57199, n57198, 
        n2_adj_5321, n29909, n57197, n57196, n57195, n29060, n29905, 
        n57194, n29726;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5322, n29901, n30006, n10_adj_5323, n6_adj_5324, \FRAME_MATCHER.i_31__N_2512 , 
        n26950, n29897, n57102, n49544, n29894, n57101, n49543;
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    
    wire n6_adj_5325, n26412, n3_adj_5326, \FRAME_MATCHER.i_31__N_2507 , 
        n65548, n65549, n65550, n65551, n57100, n49542, n23, n65552, 
        n65553, n65554, n27315, n28941, n33798, n65555, n5, n65556, 
        n65557, n65558, n52094, n6_adj_5327, n65563, n69655, n65570, 
        n29761;
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    
    wire n8_c, n57786, n3_adj_5328, n29768, n53193, n58136, n3_adj_5329, 
        n29771, n53044, n7_adj_5330;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n57870, n52022, n12, n29783, n29786, n29789, n29792, 
        n26253, n8_adj_5331, n3_adj_5332, n29880, n52986, n57867, 
        n3_adj_5333, n58074, n53003, n57522;
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    
    wire n24, n65571, n69649, n58086, n26138, n26899, n60087, 
        n22, n65572, n57845, n18, n68629, n26_c, n65581, n65582;
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    
    wire n53172, n57796, n6_adj_5334, n3_adj_5335, n65586, n58093, 
        n57467, n4_adj_5336, n51970;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    
    wire n59944, n12_adj_5337, n65592, n26539;
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    
    wire n65593;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    
    wire n53042, n53178, n16, n58083, n17, n65608, n65609, n58272, 
        n65615, n63023, n26545, n52143, n771, \FRAME_MATCHER.i_31__N_2508 , 
        n25545, n4_adj_5338, n62552, n57463, n3_adj_5339, n53077, 
        n57885, n65616, n65617, n65649, n3_adj_5340, n53159, n60167, 
        n59475, n53176, n10_adj_5341, n58049, n65660, n65661, Kp_23__N_748, 
        n52588, n26690, n14_adj_5342;
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    
    wire n2_adj_5343, n65662;
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    
    wire n2_adj_5344, n59292, n57741;
    wire [7:0]\data_out_frame[20]_c ;   // verilog/coms.v(100[12:26])
    
    wire n62504, n53137, n57812, n57805, n62510, n65663, n58090, 
        n62514, n62528, n62526, n57873, n62536, n62314, n65673, 
        n28404, n52492, n57905, n59473, n26373, n2_adj_5345, n58069, 
        n57734, n62540, n57789, n62320, n25835, n57902, n3_adj_5346, 
        n57099, tx_transmit_N_3416, n52026, n52132, n53119, n3_adj_5347, 
        n53207, n3_adj_5348, n2_adj_5349, n53107, n6_adj_5350, n3_adj_5351, 
        n2_adj_5352, n57981, n10_adj_5353, n2_adj_5354, n53093, n3_adj_5355, 
        n2_adj_5356, n2_adj_5357, n52390, n2_adj_5358, n2217, n52188, 
        n23735, n16_adj_5359, n28421, n2_adj_5360, n53209, n52516, 
        n57799, n52042, n17_adj_5361, n29828, n6_adj_5362, n52984, 
        n57839, n51944, n57876, n10_adj_5363, n52973, n51995, n10_adj_5364, 
        n25162, n59919, n40928, n7_adj_5365, n57722, n57856, n2_adj_5366, 
        n57193, n2_adj_5367, n57192, n2_adj_5368, n57191, n2_adj_5369, 
        n57190;
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    
    wire n57747, n62546, n29806, n2_adj_5370, n57189, n57531, n25734, 
        n57750, n52663, n2_adj_5371, n57188, n2_adj_5372, n57187, 
        n2_adj_5373, n57186, n2_adj_5374, n57114, n1720, n56594, 
        n2_adj_5375, n57115, n2_adj_5376, n57116, n2_adj_5377, n57117, 
        n52068, n58111, n52024, n14_adj_5378, n10_adj_5379, n58123, 
        n57709, n26731, n26432, n1699, n57470, n2_adj_5380, n57118, 
        n59803, n2_adj_5381, n57119, n57599, n2_adj_5382, n57121, 
        n2_adj_5383, n57122, n62384, n2_adj_5384, n57123, n2_adj_5385, 
        n57124, n2_adj_5386, n57125, n62386, n2076, n62394, n26664, 
        n62398, n2_adj_5387, n57126, n57455, n52198, n26279, n62404, 
        n58080, n62410, n2_adj_5388, n57127, n62562, n2_adj_5389, 
        n57128, n2_adj_5390, n57129, n57744, n57608, n62416, n51946, 
        n26896, n62566, n60272, n60035, n23733, n57782, n58056, 
        n60044, n30002, n2_adj_5391, n57130, n2_adj_5392, n57131, 
        n2_adj_5393, n57111, n2_adj_5394, n57132, n2_adj_5395, n57133, 
        n2_adj_5396, n57134, n52175, n2_adj_5397, n57135, n4_adj_5398, 
        n57571, n62322, n2_adj_5399, n57136, n2_adj_5400, n57137, 
        n2_adj_5401, n57138, n28439, n2_adj_5402, n57139, n57848, 
        n6_adj_5403, n53027, n2_adj_5405, n57140, n52236, n62376, 
        n69643, n63029, n29720, n58030, n6_adj_5406, n57953;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n69631, n36, n58008, n6_adj_5407, n29719, n57622, n26291, 
        n57604, n52107, n57936, n57516, n52684, n8_adj_5408, n60454, 
        n51960, n6_adj_5409, n57641, n57996, n57644, n69634, n52338, 
        n26623, n57833, n29679;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n29665, n2_adj_5410, n57141, n8_adj_5411, n52991, n12_adj_5412, 
        n25990, n58021, n2_adj_5414, n57142, n2_adj_5415, n57143, 
        n2_adj_5416, n57144, n2_adj_5417, n29019, n2_adj_5418, n57145, 
        n3_adj_5419, n2_adj_5420, n29017, n2_adj_5421, n57146, n2_adj_5422, 
        n57147, n2_adj_5423, n57148, n2_adj_5424, n57149, n2_adj_5425, 
        n57150, n2_adj_5426, n29011, n2_adj_5427, n57151, n2_adj_5428, 
        n57152, n53102, n57541, n24_adj_5429, n2_adj_5430, n57153, 
        n57615, n2_adj_5431, n57154, n2_adj_5432, n57155, n2_adj_5433, 
        n57156, n2_adj_5434, n57157, n2_adj_5435, n57158, n2_adj_5436, 
        n57159, n2_adj_5437, n57160, n2_adj_5438, n57161, n2_adj_5439, 
        n57162, n26795, n2_adj_5440, n58042, n12_adj_5441, n2_adj_5442, 
        n2_adj_5443, n28080, n2_adj_5444, n57163, n2_adj_5445, n57164, 
        n57165, n57166, n28082, n28084, n28086, n28088, n28090, 
        n28092, n28094, n28096, n28098, n28100, n28102, n28104, 
        n28106, n28108, n28110, n28112, n28114, n28116, n28118, 
        n28120, n28122, n28124, n28126, n28128, n28130, n28132, 
        n28134, n28136, n28138, n28140, n28142, n57167, n57476, 
        n6_adj_5446, n26380, n57939, n57950, n14_adj_5447, n58126, 
        n25702, n58017, n15_c, n57534, n26645, n4_adj_5448, n57452, 
        n57921, n60077, n57293, n57292, n57291, n57290, n58108, 
        n57289, n57288, n57287, n1516, n57574, n52635, n52209, 
        n57286;
    wire [31:0]n133;
    
    wire n50838, n50837, n57285, n50836, n57284, n50835, n50834, 
        n50833, n50832, n50831, n50830, n50829, n50828, n50827, 
        n50826, n50825, n50824, n50823, n6_adj_5449, n50822, n50821, 
        n50820, n50819, n50818, n50817, n50816, n50815, n50814, 
        n50813, n50812, n50811, n50810, n50809, n50808, n29483, 
        n29486, n29489, n29492, n29495, n29498, n56504, n26282, 
        n53133, n26104, n60324, n30466, n29504, n30414, n30413, 
        n30412, n30411, n30410, n30409, n30408, n30407;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n30406, n30405, n30404, n53199, n62454, n30403, n30402, 
        n30401, n30400, n30399;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n30398, n2_adj_5450, n57283, n30397, n30396, n30395, n30394, 
        n30393, n30392, n30391;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n30390, n62456, n30389, n62424, n30388;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n43569, \FRAME_MATCHER.i_31__N_2511 , n1, n30387, n62458, 
        n30386, n30385, n30384, n2_adj_5451, n57282, n30370, n57577, 
        n58036, n62472, n2_adj_5452, n57281, n30025, n30028, n30031, 
        n30034, n30037, n30040, n30043, n30046;
    wire [7:0]\data_in_frame[6]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30049, n56514;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n56520, n56518, n2_adj_5453, n57280, n62466, n1130, n62474, 
        n62476, n30128;
    wire [7:0]\data_in_frame[10]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58002, n57558, n57968, n62430, n30206, n30209, n30213, 
        n30216, n30219, n30223, n30226, n62482, n30260, n26461, 
        n26844, n56554;
    wire [7:0]\data_in_frame[19]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30229, n30222, n62300, n26553, n57908, n29638, n29641, 
        n29646, n29649, n29657, n29666, n2_adj_5456, n57279, n2_adj_5457, 
        n57278, n2_adj_5458, n57277, n2_adj_5459, n57276, n2_adj_5460, 
        n57275, n29680, n57590, n57496, n10_adj_5461, n29529, n2_adj_5462, 
        n57274, n58105, n10_adj_5463, n2_adj_5464, n57273, n51958, 
        n57999, n6_adj_5465, n52036, n57672, n53030, n2_adj_5466, 
        n57272, n51954, n57525, n57706, n26738, n57816, n53052, 
        n58061, n58120, n69866, n27046, n2048, n2049, n20442, 
        n56292, n2060, n27049, \FRAME_MATCHER.i_31__N_2514 , n2_adj_5467, 
        n57271, n57700, n25808, n59240, Kp_23__N_1551, n2_adj_5468, 
        n57270, n57502, n57942, n10_adj_5469, n2_adj_5470, n57269, 
        n57681, n2_adj_5471, n57268, n2_adj_5472, n57267, n2_adj_5473, 
        n57266, n25937, n2_adj_5475, n57265, n2_adj_5476, n57264, 
        n57764, n57634, n2_adj_5477, n57263, n52141, n2_adj_5478, 
        n57262, n59871, n57984, n2_adj_5479, n57261, n29684, n2_adj_5480, 
        n57260, n2_adj_5481, n57259, n2_adj_5482, n57258, n2_adj_5483, 
        n57257, n2_adj_5484, n57256, n2_adj_5485, n57255, n20, n22_adj_5486, 
        n30_c, n28, n57564, n34_adj_5487, n32_c, n36_adj_5488, n23_adj_5489, 
        n57792, n52449, n14_adj_5490, n10_adj_5491, n52147, n25207, 
        n57587, n20_adj_5492, n52995, n19_c, n58141, n57492, n57761, 
        n21_c, n58039, n26009, n26025, n6_adj_5493, n59287, n25751, 
        n57547, n6_adj_5494, n51948, n57675, n58011, n12_adj_5495, 
        n26121, n57612, n57896, n1563, n58045, n57756, n6_adj_5496, 
        n52413, n26061, n4_adj_5497, n57458, n9, n8_adj_5498, n57975, 
        n2_adj_5499, n57168, n58114, n15_adj_5500, n2_adj_5501, n57169, 
        n57859, n14_adj_5502, n59679, n25858, n6_adj_5503, n57663, 
        n26367, n58005, n10_adj_5504, n57479, n57930, n2_adj_5505, 
        n57170, n58077, n57697, n22_adj_5506, n57842, n57631, n57719, 
        n24_adj_5507, n57822, n57513, n58144, n23_adj_5508, n25_adj_5509, 
        n57927, n10_adj_5510, n51992, n8_adj_5511, n53059, n57473, 
        n52693, n57519, n25906, n22_adj_5512, n2_adj_5513, n57171, 
        n57555, n57767, n15_adj_5514, n24_adj_5515, n20_adj_5516, 
        n68627, Kp_23__N_974, n26715, n2_adj_5517, n57172, n6_adj_5518, 
        n2_adj_5519, n57173, n58053, n6_adj_5520, n14_adj_5521, n2_adj_5522, 
        n57174, n26818, n2_adj_5523, n57175, n2_adj_5524, n57176, 
        n9_adj_5525, n58072, n26487, n57443, n59598, n59447, n2_adj_5526, 
        n57177, n14_adj_5527, n53022, n9_adj_5528, n57830, n57628, 
        n25266, n2_adj_5529, n57178, n2_adj_5530, n57112, n2_adj_5531, 
        n57120, n2_adj_5532, n57179, n2_adj_5533, n57180, n2_adj_5534, 
        n57181, n2_adj_5535, n57254, n26721, n57538, n2_adj_5536, 
        n57253, n2_adj_5537, n57252, n57899, n4_adj_5538, n57461, 
        n57924, n2_adj_5539, n57251, n2_adj_5540, n57182, n25927, 
        n12_adj_5541, n15_adj_5542, n14_adj_5543, n2_adj_5544, n57183, 
        n62334, n2_adj_5545, n57184, n2_adj_5546, n57185, n2_adj_5547, 
        n57110, n3_adj_5548, n57303, n57304, n57305, n57301, n57306, 
        n57299, n3_adj_5549, n57307, n57308, n57309, n57310, n57311, 
        n57302, n57312, n57300, n57298, n62342, n28942, n57313, 
        n1_adj_5550, n1_adj_5551, n1_adj_5552, n1_adj_5553, n1_adj_5554, 
        n1_adj_5555, n1_adj_5556, n57098, n28931, n58102, n62344, 
        n57250, n62352, n62356, n1_adj_5557, n58027, n25784, n52173, 
        n26931, n62362, n62368, n57249, n57568, n57248, n57528, 
        n57891, n62292, n62298, n57893, n57247, n57246, n58099, 
        n10_adj_5558, n26853, n57852, n57731, n25769, n10_adj_5559, 
        n6_adj_5560, n12_adj_5561, n25941, n1655, Kp_23__N_760, n57506, 
        n57959, n22_adj_5562, Kp_23__N_772, n21_adj_5563, n14_adj_5564, 
        n23_adj_5565, n57666, n57561, n26_adj_5566, n19_adj_5567, 
        n58014, n16_adj_5568, n57619, n57669, n24_adj_5569, n57678, 
        n28_adj_5570, Kp_23__N_799, n57648, n26428, n57694, n58028, 
        n10_adj_5571, n52130, n26310, n6_adj_5572, n6_adj_5573, n57725, 
        n69619, n6_adj_5574, n26231, n24009, n69622, n69613, n69616, 
        n8_adj_5575, n10_adj_5576, n14_adj_5577, n10_adj_5578, n12_adj_5579, 
        n26370, n60278, n26401, n57596, Kp_23__N_872, n26508, n13, 
        n25953, n6_adj_5580, Kp_23__N_869, n59349, n62656, n20_adj_5581, 
        n18_adj_5582, n19_adj_5583, n57752, n17_adj_5584, n52194, 
        n26304, n15_adj_5586, n14_adj_5587, n24005, n6_adj_5588, n25842, 
        n25745, n57911, n52001, n7_adj_5589, n63059, n28205, n63060, 
        n63058, n69607, n6_adj_5590, n57809, n10_adj_5591, n22911, 
        n62676, n8_adj_5592, n52504, n53032, n69610, n69568, n67824, 
        n8_adj_5593, n28147, n63050, n59453, n60320, n70027, n12_adj_5594, 
        n63051, n10_adj_5595, n60373, n63049, n59724, n62682, n24_adj_5596, 
        n62684, n23_adj_5597, n8_adj_5598, n60421, n63142, n59645, 
        n63143, n63140, n63139, n19_adj_5599, n63013, n22_adj_5600, 
        n62686, n32_adj_5601, n27_c, n63014, n63017, n63016, n63151, 
        n63152, n62996, n62995, n63127, n63128, n63002, n63001, 
        n65734, n28145, n63044, n63045, n63043, n65735, n63115, 
        n1954, n1951, n1957, n59892, n63116, n63065, n63064, n25621, 
        n5_adj_5602, n15_adj_5603, n14_adj_5604, n59699, n28155, n62814, 
        Kp_23__N_878, n63074, n62844, n28_adj_5605, n63075, n63073, 
        n69538, n69526, n67267, n69556, n62812, n69502, n69550, 
        n67419, n69544, n69532, n65732, n27_adj_5606, n63022, n1_adj_5607, 
        n63028, n63163, n63164, n63005, n59374, n4452, n20437, 
        n22769, n63004, n3303, n63010, n63011, n63020, n63019, 
        n62601, n60102, n1955, n63053, n63054, n63052, n25468, 
        n65787, n27626, n59773, n25550, n63118, n57396, n10_adj_5609, 
        n57728, n63119, n14_adj_5610, n25618, n63038, n20_adj_5611, 
        n63037, n63121, n25492, n19_adj_5612, n62802, n63122, n25676, 
        n18_adj_5613, n63026, n25572, n20_adj_5614, n15_adj_5615, 
        n63025, n33795, n62917, n10_adj_5616, n62918, n14_adj_5617, 
        n63173, n15_adj_5618, n63172, n16_adj_5619, n17_adj_5620, 
        n60447, n12_adj_5622, n44, n42, n42760, n6_adj_5623, n43_adj_5624, 
        n41, n40, n39, n50, n45_adj_5625, n57399, n106, n40952, 
        n145, n40997, n51920, n4_adj_5629, n4_adj_5630, n57430, 
        n5_adj_5631, n107, n65697, n62738, n40982, n69841, n63105, 
        n69835, n63111, n65728, n69595, n69598, n69589, n69829, 
        n63114, n41131, n69592, n69583, n69586, n69823, n63126, 
        n69466, n69817, n69580, n7_adj_5635, n69577, n69571, n69574, 
        n69565, n40967, n12_adj_5636, n10_adj_5637, n11_adj_5638, 
        n9_adj_5639, n57651, n69559, n57638, n62674, n18_adj_5640, 
        n20_adj_5641, n60517, n12_adj_5642, n69553, n69547, n69805, 
        n69541, n69535, n69472, n69799, n7_adj_5643, n69529, n69523, 
        n69517, n69511, n69499, n69478, n69793, n7_adj_5644, n7_adj_5647, 
        n69487, n69484, n69787, n69481, n7_adj_5648, n69475, n69469, 
        n69463, n69781;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n58925, n29, n23_adj_5650;
    wire [24:0]o_Rx_DV_N_3488;
    
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n56422));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29997));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1099_8_lut (.I0(n57097), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n49547), .O(n57105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_8_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2), .S(n57245));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5259), .S(n57244));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29994));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15946_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n30022));
    defparam i15946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[3] [5]), .I1(n57446), .I2(n57965), 
            .I3(n57551), .O(n25962));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i52891_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[0] [6]), .I2(n7), 
            .I3(GND_net), .O(n56712));   // verilog/coms.v(94[13:20])
    defparam i52891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[9] [0]), .I1(n52555), .I2(n25891), 
            .I3(n57593), .O(n6_c));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29989));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29986));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29983));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n56418));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29979));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3]_c [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n56700));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n56414));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29966));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[9] [0]), .I1(n52555), .I2(n25891), 
            .I3(Kp_23__N_1080), .O(n52308));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i29 (.Q(\data_in_frame[3][4] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29963));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15943_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n30019));
    defparam i15943_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29957));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0][1] ), .C(clk16MHz), 
           .D(n29701));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i26 (.Q(\data_in_frame[3][1] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29953));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29950));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29947));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n56410));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29943));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29940));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29937));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n25891), .I1(n25976), .I2(\data_in_frame[10] [6]), 
            .I3(GND_net), .O(n58117));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1103 (.I0(n25891), .I1(n25976), .I2(n26324), 
            .I3(GND_net), .O(n57972));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_3_lut (.I0(n4_c), .I1(n3), .I2(n58033), .I3(GND_net), 
            .O(n11));   // verilog/coms.v(77[16:43])
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1104 (.I0(n4_c), .I1(n3), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n26069));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1105 (.I0(n26336), .I1(n26496), .I2(Kp_23__N_993), 
            .I3(n68623), .O(n58033));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1105.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1106 (.I0(n26336), .I1(n26496), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n57482));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1106.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1107 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(n57914), .O(n35692));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1108 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[0][7] ), .I3(GND_net), .O(n57580));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_adj_1108.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5260), .S(n57243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5261), .S(n57242));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_8 (.CI(n49547), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n49548));
    SB_LUT4 add_1099_7_lut (.I0(n57097), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n49546), .O(n57104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_7_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5262), .S(n57294));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2068), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i15939_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n30015));
    defparam i15939_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n56406));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27767), 
            .D(n4762[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29933));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1109 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[5] [5]), .I3(n58129), .O(n57933));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1110 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n25705));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1110.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(n57962), .I3(n25698), .O(n1168));   // verilog/coms.v(74[16:27])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1111 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[10] [5]), .I3(\data_out_frame[8] [4]), .O(n57918));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29930));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_7 (.CI(n49546), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n49547));
    SB_LUT4 i1_3_lut_4_lut_adj_1112 (.I0(n57688), .I1(n58024), .I2(\data_out_frame[16] [6]), 
            .I3(\data_out_frame[16] [4]), .O(n62436));   // verilog/coms.v(88[17:28])
    defparam i1_3_lut_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5263), .S(n57241));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n56402));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5264), .S(n57113));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i52892_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[0] [5]), .I2(n7), 
            .I3(GND_net), .O(n56714));   // verilog/coms.v(94[13:20])
    defparam i52892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52890_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[0] [4]), .I2(n7), 
            .I3(GND_net), .O(n56706));   // verilog/coms.v(94[13:20])
    defparam i52890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1113 (.I0(n57691), .I1(n10_adj_5265), .I2(\data_in_frame[8] [2]), 
            .I3(n52028), .O(n52034));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5266), .S(n57240));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5267), .S(n57239));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5268), .S(n57238));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5269), .S(n57237));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5270), .S(n57236));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5271), .S(n57235));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5272), .S(n57234));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5273), .S(n57233));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5274), .S(n57232));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5275), .S(n57231));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5276), .S(n57230));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5277), .S(n57229));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5278), .S(n57228));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5279), .S(n57227));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5280), .S(n57226));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5281), .S(n57225));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1114 (.I0(n57691), .I1(n10_adj_5265), .I2(\data_in_frame[8] [2]), 
            .I3(\data_in_frame[12] [5]), .O(n57657));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i50085_2_lut (.I0(\data_out_frame[0] [2]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65574));
    defparam i50085_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i47340_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63068));
    defparam i47340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47341_4_lut (.I0(n63068), .I1(n65574), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[1] ), .O(n63069));
    defparam i47341_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i47339_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63067));
    defparam i47339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1115 (.I0(n57691), .I1(n10_adj_5265), .I2(\data_in_frame[8] [2]), 
            .I3(\data_in_frame[14] [5]), .O(n6));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i29880110_i1_3_lut (.I0(n69520), .I1(n69514), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14));
    defparam i29880110_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5283), .S(n57224));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5284), .S(n57223));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5285), .S(n57222));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5286), .S(n57221));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5287), .S(n57220));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5288), .S(n57219));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5289), .S(n57218));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5290), .S(n57217));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5291), .S(n57216));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5292), .S(n57215));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5293), .S(n57214));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5294), .S(n57213));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5295), .S(n57212));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5296), .S(n57211));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5297), .S(n57210));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50099_2_lut (.I0(n69640), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65560));
    defparam i50099_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51530_3_lut (.I0(n69490), .I1(n69562), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n67258));
    defparam i51530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1099_6_lut (.I0(n57097), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n49545), .O(n57103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_6_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5298), .S(n29076));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29923));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_6 (.CI(n49545), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n49546));
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5299), .S(n57209));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5300), .S(n57208));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5301), .S(n57207));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5302), .S(n57206));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29920));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i23269_3_lut (.I0(n43), .I1(n379), .I2(n405), .I3(GND_net), 
            .O(n4));
    defparam i23269_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i3_4_lut (.I0(n56993), .I1(\FRAME_MATCHER.i [2]), .I2(n10_adj_5304), 
            .I3(\FRAME_MATCHER.i [0]), .O(n57427));
    defparam i3_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 select_777_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5305));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29714));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5306));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5307));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29916));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29913));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5309), .S(n57205));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23281_3_lut (.I0(n379), .I1(n459), .I2(n11610), .I3(GND_net), 
            .O(n37308));
    defparam i23281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5312), .S(n57204));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1116 (.I0(n25709), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[8] [2]), .I3(n62488), .O(n62492));
    defparam i1_3_lut_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5314), .S(n57203));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5315), .S(n57202));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n43390), .I2(\FRAME_MATCHER.i [1]), 
            .I3(GND_net), .O(n59293));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_777_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5317), .S(n57201));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15936_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n30012));
    defparam i15936_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15404_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n57425), .I3(GND_net), .O(n29480));   // verilog/coms.v(130[12] 305[6])
    defparam i15404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 select_777_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5319), .S(n57200));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15933_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n30009));
    defparam i15933_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5316), .S(n57199));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5313), .S(n57198));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5311), .S(n57197));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5310), .S(n57196));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5315));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5308), .S(n57195));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5314));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n56398));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5306), .S(n29060));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5305), .S(n57194));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5309));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29726));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29901));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15930_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n30006));
    defparam i15930_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5302));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5299));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1117 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_5323));   // verilog/coms.v(157[7:23])
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1118 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5324), .I3(\FRAME_MATCHER.i_31__N_2512 ), .O(n26950));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1118.LUT_INIT = 16'haaa8;
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29897));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1099_5_lut (.I0(n57097), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n49544), .O(n57102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1119 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [0]), 
            .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5298));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1119.LUT_INIT = 16'ha088;
    SB_CARRY add_1099_5 (.CI(n49544), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n49545));
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29894));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1099_4_lut (.I0(n57097), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n49543), .O(n57101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1099_4 (.CI(n49543), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n49544));
    SB_LUT4 select_777_Select_223_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n6_adj_5325), .I3(n26412), 
            .O(n3_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i50097_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65548));   // verilog/coms.v(158[12:15])
    defparam i50097_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50071_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65549));   // verilog/coms.v(158[12:15])
    defparam i50071_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50072_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65550));   // verilog/coms.v(158[12:15])
    defparam i50072_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50073_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65551));   // verilog/coms.v(158[12:15])
    defparam i50073_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_1099_3_lut (.I0(n57097), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n49542), .O(n57100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_3_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0][2] ), .C(clk16MHz), 
           .D(n29739));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut (.I0(LED_c), .I1(n33801), .I2(GND_net), .I3(GND_net), 
            .O(n23));   // verilog/TinyFPGA_B.v(4[10:13])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50074_2_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65552));   // verilog/coms.v(158[12:15])
    defparam i50074_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50075_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65553));   // verilog/coms.v(158[12:15])
    defparam i50075_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50076_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65554));   // verilog/coms.v(158[12:15])
    defparam i50076_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14865_4_lut (.I0(n2873), .I1(n23), .I2(n27315), .I3(\FRAME_MATCHER.i_31__N_2513 ), 
            .O(n28941));   // verilog/coms.v(130[12] 305[6])
    defparam i14865_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i19722_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n33798));   // verilog/coms.v(118[11:12])
    defparam i19722_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i50077_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65555));   // verilog/coms.v(158[12:15])
    defparam i50077_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(n33798), .I1(n27726), .I2(GND_net), 
            .I3(GND_net), .O(n5));
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'heeee;
    SB_LUT4 i50078_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65556));   // verilog/coms.v(158[12:15])
    defparam i50078_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50079_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65557));   // verilog/coms.v(158[12:15])
    defparam i50079_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50080_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65558));   // verilog/coms.v(158[12:15])
    defparam i50080_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[13] [7]), .I3(n52094), .O(n6_adj_5327));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i50562_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65563));   // verilog/coms.v(158[12:15])
    defparam i50562_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53994 (.I0(byte_transmit_counter[3]), 
            .I1(n67258), .I2(n65560), .I3(byte_transmit_counter[4]), .O(n69655));
    defparam byte_transmit_counter_3__bdd_4_lut_53994.LUT_INIT = 16'he4aa;
    SB_LUT4 i50688_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65570));   // verilog/coms.v(158[12:15])
    defparam i50688_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29761));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0][3] ), .C(clk16MHz), 
           .D(n29764));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_222_i3_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n8_c), .I3(n57786), .O(n3_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n29768));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_221_i3_4_lut (.I0(n53193), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n58136), .I3(\data_out_frame[25] [4]), .O(n3_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_221_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29771));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_out_frame[25] [3]), .I1(n53044), 
            .I2(GND_net), .I3(GND_net), .O(n53193));
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 n69655_bdd_4_lut (.I0(n69655), .I1(n14), .I2(n7_adj_5330), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n69655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n56706));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n56714));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[20] [7]), .I1(n57870), .I2(n53193), 
            .I3(n52022), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29783));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29786));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n29789));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29792));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n56712));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0][7] ), .C(clk16MHz), 
           .D(n29802));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_220_i3_4_lut (.I0(n26253), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n12), .I3(n8_adj_5331), .O(n3_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29880), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29879), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29878), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29877), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_219_i3_3_lut (.I0(n52986), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n57867), .I3(GND_net), .O(n3_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_219_i3_3_lut.LUT_INIT = 16'h4848;
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29876), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29875), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i10_4_lut (.I0(n58074), .I1(n53003), .I2(n57522), .I3(\data_out_frame[18] [5]), 
            .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i50086_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65571));   // verilog/coms.v(158[12:15])
    defparam i50086_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29874), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29873), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29872), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29871), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29870), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29869), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29868), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29867), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29866), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29865), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29864), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29863), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29862), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29861), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54014 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[6] [4]), .I2(\data_out_frame[7] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n69649));
    defparam byte_transmit_counter_0__bdd_4_lut_54014.LUT_INIT = 16'he4aa;
    SB_LUT4 i8_4_lut (.I0(n58086), .I1(n26138), .I2(n26899), .I3(n60087), 
            .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i50087_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65572));   // verilog/coms.v(158[12:15])
    defparam i50087_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut (.I0(n57845), .I1(n24), .I2(n18), .I3(n68629), 
            .O(n26_c));
    defparam i12_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i50107_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65581));   // verilog/coms.v(158[12:15])
    defparam i50107_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29860), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50108_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65582));   // verilog/coms.v(158[12:15])
    defparam i50108_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[17] [0]), .I1(n26_c), .I2(n22), 
            .I3(n53172), .O(n52022));
    defparam i13_4_lut.LUT_INIT = 16'h9669;
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29859), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29858), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut (.I0(n57796), .I1(\data_out_frame[25] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5334));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_218_i3_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n6_adj_5334), .I3(n52022), 
            .O(n3_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29857), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29856), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29855), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29854), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50141_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65586));   // verilog/coms.v(158[12:15])
    defparam i50141_2_lut.LUT_INIT = 16'h2222;
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29853), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1122 (.I0(n53095), .I1(n58093), .I2(GND_net), 
            .I3(GND_net), .O(n58074));
    defparam i1_2_lut_adj_1122.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(n57467), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5336));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(n51970), .I1(\data_out_frame[16] [4]), .I2(n52011), 
            .I3(n4_adj_5336), .O(n57870));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1124 (.I0(\data_out_frame[22] [5]), .I1(n57870), 
            .I2(\data_out_frame[23] [1]), .I3(n59944), .O(n12_adj_5337));
    defparam i5_4_lut_adj_1124.LUT_INIT = 16'h9669;
    SB_LUT4 i50251_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65592));   // verilog/coms.v(158[12:15])
    defparam i50251_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut (.I0(n26539), .I1(n12_adj_5337), .I2(n58086), .I3(\data_out_frame[24] [7]), 
            .O(n52986));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29852), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50166_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65593));   // verilog/coms.v(158[12:15])
    defparam i50166_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1125 (.I0(\data_out_frame[21] [1]), .I1(n53042), 
            .I2(n58074), .I3(n53178), .O(n16));
    defparam i6_4_lut_adj_1125.LUT_INIT = 16'h9669;
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29851), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut (.I0(\data_out_frame[23] [2]), .I1(n57836), .I2(n58083), 
            .I3(\data_out_frame[18][3] ), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_out_frame[16] [1]), .I2(n16), 
            .I3(\data_out_frame[23] [1]), .O(n53044));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i50207_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65608));   // verilog/coms.v(158[12:15])
    defparam i50207_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50225_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65609));   // verilog/coms.v(158[12:15])
    defparam i50225_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i42588_2_lut_3_lut (.I0(n3470), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n58272));
    defparam i42588_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i50232_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65615));   // verilog/coms.v(158[12:15])
    defparam i50232_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n69649_bdd_4_lut (.I0(n69649), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n63023));
    defparam n69649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(n26545), .I1(\data_out_frame[23][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n52143));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1127 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25545), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n4_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1127.LUT_INIT = 16'hfff4;
    SB_LUT4 i1_3_lut (.I0(n58136), .I1(n53044), .I2(n52986), .I3(GND_net), 
            .O(n62552));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 select_777_Select_217_i3_4_lut (.I0(n52143), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n57463), .I3(n62552), .O(n3_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i3_4_lut_adj_1128 (.I0(\data_out_frame[24] [6]), .I1(n53077), 
            .I2(\data_out_frame[25] [0]), .I3(n57885), .O(n57796));
    defparam i3_4_lut_adj_1128.LUT_INIT = 16'h9669;
    SB_LUT4 i50236_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65616));   // verilog/coms.v(158[12:15])
    defparam i50236_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50235_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65617));   // verilog/coms.v(158[12:15])
    defparam i50235_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50367_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65649));   // verilog/coms.v(158[12:15])
    defparam i50367_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_777_Select_216_i3_3_lut (.I0(n57463), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n57796), .I3(GND_net), .O(n3_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_216_i3_3_lut.LUT_INIT = 16'h8484;
    SB_LUT4 i3_4_lut_adj_1129 (.I0(n53159), .I1(\data_out_frame[16][3] ), 
            .I2(n60167), .I3(\data_out_frame[14] [3]), .O(n57467));
    defparam i3_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut (.I0(n59475), .I1(\data_out_frame[20] [7]), .I2(n53176), 
            .I3(n57467), .O(n10_adj_5341));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29850), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut (.I0(n53095), .I1(n10_adj_5341), .I2(\data_out_frame[21] [1]), 
            .I3(GND_net), .O(n26545));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29849), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n58049));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i50310_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65660));   // verilog/coms.v(158[12:15])
    defparam i50310_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26253));
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29848), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29847), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n57867));
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29846), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50311_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65661));   // verilog/coms.v(158[12:15])
    defparam i50311_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29845), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29844), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57786));
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29843), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1134 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0][0] ), 
            .I2(Kp_23__N_748), .I3(GND_net), .O(n52588));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut (.I0(n26690), .I1(\data_in_frame[1] [0]), .I2(\data_in_frame[0][7] ), 
            .I3(\data_in_frame[0] [6]), .O(n14_adj_5342));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h4114;
    SB_LUT4 select_777_Select_25_i2_3_lut (.I0(\data_out_frame[3] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_adj_1135 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[22] [6]), 
            .I2(\data_out_frame[22] [7]), .I3(GND_net), .O(n58086));
    defparam i2_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 i50312_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65662));   // verilog/coms.v(158[12:15])
    defparam i50312_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1136 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n26690));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_15_i2_3_lut (.I0(\data_out_frame[1] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1137 (.I0(n59292), .I1(n57741), .I2(n58086), 
            .I3(\data_out_frame[20]_c [1]), .O(n62504));
    defparam i1_4_lut_adj_1137.LUT_INIT = 16'h9669;
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29842), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_3 (.CI(n49542), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n49543));
    SB_LUT4 i1_4_lut_adj_1138 (.I0(n53137), .I1(n57812), .I2(n57805), 
            .I3(n62504), .O(n62510));
    defparam i1_4_lut_adj_1138.LUT_INIT = 16'h9669;
    SB_LUT4 i50313_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65663));   // verilog/coms.v(158[12:15])
    defparam i50313_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1139 (.I0(n58090), .I1(n62510), .I2(n52011), 
            .I3(GND_net), .O(n62514));
    defparam i1_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1140 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[23] [5]), 
            .I2(\data_out_frame[24] [7]), .I3(\data_out_frame[24] [5]), 
            .O(n62528));
    defparam i1_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1141 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[24] [1]), 
            .I2(\data_out_frame[23] [7]), .I3(GND_net), .O(n62526));
    defparam i1_3_lut_adj_1141.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1142 (.I0(n57873), .I1(n62526), .I2(n58049), 
            .I3(n62528), .O(n62536));
    defparam i1_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1143 (.I0(n57786), .I1(n57867), .I2(\data_out_frame[25] [6]), 
            .I3(\data_out_frame[25] [3]), .O(n62314));
    defparam i1_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i50345_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65673));   // verilog/coms.v(158[12:15])
    defparam i50345_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14329_1_lut (.I0(n3470), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28404));   // verilog/coms.v(148[4] 304[11])
    defparam i14329_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1144 (.I0(n52492), .I1(n57905), .I2(n26545), 
            .I3(n62514), .O(n59473));
    defparam i1_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1145 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0][2] ), 
            .I2(\data_in_frame[0][1] ), .I3(GND_net), .O(n26373));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1145.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_14_i2_3_lut (.I0(\data_out_frame[1] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29841), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1146 (.I0(n58069), .I1(n62536), .I2(n26253), 
            .I3(n57734), .O(n62540));
    defparam i1_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1147 (.I0(n57789), .I1(n26412), .I2(n53077), 
            .I3(n62314), .O(n62320));
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1148 (.I0(n62320), .I1(n62540), .I2(n59473), 
            .I3(n53077), .O(n57463));
    defparam i1_4_lut_adj_1148.LUT_INIT = 16'h9669;
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29840), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29839), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1149 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0][3] ), .I3(GND_net), .O(n25835));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_215_i3_4_lut (.I0(n57902), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n57463), .I3(\data_out_frame[25] [0]), .O(n3_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29838), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29837), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29836), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29835), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1099_2_lut (.I0(n57097), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n57099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_out_frame[24] [4]), .I1(n52026), 
            .I2(GND_net), .I3(GND_net), .O(n52132));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_213_i3_4_lut (.I0(n53119), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\data_out_frame[24] [3]), .I3(n52132), .O(n3_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_213_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29834), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n57734));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29833), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_212_i3_4_lut (.I0(n53119), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n57734), .I3(n53207), .O(n3_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_212_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_777_Select_13_i2_3_lut (.I0(\data_out_frame[1] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_2_lut_adj_1152 (.I0(n53107), .I1(\data_out_frame[24][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5350));
    defparam i2_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_211_i3_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n6_adj_5350), .I3(n53207), 
            .O(n3_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_211_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29832), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_11_i2_3_lut (.I0(\data_out_frame[1] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i4_4_lut_adj_1153 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[24] [0]), 
            .I2(\data_out_frame[24] [1]), .I3(n57981), .O(n10_adj_5353));
    defparam i4_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_9_i2_3_lut (.I0(\data_out_frame[1] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_777_Select_210_i3_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n10_adj_5353), .I3(n53093), 
            .O(n3_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_777_Select_8_i2_3_lut (.I0(\data_out_frame[1] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_777_Select_4_i2_3_lut (.I0(\data_out_frame[0] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29831), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29830), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1154 (.I0(n52390), .I1(n53093), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n26412));
    defparam i2_3_lut_adj_1154.LUT_INIT = 16'h6969;
    SB_LUT4 select_777_Select_3_i2_3_lut (.I0(\data_out_frame[0] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i6_4_lut_adj_1155 (.I0(n2217), .I1(n52188), .I2(n57741), .I3(n23735), 
            .O(n16_adj_5359));
    defparam i6_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(n3470), .I1(n10_adj_5323), .I2(n59293), 
            .I3(GND_net), .O(n28421));
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 select_777_Select_2_i2_3_lut (.I0(\data_out_frame[0] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i7_4_lut_adj_1156 (.I0(n53209), .I1(n52516), .I2(n57799), 
            .I3(n52042), .O(n17_adj_5361));
    defparam i7_4_lut_adj_1156.LUT_INIT = 16'h9669;
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29829), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1157 (.I0(n17_adj_5361), .I1(n53172), .I2(n16_adj_5359), 
            .I3(n53137), .O(n53207));
    defparam i9_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1158 (.I0(n3470), .I1(n10_adj_5323), 
            .I2(rx_data_ready), .I3(\FRAME_MATCHER.rx_data_ready_prev ), 
            .O(n57437));
    defparam i1_2_lut_3_lut_4_lut_adj_1158.LUT_INIT = 16'hffdf;
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29828), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29827), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1159 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[21] [7]), 
            .I2(n53137), .I3(n6_adj_5362), .O(n57981));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h9669;
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29826), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1160 (.I0(n57981), .I1(n52188), .I2(\data_out_frame[23] [7]), 
            .I3(n52984), .O(n53107));
    defparam i3_4_lut_adj_1160.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1161 (.I0(n57839), .I1(\data_out_frame[15] [6]), 
            .I2(n51944), .I3(n57876), .O(n10_adj_5363));
    defparam i4_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(n51970), .I1(n52973), .I2(GND_net), 
            .I3(GND_net), .O(n53172));
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29825), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1163 (.I0(n51995), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[13] [5]), .I3(n57876), .O(n10_adj_5364));
    defparam i4_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1164 (.I0(n25162), .I1(n10_adj_5364), .I2(\data_out_frame[17] [7]), 
            .I3(GND_net), .O(n59919));
    defparam i5_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29824), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1165 (.I0(n40928), .I1(n3470), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n10), .O(n172));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1165.LUT_INIT = 16'hfffb;
    SB_LUT4 i4_4_lut_adj_1166 (.I0(n7_adj_5365), .I1(n57722), .I2(n57856), 
            .I3(n59919), .O(n52042));
    defparam i4_4_lut_adj_1166.LUT_INIT = 16'h9669;
    SB_LUT4 i23_2_lut (.I0(n23735), .I1(\data_out_frame[20][3] ), .I2(GND_net), 
            .I3(GND_net), .O(n26539));   // verilog/coms.v(100[12:26])
    defparam i23_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29823), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29822), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1167 (.I0(n40928), .I1(n3470), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n10_adj_5304), .O(n28413));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1167.LUT_INIT = 16'hfffb;
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29821), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29820), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29819), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29818), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29817), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29816), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29815), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29814), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29813), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29812), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29811), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_out_frame[15] [7]), .I1(n57839), 
            .I2(GND_net), .I3(GND_net), .O(n53042));
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29810), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5366), .S(n57193));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5367), .S(n57192));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29809), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5368), .S(n57191));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5369), .S(n57190));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29808), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1169 (.I0(\data_out_frame[19] [0]), .I1(n57747), 
            .I2(n68629), .I3(n62546), .O(n58093));
    defparam i1_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29807), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29806), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29805), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5370), .S(n57189));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1170 (.I0(\data_out_frame[17] [4]), .I1(n57531), 
            .I2(n25734), .I3(n57750), .O(n52663));
    defparam i3_4_lut_adj_1170.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5371), .S(n57188));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5372), .S(n57187));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5373), .S(n57186));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5374), .S(n57114));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(GND_net), .I3(GND_net), .O(n57722));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i52884_3_lut_4_lut (.I0(rx_data[7]), .I1(\data_in_frame[16] [7]), 
            .I2(reset), .I3(n105), .O(n56594));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i52884_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5375), .S(n57115));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5376), .S(n57116));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5377), .S(n57117));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1172 (.I0(\data_out_frame[13] [7]), .I1(n52068), 
            .I2(n58111), .I3(n52024), .O(n14_adj_5378));
    defparam i6_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1173 (.I0(\data_out_frame[14] [1]), .I1(n14_adj_5378), 
            .I2(n10_adj_5379), .I3(n58123), .O(n60167));
    defparam i7_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(n60167), .I1(n57709), .I2(GND_net), 
            .I3(GND_net), .O(n53003));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1175 (.I0(n60167), .I1(n26731), .I2(n26432), 
            .I3(n1699), .O(n57470));
    defparam i3_4_lut_adj_1175.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5380), .S(n57118));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1176 (.I0(\data_out_frame[16] [2]), .I1(n57470), 
            .I2(n53178), .I3(GND_net), .O(n59803));
    defparam i2_3_lut_adj_1176.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5381), .S(n57119));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1177 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57599));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5382), .S(n57121));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5383), .S(n57122));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57856));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[18][4] ), .I1(n59803), 
            .I2(GND_net), .I3(GND_net), .O(n57845));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n62384));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5384), .S(n57123));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5385), .S(n57124));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5386), .S(n57125));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1181 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[19] [5]), .I3(GND_net), .O(n62386));
    defparam i1_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1182 (.I0(n57856), .I1(n62386), .I2(n2076), .I3(n62384), 
            .O(n62394));
    defparam i1_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1183 (.I0(n62394), .I1(n26664), .I2(n25848), 
            .I3(n57599), .O(n62398));
    defparam i1_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5387), .S(n57126));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1184 (.I0(n57455), .I1(n52198), .I2(n26279), 
            .I3(n62398), .O(n62404));
    defparam i1_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1185 (.I0(n58080), .I1(n51995), .I2(n26899), 
            .I3(n62404), .O(n62410));
    defparam i1_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5388), .S(n57127));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1186 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[17][3] ), .I3(\data_out_frame[17] [1]), 
            .O(n62562));   // verilog/coms.v(79[16:43])
    defparam i1_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5389), .S(n57128));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5390), .S(n57129));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1187 (.I0(n57744), .I1(n57608), .I2(n53178), 
            .I3(n62410), .O(n62416));
    defparam i1_4_lut_adj_1187.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1188 (.I0(n51946), .I1(n68629), .I2(n26896), 
            .I3(n62566), .O(n60272));   // verilog/coms.v(79[16:43])
    defparam i1_4_lut_adj_1188.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1189 (.I0(n60272), .I1(n59475), .I2(n62416), 
            .I3(n60035), .O(n23733));
    defparam i1_4_lut_adj_1189.LUT_INIT = 16'h9669;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29767));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1190 (.I0(n57782), .I1(n58056), .I2(\data_in_frame[14] [7]), 
            .I3(n26517), .O(n60044));
    defparam i2_3_lut_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i15926_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n30002));
    defparam i15926_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5391), .S(n57130));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3416), .CO(n49542));
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5392), .S(n57131));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5393), .S(n57111));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18][4] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5394), .S(n57132));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5395), .S(n57133));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5396), .S(n57134));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29760));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29759));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29758));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29757));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1191 (.I0(n52663), .I1(\data_out_frame[19] [5]), 
            .I2(n52175), .I3(GND_net), .O(n52984));
    defparam i1_3_lut_adj_1191.LUT_INIT = 16'h6969;
    SB_LUT4 select_777_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5297));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5296));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29756));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29755));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29754));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29753));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5397), .S(n57135));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1192 (.I0(\data_out_frame[20]_c [4]), .I1(\data_out_frame[20]_c [2]), 
            .I2(n4_adj_5398), .I3(n57571), .O(n2217));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(n2217), .I1(\data_out_frame[20]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n62322));
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1194 (.I0(n52984), .I1(n23733), .I2(n57845), 
            .I3(n62322), .O(n52492));
    defparam i1_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29752));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29750));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29749));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29748));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5399), .S(n57136));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29747));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5295));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5294));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5400), .S(n57137));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29746));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29745));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29744));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29743));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29742));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5401), .S(n57138));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1195 (.I0(n10), .I1(n3470), .I2(n161), 
            .I3(n31), .O(n28439));
    defparam i1_2_lut_3_lut_4_lut_adj_1195.LUT_INIT = 16'hffbf;
    SB_LUT4 select_777_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5293));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5402), .S(n57139));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1196 (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[20]_c [0]), 
            .I2(n57848), .I3(n6_adj_5403), .O(n53027));
    defparam i4_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(n59944), .I1(n52492), .I2(GND_net), 
            .I3(GND_net), .O(n53209));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h9999;
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29738));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14412_4_lut_4_lut (.I0(n3470), .I1(reset), .I2(n59293), .I3(n10), 
            .O(n7_adj_10));
    defparam i14412_4_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 select_777_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5292));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5291));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5405), .S(n57140));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5290));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29735));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5289));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1198 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[11] [6]), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5288));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1198.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5287));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n57245));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1199 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n57244));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1199.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5286));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1200 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n57243));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1200.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5285));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1201 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n57242));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1201.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5284));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1202 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n57294));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1202.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_out_frame[22] [1]), .I1(n23733), 
            .I2(GND_net), .I3(GND_net), .O(n57799));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5283));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1204 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n57241));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1204.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1205 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n57113));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1205.LUT_INIT = 16'h4500;
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29734));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29733));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29732));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1206 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n57240));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1206.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1207 (.I0(n52236), .I1(n25), .I2(\data_out_frame[20]_c [5]), 
            .I3(\data_out_frame[21] [7]), .O(n62376));
    defparam i1_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29730));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1208 (.I0(n57799), .I1(n53209), .I2(n53027), 
            .I3(n62376), .O(n57905));
    defparam i1_4_lut_adj_1208.LUT_INIT = 16'h9669;
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29729));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29725));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1209 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n57239));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1209.LUT_INIT = 16'h4500;
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29721));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53886 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n69643));
    defparam byte_transmit_counter_0__bdd_4_lut_53886.LUT_INIT = 16'he4aa;
    SB_LUT4 n69643_bdd_4_lut (.I0(n69643), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n63029));
    defparam n69643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29720));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5281));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1210 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n57238));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1210.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5280));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1211 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n57237));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1211.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_out_frame[9] [0]), .I1(n58030), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5406));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1213 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[11] [1]), 
            .I2(n57953), .I3(n6_adj_5406), .O(n25734));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1214 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n57236));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1214.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5279));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1215 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n57235));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1215.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5278));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5277));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53876 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n69631));
    defparam byte_transmit_counter_0__bdd_4_lut_53876.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1216 (.I0(n36), .I1(n58008), .I2(\data_out_frame[11] [2]), 
            .I3(n6_adj_5407), .O(n51944));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5276));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1217 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n57234));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1217.LUT_INIT = 16'h4500;
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29719));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1218 (.I0(\data_out_frame[19] [7]), .I1(n51944), 
            .I2(n57622), .I3(n25734), .O(n57848));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5275));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1219 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n57233));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1219.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1220 (.I0(n26291), .I1(\data_out_frame[15] [3]), 
            .I2(n25734), .I3(GND_net), .O(n57604));
    defparam i2_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1221 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n57232));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1221.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1222 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n57231));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1222.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5274));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1223 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n57230));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1223.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5273));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(n57604), .I1(n57848), .I2(GND_net), 
            .I3(GND_net), .O(n58080));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1225 (.I0(n52107), .I1(n57936), .I2(n57516), 
            .I3(\data_in_frame[13] [4]), .O(n52684));
    defparam i2_3_lut_4_lut_adj_1225.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5272));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5271));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_3_lut_4_lut (.I0(n52107), .I1(n57936), .I2(\data_in_frame[13] [3]), 
            .I3(n8_adj_5408), .O(n60454));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29718));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5270));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5269));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1226 (.I0(\data_out_frame[17] [7]), .I1(n51960), 
            .I2(\data_out_frame[18] [0]), .I3(n6_adj_5409), .O(n52516));
    defparam i4_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5268));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1227 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22][3] ), 
            .I2(n52516), .I3(GND_net), .O(n59292));
    defparam i2_3_lut_adj_1227.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_out_frame[20]_c [1]), .I1(\data_out_frame[20][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n57571));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1229 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n57229));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1229.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1230 (.I0(n59919), .I1(\data_out_frame[18] [1]), 
            .I2(n52973), .I3(GND_net), .O(n23735));
    defparam i2_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1231 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n57228));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1231.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5267));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1232 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n57227));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1232.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1233 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n57226));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1233.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1234 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n57225));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1234.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5266));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1235 (.I0(n57641), .I1(n57996), .I2(n57879), 
            .I3(n59684), .O(n57644));
    defparam i1_2_lut_3_lut_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1236 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n57224));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1236.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1237 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [0]), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5264));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1237.LUT_INIT = 16'ha088;
    SB_LUT4 n69631_bdd_4_lut (.I0(n69631), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n69634));
    defparam n69631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1238 (.I0(\data_out_frame[25] [7]), .I1(n26412), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n57789));
    defparam i2_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1239 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n57223));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1239.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5263));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(n52338), .I1(n26623), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n57833));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1241 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n57222));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1241.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_3_lut_adj_1242 (.I0(n52338), .I1(n26623), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n57499));
    defparam i1_2_lut_3_lut_adj_1242.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1243 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n57221));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1243.LUT_INIT = 16'h4500;
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29700));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29699));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n29692));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29679));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29673), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29665), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29664));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29663));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29662));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29661), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29660), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29644), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5410), .S(n57141));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1244 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n57220));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1244.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(n57885), .I1(n53107), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5411));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1246 (.I0(n53119), .I1(n57789), .I2(n52026), 
            .I3(n52991), .O(n12_adj_5412));
    defparam i5_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1247 (.I0(n25990), .I1(n57936), .I2(\data_in_frame[13] [4]), 
            .I3(\data_in_frame[18] [0]), .O(n58021));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i13_2_lut (.I0(pwm_setpoint[22]), .I1(\pwm_counter[22] ), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/pwm.v(11[19:30])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1248 (.I0(n25990), .I1(n57936), .I2(\data_in_frame[13] [3]), 
            .I3(GND_net), .O(n57516));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_LUT4 i15_2_lut (.I0(pwm_setpoint[21]), .I1(\pwm_counter[21] ), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_11));   // verilog/pwm.v(11[19:30])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5414), .S(n57142));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5415), .S(n57143));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20]_c [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5416), .S(n57144));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20]_c [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5417), .S(n29019));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20]_c [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5418), .S(n57145));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_209_i3_4_lut (.I0(n53207), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n12_adj_5412), .I3(n8_adj_5411), .O(n3_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5420), .S(n29017));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20]_c [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5421), .S(n57146));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20]_c [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5422), .S(n57147));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5423), .S(n57148));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5424), .S(n57149));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21][0] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5425), .S(n57150));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5426), .S(n29011));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5427), .S(n57151));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5428), .S(n57152));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_2_lut_4_lut (.I0(\data_in_frame[19] [2]), .I1(n53127), .I2(n53102), 
            .I3(n57541), .O(n24_adj_5429));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5430), .S(n57153));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1249 (.I0(\data_in_frame[19] [2]), .I1(n53127), 
            .I2(n53102), .I3(\data_in_frame[21] [4]), .O(n57615));
    defparam i1_2_lut_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5431), .S(n57154));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5432), .S(n57155));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5433), .S(n57156));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5434), .S(n57157));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5435), .S(n57158));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5436), .S(n57159));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5437), .S(n57160));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5438), .S(n57161));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5439), .S(n57162));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1250 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n57219));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1250.LUT_INIT = 16'h4500;
    SB_LUT4 i1288_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(88[17:28])
    defparam i1288_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_out_frame[16] [6]), .I1(n26795), 
            .I2(GND_net), .I3(GND_net), .O(n57522));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1252 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n57218));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1252.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1253 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n57217));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1253.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1254 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n57216));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1254.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1255 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n57215));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1255.LUT_INIT = 16'h4500;
    SB_LUT4 i5_4_lut_adj_1256 (.I0(n26896), .I1(n57688), .I2(n58042), 
            .I3(n53095), .O(n12_adj_5441));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1256.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1257 (.I0(n57522), .I1(n12_adj_5441), .I2(n57747), 
            .I3(\data_out_frame[19] [0]), .O(n60087));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1258 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n57214));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1258.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1259 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n57213));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1259.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1260 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n57212));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1260.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1261 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n57211));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1261.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5442));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1262 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n57210));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1262.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1263 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n29076));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1263.LUT_INIT = 16'h4500;
    SB_DFFR \FRAME_MATCHER.i_1942__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n28080), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1264 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n57209));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1264.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1265 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n57208));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1265.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5444), .S(n57163));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5445), .S(n57164));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5443), .S(n57165));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[17] [0]), .I1(n57455), 
            .I2(GND_net), .I3(GND_net), .O(n26896));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5442), .S(n57166));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1942__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n28082), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n28084), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n28086), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n28088), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n28090), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n28092), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n28094), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n28096), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n28098), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n28100), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n28102), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n28104), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n28106), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28108), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28110), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28112), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28114), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28116), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28118), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28120), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28122), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28124), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28126), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28128), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28130), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28132), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i5  (.Q(\FRAME_MATCHER.i[5] ), .C(clk16MHz), 
            .D(n28134), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i4  (.Q(\FRAME_MATCHER.i[4] ), .C(clk16MHz), 
            .D(n28136), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n28138), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n28140), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n28142), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5440), .S(n57167));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1267 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n57207));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1267.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1268 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n57206));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1268.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_adj_1269 (.I0(n1168), .I1(n57476), .I2(\data_out_frame[7] [0]), 
            .I3(n58030), .O(n6_adj_5446));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1270 (.I0(n1168), .I1(n57476), .I2(\data_out_frame[7] [0]), 
            .I3(n26380), .O(n57939));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1271 (.I0(\data_out_frame[12] [7]), .I1(n36), .I2(n57950), 
            .I3(GND_net), .O(n14_adj_5447));
    defparam i5_3_lut_adj_1271.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1272 (.I0(n58126), .I1(\data_out_frame[13] [1]), 
            .I2(n25702), .I3(n58017), .O(n15_c));
    defparam i6_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1273 (.I0(n15_c), .I1(n57534), .I2(n14_adj_5447), 
            .I3(n26645), .O(n26291));
    defparam i8_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5448));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1275 (.I0(n57452), .I1(n57921), .I2(\data_out_frame[10] [4]), 
            .I3(GND_net), .O(n60077));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1275.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5360), .S(n57293));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5358), .S(n57292));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5357), .S(n57291));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5356), .S(n57290));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1276 (.I0(\data_out_frame[7] [7]), .I1(n58108), 
            .I2(\data_out_frame[14] [4]), .I3(n26279), .O(n57455));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5354), .S(n57289));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5352), .S(n57288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5349), .S(n57287));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1277 (.I0(n1516), .I1(\data_out_frame[12] [4]), 
            .I2(n60077), .I3(n4_adj_5448), .O(n26795));
    defparam i2_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(n26795), .I1(n57574), .I2(GND_net), 
            .I3(GND_net), .O(n52635));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1279 (.I0(\data_out_frame[7] [7]), .I1(n58108), 
            .I2(n52198), .I3(GND_net), .O(n53159));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1280 (.I0(\data_out_frame[7] [7]), .I1(n58108), 
            .I2(n52209), .I3(n26279), .O(n53095));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5345), .S(n57286));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14005_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3470), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n28080));   // verilog/coms.v(158[12:15])
    defparam i14005_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_33_lut  (.I0(n65673), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n50838), .O(n28082)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_32_lut  (.I0(n65663), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n50837), .O(n28084)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_32  (.CI(n50837), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n50838));
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5344), .S(n57285));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_31_lut  (.I0(n65662), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n50836), .O(n28086)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5343), .S(n57284));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_31  (.CI(n50836), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n50837));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_30_lut  (.I0(n65661), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n50835), .O(n28088)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_30  (.CI(n50835), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n50836));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_29_lut  (.I0(n65660), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n50834), .O(n28090)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_29  (.CI(n50834), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n50835));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_28_lut  (.I0(n65649), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n50833), .O(n28092)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_28  (.CI(n50833), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n50834));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_27_lut  (.I0(n65617), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n50832), .O(n28094)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_27  (.CI(n50832), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n50833));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_26_lut  (.I0(n65616), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n50831), .O(n28096)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_26  (.CI(n50831), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n50832));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_25_lut  (.I0(n65615), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n50830), .O(n28098)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_25  (.CI(n50830), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n50831));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_24_lut  (.I0(n65609), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n50829), .O(n28100)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_24  (.CI(n50829), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n50830));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_23_lut  (.I0(n65608), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n50828), .O(n28102)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_23  (.CI(n50828), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n50829));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_22_lut  (.I0(n65593), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n50827), .O(n28104)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_22  (.CI(n50827), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n50828));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_21_lut  (.I0(n65592), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n50826), .O(n28106)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_21  (.CI(n50826), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n50827));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_20_lut  (.I0(n65586), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n50825), .O(n28108)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_20  (.CI(n50825), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n50826));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_19_lut  (.I0(n65582), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n50824), .O(n28110)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_19  (.CI(n50824), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n50825));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_18_lut  (.I0(n65581), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n50823), .O(n28112)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_18  (.CI(n50823), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n50824));
    SB_LUT4 i4_4_lut_adj_1281 (.I0(\data_out_frame[17][3] ), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(n6_adj_5449), .O(n52175));
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_17_lut  (.I0(n65572), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n50822), .O(n28114)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_17  (.CI(n50822), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n50823));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_16_lut  (.I0(n65571), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n50821), .O(n28116)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_16  (.CI(n50821), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n50822));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_15_lut  (.I0(n65570), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n50820), .O(n28118)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_15  (.CI(n50820), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n50821));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_14_lut  (.I0(n65563), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n50819), .O(n28120)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_14  (.CI(n50819), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n50820));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_13_lut  (.I0(n65558), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n50818), .O(n28122)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_13  (.CI(n50818), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n50819));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_12_lut  (.I0(n65557), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n50817), .O(n28124)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_12  (.CI(n50817), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n50818));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_11_lut  (.I0(n65556), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n50816), .O(n28126)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_11  (.CI(n50816), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n50817));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_10_lut  (.I0(n65555), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n50815), .O(n28128)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_10  (.CI(n50815), .I0(n28404), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n50816));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_9_lut  (.I0(n65554), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n50814), .O(n28130)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_9  (.CI(n50814), .I0(n28404), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n50815));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_8_lut  (.I0(n65553), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n50813), .O(n28132)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_8  (.CI(n50813), .I0(n28404), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n50814));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_7_lut  (.I0(n65552), .I1(n28404), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n50812), .O(n28134)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_7  (.CI(n50812), .I0(n28404), .I1(\FRAME_MATCHER.i[5] ), 
            .CO(n50813));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_6_lut  (.I0(n65551), .I1(n28404), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(n50811), .O(n28136)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_6  (.CI(n50811), .I0(n28404), .I1(\FRAME_MATCHER.i[4] ), 
            .CO(n50812));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_5_lut  (.I0(n65550), .I1(n28404), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n50810), .O(n28138)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_5  (.CI(n50810), .I0(n28404), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n50811));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_4_lut  (.I0(n65549), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n50809), .O(n28140)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_4  (.CI(n50809), .I0(n28404), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n50810));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_3_lut  (.I0(n65548), .I1(n28404), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n50808), .O(n28142)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_3  (.CI(n50808), .I0(n28404), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n50809));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n50808));
    SB_LUT4 i2_3_lut_adj_1282 (.I0(n52175), .I1(\data_out_frame[19] [4]), 
            .I2(n52635), .I3(GND_net), .O(n52188));
    defparam i2_3_lut_adj_1282.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n29471));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57688));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26138));
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n30549), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n30548), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n30547), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n30546), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n30545), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n30544), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n30543), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n29474));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n30534));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n29477));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1285 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n57205));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1285.LUT_INIT = 16'h4500;
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n29480));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_out_frame[6] [1]), .I1(n25705), 
            .I2(GND_net), .I3(GND_net), .O(n25702));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n29483));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30512));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n29486));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n29489));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n29492));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30506));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n29495));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n30504), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n30503), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n29498));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n30501));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n30500), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n30499), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n30498), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n56504));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n30490), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1287 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n57953));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1287.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1288 (.I0(n26282), .I1(\data_out_frame[10] [2]), 
            .I2(n53133), .I3(n26104), .O(n60324));
    defparam i1_3_lut_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n30466), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30439), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n30431), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n29504));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30429), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30428), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n30002));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n30415));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30414));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30413));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30412));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30411));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30410));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30409));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30408));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30407));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30406));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30405));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30404));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[19] [1]), .I1(n53199), .I2(\data_out_frame[18] [7]), 
            .I3(\data_out_frame[20]_c [4]), .O(n18));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58017));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1290 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[6] [4]), .O(n62454));
    defparam i1_4_lut_adj_1290.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30403));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30402));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30401));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30400));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30399));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30398));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5450), .S(n57283));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30397));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30396));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30395));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30394));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30393));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30392));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30391));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30390));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1291 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[7] [4]), .O(n62456));
    defparam i1_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30389));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1292 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[9] [1]), .I3(\data_out_frame[9] [6]), .O(n62424));
    defparam i1_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30388));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_1650_Select_0_i1_2_lut_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n43569), .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n1));   // verilog/coms.v(148[4] 304[11])
    defparam select_1650_Select_0_i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1293 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n57204));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1293.LUT_INIT = 16'h4500;
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30387));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1294 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[8] [4]), .O(n62458));
    defparam i1_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30386));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30385));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30384));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1295 (.I0(\data_out_frame[19] [1]), .I1(n53199), 
            .I2(\data_out_frame[18] [7]), .I3(\data_out_frame[16] [4]), 
            .O(n58042));
    defparam i1_2_lut_4_lut_adj_1295.LUT_INIT = 16'h9669;
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30383), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30382), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n30381));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30380), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5451), .S(n57282));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n30006));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30378), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n30009));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n56568));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n30012));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30372));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n30371));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n30370));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n56566));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n29520));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1296 (.I0(n58129), .I1(n57577), .I2(n62458), 
            .I3(n58036), .O(n62472));
    defparam i1_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n29523));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n29526));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n29530));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n56594));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n56478));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n56474));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n56470));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n56466));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n56462));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n30015));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n30019));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n30022));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5452), .S(n57281));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n56458));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30343));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n56454));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n56450));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n56446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n30025));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n30028));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n30336));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n30031));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
           .D(n30034));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
           .D(n30037));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
           .D(n30040));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
           .D(n30043));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6]_c [6]), .C(clk16MHz), 
           .D(n30046));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1297 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n57203));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1297.LUT_INIT = 16'h4500;
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6]_c [7]), .C(clk16MHz), 
           .D(n30049));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n56514));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7][1] ), .C(clk16MHz), 
           .D(n30055));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7][2] ), .C(clk16MHz), 
           .D(n30059));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7][3] ), .C(clk16MHz), 
           .D(n30062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7][4] ), .C(clk16MHz), 
           .D(n30065));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7][5] ), .C(clk16MHz), 
           .D(n30068));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n56520));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
           .D(n56518));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n30077));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n30080));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n30083));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n30317));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n30316));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5453), .S(n57280));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
           .D(n30087));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
           .D(n30314));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1298 (.I0(n62456), .I1(n62466), .I2(n1130), .I3(n62454), 
            .O(n62474));
    defparam i1_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1299 (.I0(n62472), .I1(n26645), .I2(n57953), 
            .I3(GND_net), .O(n62476));
    defparam i1_3_lut_adj_1299.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
           .D(n30093));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
           .D(n30096));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
           .D(n30099));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n30102));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n30105));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n30108));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n30112));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n30115));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n30118));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n30122));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n30125));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10]_c [0]), .C(clk16MHz), 
           .D(n30128));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10][1] ), .C(clk16MHz), 
           .D(n30131));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10][2] ), .C(clk16MHz), 
           .D(n30134));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10][3] ), .C(clk16MHz), 
           .D(n30138));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n30141));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1300 (.I0(n58002), .I1(n57558), .I2(n57968), 
            .I3(n62424), .O(n62430));
    defparam i1_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10][5] ), .C(clk16MHz), 
           .D(n30144));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n30148));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10][7] ), .C(clk16MHz), 
           .D(n30151));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n30154));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n56662));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n56678));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n56604));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n30167));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n30170));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n30173));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n30287));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30177));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30180));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n30183));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n30186));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n56636));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n56690));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n30196));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n30199));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n30203));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n30206));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30209));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n30213));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30216));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n30219));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n30223));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1301 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n57202));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1301.LUT_INIT = 16'h4500;
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n30226));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1302 (.I0(n25702), .I1(n57962), .I2(n62476), 
            .I3(n62474), .O(n62482));
    defparam i1_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n30260));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n56442));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n56438));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n30265));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1303 (.I0(n26461), .I1(n62482), .I2(n62430), 
            .I3(n26844), .O(n53133));
    defparam i1_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29570));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n29573));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29576));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n56434));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n56430));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n56546));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n56542));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1304 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n57201));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1304.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_179_i2_4_lut (.I0(\data_out_frame[22][3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n56540));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29594));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n56538));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n56536));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n56534));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19]_c [7]), .C(clk16MHz), 
           .D(n56554));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n29609));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n30229));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n30222));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29618));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1305 (.I0(n26461), .I1(n53133), .I2(n62300), 
            .I3(n58017), .O(n58123));
    defparam i1_4_lut_adj_1305.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29621));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1306 (.I0(n26553), .I1(n58123), .I2(\data_out_frame[10] [2]), 
            .I3(\data_out_frame[10] [1]), .O(n52068));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5436));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1307 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n57200));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1307.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n29624));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1308 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n57199));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1308.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5434));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1309 (.I0(n60324), .I1(n52068), .I2(\data_out_frame[8] [3]), 
            .I3(GND_net), .O(n57950));
    defparam i1_3_lut_adj_1309.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1310 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n57198));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1310.LUT_INIT = 16'h4500;
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n30176));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1311 (.I0(n52635), .I1(n57908), .I2(\data_out_frame[19][3] ), 
            .I3(\data_out_frame[21] [5]), .O(n57812));
    defparam i2_3_lut_4_lut_adj_1311.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n29632));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1312 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n57197));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1312.LUT_INIT = 16'h4500;
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29638));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1313 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[10] [7]), .I3(\data_out_frame[12] [6]), 
            .O(n62488));
    defparam i1_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1314 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [5]), 
            .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1314.LUT_INIT = 16'ha088;
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29641));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29646));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1315 (.I0(n10_adj_5323), .I1(reset), 
            .I2(n58272), .I3(n8), .O(n57425));
    defparam i1_2_lut_3_lut_4_lut_adj_1315.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1316 (.I0(\data_out_frame[20]_c [5]), 
            .I1(\data_out_frame[20] [6]), .I2(\data_out_frame[20] [7]), 
            .I3(\data_out_frame[22] [7]), .O(n58083));
    defparam i1_2_lut_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1317 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [4]), 
            .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5430));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1317.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1318 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n57196));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1318.LUT_INIT = 16'h4500;
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29649));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1319 (.I0(\data_out_frame[13] [0]), .I1(n62492), 
            .I2(n57950), .I3(n57918), .O(n57750));
    defparam i1_4_lut_adj_1319.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29657));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57531));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1321 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21][3] ), 
            .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5428));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1322 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n57195));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1322.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5427));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i53010_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n43569), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i53010_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29666));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5426));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1323 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n29060));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1323.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1324 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n57194));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1324.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1325 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n57193));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1325.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_168_i2_4_lut (.I0(\data_out_frame[21][0] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5425));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1326 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n57192));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1326.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5424));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1327 (.I0(n10_adj_5323), .I1(reset), 
            .I2(n58272), .I3(n8_adj_12), .O(n57426));
    defparam i1_2_lut_3_lut_4_lut_adj_1327.LUT_INIT = 16'hffef;
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5456), .S(n57279));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1328 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [6]), 
            .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5423));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1328.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_adj_1329 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n57534));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1329.LUT_INIT = 16'h9696;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1330 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n57191));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1330.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5457), .S(n57278));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5458), .S(n57277));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5459), .S(n57276));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1331 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20]_c [5]), 
            .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1331.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5460), .S(n57275));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1332 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n57190));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1332.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_164_i2_4_lut (.I0(\data_out_frame[20]_c [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5421));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1333 (.I0(n1130), .I1(n57534), .I2(n25705), .I3(\data_out_frame[13] [2]), 
            .O(n58030));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1334 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n57189));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1334.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1335 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20][3] ), 
            .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5420));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1335.LUT_INIT = 16'ha088;
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29680));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57590));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1337 (.I0(n57496), .I1(n1130), .I2(\data_out_frame[11] [4]), 
            .I3(n57939), .O(n10_adj_5461));
    defparam i4_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29536));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1338 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n57188));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1338.LUT_INIT = 16'h4500;
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29529), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1339 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n57187));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1339.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_162_i2_4_lut (.I0(\data_out_frame[20]_c [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5462), .S(n57274));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1340 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n57186));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1340.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1341 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20]_c [1]), 
            .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1341.LUT_INIT = 16'ha088;
    SB_LUT4 i4_4_lut_adj_1342 (.I0(n57590), .I1(n58105), .I2(n57939), 
            .I3(\data_out_frame[13] [4]), .O(n10_adj_5463));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5464), .S(n57273));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27767), 
            .D(n4762[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27767), 
            .D(n4762[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27767), 
            .D(n4762[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27767), 
            .D(n4762[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27767), 
            .D(n4762[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27767), 
            .D(n4762[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27767), 
            .D(n4762[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1343 (.I0(\data_in_frame[18] [7]), .I1(n51958), 
            .I2(n57999), .I3(n6_adj_5465), .O(n52036));
    defparam i4_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27767), 
            .D(n4762[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27767), 
            .D(n4762[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1344 (.I0(\data_out_frame[5] [0]), .I1(n10_adj_5463), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n57672));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1344.LUT_INIT = 16'h9696;
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27767), 
            .D(n4762[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1345 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n57114));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1345.LUT_INIT = 16'h4500;
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27767), 
            .D(n4762[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1346 (.I0(n26432), .I1(n52024), .I2(GND_net), 
            .I3(GND_net), .O(n53030));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27767), 
            .D(n4762[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_160_i2_4_lut (.I0(\data_out_frame[20]_c [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27767), 
            .D(n4762[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1347 (.I0(\data_in_frame[20] [0]), .I1(\data_in_frame[19]_c [7]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n57541));
    defparam i2_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27767), 
            .D(n4762[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27767), 
            .D(n4762[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27767), 
            .D(n4762[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27767), 
            .D(n4762[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27767), 
            .D(n4762[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27767), 
            .D(n4762[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27767), 
            .D(n4762[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27767), 
            .D(n4762[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57999));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27767), 
            .D(n4762[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27767), 
            .D(n4762[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5466), .S(n57272));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1349 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16][3] ), 
            .O(n57115));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1349.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1350 (.I0(n51954), .I1(\data_in_frame[20] [3]), 
            .I2(n57525), .I3(\data_in_frame[20] [4]), .O(n57706));
    defparam i3_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1351 (.I0(n26738), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[18] [4]), .O(n57816));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1352 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[18] [5]), 
            .I2(n53052), .I3(GND_net), .O(n58061));
    defparam i1_3_lut_adj_1352.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1353 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n57116));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1353.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1354 (.I0(\data_in_frame[20] [7]), .I1(n57644), 
            .I2(GND_net), .I3(GND_net), .O(n58120));
    defparam i1_2_lut_adj_1354.LUT_INIT = 16'h6666;
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n69866), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n27046), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2048), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state [3]), .C(clk16MHz), 
            .D(n2049), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20442), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n56292), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2060), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n27049), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5467), .S(n57271));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1355 (.I0(\data_out_frame[11] [2]), .I1(n25709), 
            .I2(n57700), .I3(n6_adj_5446), .O(n1720));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1356 (.I0(\data_in_frame[15] [5]), .I1(n52684), 
            .I2(n60454), .I3(GND_net), .O(n25808));
    defparam i2_3_lut_adj_1356.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57622));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1358 (.I0(n59240), .I1(n25808), .I2(Kp_23__N_1551), 
            .I3(GND_net), .O(n57956));
    defparam i2_3_lut_adj_1358.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5468), .S(n57270));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1359 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26282));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1359.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1360 (.I0(n57502), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(n57942), .O(n10_adj_5469));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5470), .S(n57269));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1361 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57681));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1361.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5471), .S(n57268));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5472), .S(n57267));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5473), .S(n57266));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1362 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n57117));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1362.LUT_INIT = 16'h4500;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1363 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n57118));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1363.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1364 (.I0(n10_adj_5323), .I1(reset), 
            .I2(n58272), .I3(n8_adj_13), .O(n57424));
    defparam i1_2_lut_3_lut_4_lut_adj_1364.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1365 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n57119));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1365.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1366 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n25937));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1366.LUT_INIT = 16'h6666;
    SB_LUT4 i23277_3_lut (.I0(n380), .I1(n460), .I2(n11610), .I3(GND_net), 
            .O(n27722));
    defparam i23277_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5475), .S(n57265));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1367 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n57121));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1367.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5476), .S(n57264));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1368 (.I0(\data_in_frame[21] [2]), .I1(n57644), 
            .I2(n25937), .I3(n57764), .O(n57634));
    defparam i1_4_lut_adj_1368.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5477), .S(n57263));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\data_in_frame[19] [0]), .I1(n52141), 
            .I2(GND_net), .I3(GND_net), .O(n57764));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5478), .S(n57262));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1370 (.I0(n53102), .I1(\data_in_frame[21] [5]), 
            .I2(n59871), .I3(GND_net), .O(n57984));
    defparam i2_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5479), .S(n57261));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29684));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5480), .S(n57260));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5481), .S(n57259));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5482), .S(n57258));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1371 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n57122));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1371.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5483), .S(n57257));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5484), .S(n57256));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5485), .S(n57255));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29510));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1372 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[21] [6]), 
            .I2(n57984), .I3(GND_net), .O(n20));
    defparam i1_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[21] [1]), .I1(n22_adj_5486), .I2(n57764), 
            .I3(n57634), .O(n30_c));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57476));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1374 (.I0(\data_out_frame[10] [0]), .I1(n26104), 
            .I2(GND_net), .I3(GND_net), .O(n26553));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1374.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1375 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57968));
    defparam i1_2_lut_adj_1375.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1376 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n57942));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1377 (.I0(\data_in_frame[20] [2]), .I1(n33), .I2(n38), 
            .I3(n34), .O(n28));
    defparam i9_4_lut_adj_1377.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut (.I0(n57564), .I1(n30_c), .I2(n20), .I3(n57615), 
            .O(n34_adj_5487));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1378 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n57123));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1378.LUT_INIT = 16'h4500;
    SB_LUT4 i13_4_lut_adj_1379 (.I0(n58120), .I1(n58021), .I2(n58061), 
            .I3(n57816), .O(n32_c));
    defparam i13_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n57706), .I1(n34_adj_5487), .I2(n28), .I3(\data_in_frame[15] [6]), 
            .O(n36_adj_5488));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1380 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17][3] ), 
            .O(n57124));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1380.LUT_INIT = 16'h4500;
    SB_LUT4 i18_4_lut (.I0(n23_adj_5489), .I1(n36_adj_5488), .I2(n32_c), 
            .I3(n24_adj_5429), .O(n57792));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1381 (.I0(n57999), .I1(\data_in_frame[20] [6]), 
            .I2(n25937), .I3(n52449), .O(n14_adj_5490));
    defparam i6_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1382 (.I0(\data_in_frame[21] [0]), .I1(n14_adj_5490), 
            .I2(n10_adj_5491), .I3(\data_in_frame[18] [4]), .O(n52147));
    defparam i7_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(\data_in_frame[18] [3]), .I1(n25207), 
            .I2(GND_net), .I3(GND_net), .O(n51954));
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1384 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n57990));
    defparam i2_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1385 (.I0(\data_in_frame[9] [5]), .I1(n57972), 
            .I2(n57587), .I3(n57482), .O(n20_adj_5492));
    defparam i8_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1386 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[14] [7]), 
            .I2(n57737), .I3(n52995), .O(n19_c));
    defparam i7_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1387 (.I0(n57942), .I1(n57968), .I2(\data_out_frame[12] [0]), 
            .I3(GND_net), .O(n58111));
    defparam i2_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1388 (.I0(n58141), .I1(n57492), .I2(n57761), 
            .I3(\data_in_frame[10] [6]), .O(n21_c));
    defparam i9_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(n21_c), .I1(n19_c), .I2(n20_adj_5492), .I3(GND_net), 
            .O(n58039));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i21825_3_lut_4_lut (.I0(\Kp[7] ), .I1(\data_in_frame[3]_c [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29828));
    defparam i21825_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i2_3_lut_adj_1389 (.I0(n25990), .I1(n26009), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n26025));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1390 (.I0(n26069), .I1(n25891), .I2(n57990), 
            .I3(n6_adj_5493), .O(n52995));
    defparam i4_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1391 (.I0(\data_in_frame[15] [3]), .I1(n52995), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n59287));
    defparam i2_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1392 (.I0(\data_out_frame[11] [7]), .I1(n25751), 
            .I2(n57547), .I3(n6_adj_5494), .O(n52198));   // verilog/coms.v(74[16:62])
    defparam i4_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1393 (.I0(n51948), .I1(\data_in_frame[19] [4]), 
            .I2(n59240), .I3(GND_net), .O(n59871));
    defparam i2_3_lut_adj_1393.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1394 (.I0(n26025), .I1(n58039), .I2(n52684), 
            .I3(GND_net), .O(n59240));
    defparam i2_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29508));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1395 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n57125));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1395.LUT_INIT = 16'h4500;
    SB_LUT4 i5_4_lut_adj_1396 (.I0(n57675), .I1(n58011), .I2(\data_in_frame[17] [2]), 
            .I3(\data_in_frame[14] [6]), .O(n12_adj_5495));
    defparam i5_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1397 (.I0(\data_out_frame[9] [4]), .I1(n26121), 
            .I2(n57612), .I3(n25698), .O(n57896));
    defparam i3_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(74[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1398 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_5495), 
            .I2(n58045), .I3(n60044), .O(n51948));
    defparam i6_4_lut_adj_1398.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1399 (.I0(\data_in_frame[17] [1]), .I1(n51948), 
            .I2(GND_net), .I3(GND_net), .O(n52054));
    defparam i1_2_lut_adj_1399.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1400 (.I0(n52054), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[16] [7]), .I3(n58132), .O(n53102));
    defparam i2_4_lut_adj_1400.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1401 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n58045));
    defparam i1_2_lut_adj_1401.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1402 (.I0(n57756), .I1(n58045), .I2(n53024), 
            .I3(\data_in_frame[14] [5]), .O(n58132));
    defparam i3_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1403 (.I0(n59684), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[17] [0]), .I3(GND_net), .O(n57862));
    defparam i2_3_lut_adj_1403.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1404 (.I0(n57896), .I1(n52198), .I2(n58111), 
            .I3(n6_adj_5496), .O(n57709));
    defparam i4_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1405 (.I0(\data_in_frame[16] [6]), .I1(n52413), 
            .I2(GND_net), .I3(GND_net), .O(n57879));
    defparam i1_2_lut_adj_1405.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1406 (.I0(\data_in_frame[14] [6]), .I1(n26061), 
            .I2(\data_in_frame[12] [4]), .I3(n52034), .O(n52186));
    defparam i3_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(n51958), .I1(n52186), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5497));
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1408 (.I0(\data_in_frame[18] [7]), .I1(n57862), 
            .I2(\data_in_frame[19] [1]), .I3(n4_adj_5497), .O(n52141));
    defparam i2_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1409 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n57126));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1409.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1410 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n57127));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1410.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1411 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57458));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1411.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n58002));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1413 (.I0(n9), .I1(\data_out_frame[11] [5]), .I2(n8_adj_5498), 
            .I3(n57458), .O(n52024));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1414 (.I0(\data_out_frame[14] [0]), .I1(n57896), 
            .I2(\data_out_frame[11] [6]), .I3(n26104), .O(n26731));
    defparam i3_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1415 (.I0(\data_out_frame[14] [4]), .I1(n57709), 
            .I2(GND_net), .I3(GND_net), .O(n52209));
    defparam i1_2_lut_adj_1415.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1416 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[19] [2]), 
            .I2(n53127), .I3(n52141), .O(n57564));
    defparam i1_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1417 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n57128));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1417.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1418 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n57129));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1418.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1419 (.I0(\data_in_frame[9] [2]), .I1(n57482), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n26009));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1420 (.I0(\data_in_frame[16] [2]), .I1(n26009), 
            .I2(n57975), .I3(n57587), .O(n57625));
    defparam i3_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1421 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58008));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1421.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1422 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n57130));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1422.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5499), .S(n57168));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1423 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n57131));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1423.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1424 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26645));
    defparam i2_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1425 (.I0(n58114), .I1(n52094), .I2(n57516), 
            .I3(n57975), .O(n15_adj_5500));
    defparam i6_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5501), .S(n57169));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i8_4_lut_adj_1426 (.I0(n15_adj_5500), .I1(n57859), .I2(n14_adj_5502), 
            .I3(\data_in_frame[13] [6]), .O(n59679));
    defparam i8_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(n26623), .I1(n57625), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n52449));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(n25858), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5503));
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1428 (.I0(\data_in_frame[14] [4]), .I1(n52028), 
            .I2(\data_in_frame[12] [2]), .I3(n6_adj_5503), .O(n52413));
    defparam i4_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1429 (.I0(n57663), .I1(n26367), .I2(\data_in_frame[11] [3]), 
            .I3(n58005), .O(n10_adj_5504));
    defparam i4_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1430 (.I0(n57479), .I1(n10_adj_5504), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(n25990));
    defparam i5_3_lut_adj_1430.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1431 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57930));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1431.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5505), .S(n57170));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i8_4_lut_adj_1432 (.I0(n58077), .I1(n57697), .I2(\data_in_frame[5] [0]), 
            .I3(n25858), .O(n22_adj_5506));
    defparam i8_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1433 (.I0(n57842), .I1(n57631), .I2(n57719), 
            .I3(n57479), .O(n24_adj_5507));
    defparam i10_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1434 (.I0(n57822), .I1(\data_in_frame[9] [3]), 
            .I2(n57513), .I3(n58144), .O(n23_adj_5508));
    defparam i9_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1435 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18][3] ), 
            .O(n57111));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1435.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1436 (.I0(\data_in_frame[14] [2]), .I1(n25_adj_5509), 
            .I2(n23_adj_5508), .I3(n24_adj_5507), .O(n26623));
    defparam i1_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1437 (.I0(n31), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(n57410), .I3(GND_net), .O(n28409));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1437.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1438 (.I0(n57927), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[9] [3]), .I3(n57930), .O(n10_adj_5510));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1439 (.I0(\data_in_frame[11] [7]), .I1(n51992), 
            .I2(n6_c), .I3(\data_in_frame[12] [1]), .O(n57842));
    defparam i1_4_lut_adj_1439.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_1440 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[10][1] ), 
            .I2(n57842), .I3(GND_net), .O(n8_adj_5511));
    defparam i3_3_lut_adj_1440.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1441 (.I0(\data_in_frame[14] [3]), .I1(n53059), 
            .I2(n8_adj_5511), .I3(n53024), .O(n57996));
    defparam i1_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_in_frame[16] [4]), .I1(n26623), 
            .I2(GND_net), .I3(GND_net), .O(n57641));
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1443 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18][4] ), 
            .O(n57132));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1443.LUT_INIT = 16'h4500;
    SB_LUT4 i5_3_lut_adj_1444 (.I0(n57473), .I1(n10_adj_5510), .I2(\data_out_frame[9] [1]), 
            .I3(GND_net), .O(n25162));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1445 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n57133));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1445.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(n52693), .I1(n52308), .I2(GND_net), 
            .I3(GND_net), .O(n53059));
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1447 (.I0(\data_in_frame[8] [0]), .I1(n57519), 
            .I2(n25906), .I3(\data_in_frame[8] [3]), .O(n22_adj_5512));
    defparam i9_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5513), .S(n57171));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1448 (.I0(n57555), .I1(n53059), .I2(n57767), 
            .I3(GND_net), .O(n15_adj_5514));
    defparam i2_3_lut_adj_1448.LUT_INIT = 16'h6969;
    SB_LUT4 i11_4_lut_adj_1449 (.I0(n15_adj_5514), .I1(n22_adj_5512), .I2(\data_in_frame[8] [4]), 
            .I3(\data_in_frame[8] [2]), .O(n24_adj_5515));
    defparam i11_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1450 (.I0(\data_in_frame[1] [6]), .I1(n24_adj_5515), 
            .I2(n20_adj_5516), .I3(n68627), .O(n57719));
    defparam i12_4_lut_adj_1450.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(GND_net), .I3(GND_net), .O(n26715));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57492));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1453 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57558));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1453.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57612));
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1455 (.I0(\data_out_frame[7] [4]), .I1(n57612), 
            .I2(n57558), .I3(\data_out_frame[5] [1]), .O(n26104));   // verilog/coms.v(76[16:34])
    defparam i3_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5517), .S(n57172));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1456 (.I0(\data_in_frame[8] [6]), .I1(n57492), 
            .I2(n26715), .I3(n26336), .O(n57936));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1457 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n57134));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1457.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1458 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5518));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1458.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1459 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n57135));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1459.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5519), .S(n57173));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1460 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n57136));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1460.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n57097));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h4444;
    SB_LUT4 i4_4_lut_adj_1462 (.I0(n52107), .I1(Kp_23__N_974), .I2(\data_in_frame[8] [6]), 
            .I3(n6_adj_5518), .O(n58053));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1463 (.I0(\data_in_frame[10] [6]), .I1(n25976), 
            .I2(GND_net), .I3(GND_net), .O(n57782));
    defparam i1_2_lut_adj_1463.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1464 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n57137));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1464.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1465 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n57138));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1465.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1466 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(n6_adj_5520), .I3(n52107), .O(n53215));
    defparam i1_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1467 (.I0(n57782), .I1(\data_in_frame[15] [4]), 
            .I2(n58053), .I3(\data_in_frame[13] [2]), .O(n8_adj_5408));
    defparam i3_4_lut_adj_1467.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1468 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19][3] ), 
            .O(n57139));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1468.LUT_INIT = 16'h4500;
    SB_LUT4 i6_4_lut_adj_1469 (.I0(n58033), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[13] [7]), .O(n14_adj_5521));
    defparam i6_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5522), .S(n57174));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1470 (.I0(\data_out_frame[13] [5]), .I1(n25162), 
            .I2(GND_net), .I3(GND_net), .O(n26818));
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1471 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57921));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1471.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57547));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24][2] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5523), .S(n57175));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5524), .S(n57176));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5525));
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1474 (.I0(n9_adj_5525), .I1(n14_adj_5521), .I2(n57719), 
            .I3(n58072), .O(n52338));
    defparam i7_4_lut_adj_1474.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1475 (.I0(\data_in_frame[16] [1]), .I1(n26487), 
            .I2(n57443), .I3(n25990), .O(n57859));
    defparam i3_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1476 (.I0(n59598), .I1(n57859), .I2(\data_in_frame[16] [2]), 
            .I3(n52338), .O(n25207));
    defparam i3_4_lut_adj_1476.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1477 (.I0(n60454), .I1(n53215), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n59447));
    defparam i2_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25698));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1479 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n9));   // verilog/coms.v(88[17:70])
    defparam i3_3_lut_adj_1479.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5526), .S(n57177));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1480 (.I0(n57996), .I1(\data_in_frame[16] [5]), 
            .I2(n52413), .I3(GND_net), .O(n51958));
    defparam i2_3_lut_adj_1480.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1481 (.I0(n51958), .I1(n53052), .I2(n59447), 
            .I3(n25207), .O(n14_adj_5527));
    defparam i6_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1482 (.I0(n52413), .I1(n53022), .I2(n57641), 
            .I3(\data_in_frame[16] [5]), .O(n9_adj_5528));
    defparam i1_4_lut_adj_1482.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1483 (.I0(n9_adj_5528), .I1(n14_adj_5527), .I2(n26738), 
            .I3(\data_in_frame[18] [0]), .O(n57830));
    defparam i7_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57628));
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1485 (.I0(n25266), .I1(n57628), .I2(n26061), 
            .I3(\data_in_frame[15] [7]), .O(n52094));
    defparam i3_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57767));
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5529), .S(n57178));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1487 (.I0(\data_out_frame[6] [6]), .I1(n57496), 
            .I2(GND_net), .I3(GND_net), .O(n26844));
    defparam i1_2_lut_adj_1487.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5530), .S(n57112));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5531), .S(n57120));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5532), .S(n57179));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5533), .S(n57180));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25][2] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5534), .S(n57181));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5535), .S(n57254));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1488 (.I0(n26721), .I1(\data_in_frame[12] [7]), 
            .I2(n25891), .I3(GND_net), .O(n58056));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1488.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1489 (.I0(\data_out_frame[13] [3]), .I1(n58105), 
            .I2(\data_out_frame[9] [1]), .I3(\data_out_frame[10] [7]), .O(n57700));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(n26069), .I1(n57657), .I2(GND_net), 
            .I3(GND_net), .O(n26061));
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1491 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57927));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1491.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1492 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n26487));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1492.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1493 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n57538));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1493.LUT_INIT = 16'h9696;
    SB_LUT4 i19_2_lut (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26380));   // verilog/coms.v(100[12:26])
    defparam i19_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5536), .S(n57253));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5537), .S(n57252));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1494 (.I0(\data_in_frame[11] [5]), .I1(n51992), 
            .I2(GND_net), .I3(GND_net), .O(n57899));
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1495 (.I0(n58072), .I1(n4_adj_5538), .I2(GND_net), 
            .I3(GND_net), .O(n57461));
    defparam i2_2_lut_adj_1495.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57924));
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5539), .S(n57251));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5540), .S(n57182));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1497 (.I0(n57461), .I1(n57924), .I2(\data_in_frame[10][2] ), 
            .I3(n25927), .O(n12_adj_5541));
    defparam i5_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1498 (.I0(n57927), .I1(\data_out_frame[15] [5]), 
            .I2(n1168), .I3(n57700), .O(n15_adj_5542));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1499 (.I0(n15_adj_5542), .I1(\data_out_frame[13] [4]), 
            .I2(n14_adj_5543), .I3(\data_out_frame[11] [1]), .O(n51946));   // verilog/coms.v(88[17:70])
    defparam i8_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(\data_out_frame[16] [0]), .I1(n51946), 
            .I2(GND_net), .I3(GND_net), .O(n51995));
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5544), .S(n57183));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1501 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[14] [1]), 
            .O(n62334));
    defparam i1_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5545), .S(n57184));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5546), .S(n57185));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5547), .S(n57110));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5548), .S(n57303));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5419), .S(n57304));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26][2] ), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5355), .S(n57305));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5351), .S(n57301));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5348), .S(n57306));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5347), .S(n57299));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5549), .S(n57307));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5346), .S(n57308));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5340), .S(n57309));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5339), .S(n57310));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27][2] ), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5335), .S(n57311));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5333), .S(n57302));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5332), .S(n57312));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5329), .S(n57300));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5328), .S(n57298));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1502 (.I0(n62334), .I1(n57921), .I2(\data_out_frame[14] [3]), 
            .I3(\data_out_frame[11] [1]), .O(n62342));
    defparam i1_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2873), .D(n1), .S(n28942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2873), .D(n5), 
            .S(n28941));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5326), .S(n57313));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5550), .S(n57100));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5551), .S(n57101));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5552), .S(n57102));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5553), .S(n57103));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5554), .S(n57104));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5555), .S(n57105));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5556), .S(n57098));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2873), .D(n26950), 
            .S(n28931));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1503 (.I0(n1699), .I1(n58102), .I2(n1563), .I3(n57681), 
            .O(n62344));
    defparam i1_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5322), .S(n57250));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1504 (.I0(n57933), .I1(n58108), .I2(n62344), 
            .I3(n62342), .O(n62352));
    defparam i1_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1505 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n57140));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1505.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1506 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n57141));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1506.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1507 (.I0(n26818), .I1(n62352), .I2(n57473), 
            .I3(n26104), .O(n62356));
    defparam i1_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1508 (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n40928));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1508.LUT_INIT = 16'hffdf;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5557), .S(n57099));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1509 (.I0(\data_in_frame[7] [6]), .I1(n12_adj_5541), 
            .I2(n58027), .I3(n25784), .O(n52028));
    defparam i6_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1510 (.I0(n52209), .I1(n52173), .I2(n26931), 
            .I3(n62356), .O(n62362));
    defparam i1_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1511 (.I0(n1720), .I1(n53030), .I2(n57672), .I3(n62362), 
            .O(n62368));
    defparam i1_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5321), .S(n57249));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1512 (.I0(n57924), .I1(n57568), .I2(\data_in_frame[10][3] ), 
            .I3(n57965), .O(n10_adj_5265));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5320), .S(n57248));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1513 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n57142));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1513.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1514 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n57143));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1514.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1515 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20]_c [0]), 
            .O(n57144));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1515.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1516 (.I0(n26721), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n58011));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1516.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1517 (.I0(n57528), .I1(n57891), .I2(n62292), 
            .I3(n57531), .O(n62298));
    defparam i1_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1518 (.I0(n62298), .I1(n60324), .I2(n57750), 
            .I3(n62368), .O(n57893));
    defparam i1_4_lut_adj_1518.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5318), .S(n57247));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29999));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1519 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20]_c [1]), 
            .O(n29019));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1519.LUT_INIT = 16'h4500;
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5307), .S(n57246));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1520 (.I0(\data_in_frame[3][1] ), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[7][5] ), .I3(n58099), .O(n10_adj_5558));
    defparam i4_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1521 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20]_c [2]), 
            .O(n57145));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1521.LUT_INIT = 16'h4500;
    SB_LUT4 i5_3_lut_adj_1522 (.I0(\data_in_frame[3][3] ), .I1(n10_adj_5558), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n52693));
    defparam i5_3_lut_adj_1522.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1523 (.I0(n51944), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[13] [5]), .I3(n25162), .O(n51960));
    defparam i1_2_lut_3_lut_4_lut_adj_1523.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1524 (.I0(n52693), .I1(n26853), .I2(n25927), 
            .I3(GND_net), .O(n57852));
    defparam i2_3_lut_adj_1524.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1525 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20][3] ), 
            .O(n29017));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1525.LUT_INIT = 16'h4500;
    SB_LUT4 i52901_4_lut (.I0(n26931), .I1(n26899), .I2(n53199), .I3(n62436), 
            .O(n68629));
    defparam i52901_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1526 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20]_c [4]), 
            .O(n57146));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1526.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1527 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20]_c [5]), 
            .O(n57147));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1527.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1528 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n57148));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1528.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1529 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57502));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1529.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1530 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58036));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1530.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57731));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1532 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n25769));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1532.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1533 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n57149));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1533.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1534 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21][0] ), 
            .O(n57150));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1534.LUT_INIT = 16'h4500;
    SB_LUT4 i4_4_lut_adj_1535 (.I0(n57731), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[4] [0]), .I3(n58036), .O(n10_adj_5559));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1536 (.I0(n25769), .I1(n10_adj_5559), .I2(\data_out_frame[5] [4]), 
            .I3(GND_net), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1536.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1537 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[7] [7]), 
            .I2(n6_adj_5560), .I3(n57580), .O(n4_adj_5538));
    defparam i1_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1538 (.I0(\data_in_frame[1] [5]), .I1(n4_adj_5538), 
            .I2(GND_net), .I3(GND_net), .O(n25906));
    defparam i2_2_lut_adj_1538.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1539 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[12] [3]), .I3(n25769), .O(n12_adj_5561));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25941));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1541 (.I0(n25751), .I1(n12_adj_5561), .I2(\data_out_frame[5] [3]), 
            .I3(\data_out_frame[8] [1]), .O(n26279));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1542 (.I0(n26279), .I1(n1516), .I2(\data_out_frame[12] [4]), 
            .I3(GND_net), .O(n1655));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1542.LUT_INIT = 16'h9696;
    SB_LUT4 add_1099_9_lut (.I0(n57097), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n49548), .O(n57098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1543 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6]_c [7]), 
            .I2(n25941), .I3(\data_in_frame[6] [4]), .O(n58144));
    defparam i3_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1544 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57577));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1544.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1545 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n29011));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1545.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1546 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n57151));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1546.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1547 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n58129));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1547.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1548 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21][3] ), 
            .O(n57152));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1548.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1549 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n57153));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1549.LUT_INIT = 16'h4500;
    SB_LUT4 i9_4_lut_adj_1550 (.I0(Kp_23__N_760), .I1(n57506), .I2(n57959), 
            .I3(n57446), .O(n22_adj_5562));   // verilog/coms.v(73[16:69])
    defparam i9_4_lut_adj_1550.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1551 (.I0(\data_in_frame[1] [0]), .I1(n57580), 
            .I2(n26373), .I3(Kp_23__N_772), .O(n21_adj_5563));   // verilog/coms.v(73[16:69])
    defparam i8_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1552 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[2] [4]), .I3(n14_adj_5564), .O(n23_adj_5565));   // verilog/coms.v(73[16:69])
    defparam i10_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1553 (.I0(n57666), .I1(\data_in_frame[5] [6]), 
            .I2(n57561), .I3(\data_in_frame[4] [4]), .O(n26_adj_5566));   // verilog/coms.v(73[16:69])
    defparam i11_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1554 (.I0(\data_in_frame[3] [5]), .I1(n23_adj_5565), 
            .I2(n21_adj_5563), .I3(n22_adj_5562), .O(n19_adj_5567));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1555 (.I0(\data_in_frame[4] [5]), .I1(n58014), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5568));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1555.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1556 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[3][3] ), 
            .I2(n57619), .I3(n57669), .O(n24_adj_5569));   // verilog/coms.v(73[16:69])
    defparam i9_4_lut_adj_1556.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1557 (.I0(n19_adj_5567), .I1(n26_adj_5566), .I2(\data_in_frame[4] [0]), 
            .I3(n57678), .O(n28_adj_5570));   // verilog/coms.v(73[16:69])
    defparam i13_4_lut_adj_1557.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1558 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n57154));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1558.LUT_INIT = 16'h4500;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[3]_c [7]), .I1(n28_adj_5570), 
            .I2(n24_adj_5569), .I3(n16_adj_5568), .O(n57822));   // verilog/coms.v(73[16:69])
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1559 (.I0(n57822), .I1(\data_in_frame[6] [0]), 
            .I2(Kp_23__N_799), .I3(n57648), .O(n58072));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1560 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n57155));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1560.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1561 (.I0(\data_in_frame[8] [0]), .I1(n57568), 
            .I2(\data_in_frame[3] [5]), .I3(n26428), .O(n25927));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1562 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4] [0]), 
            .I2(n25705), .I3(n25709), .O(n58126));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1563 (.I0(\data_out_frame[7] [7]), .I1(n57933), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n57452));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1563.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(n57694), .I1(n58027), .I2(GND_net), 
            .I3(GND_net), .O(n58028));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n58102));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1566 (.I0(n58102), .I1(n57452), .I2(\data_out_frame[12] [6]), 
            .I3(n58126), .O(n10_adj_5571));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1566.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1567 (.I0(n57918), .I1(n10_adj_5571), .I2(\data_out_frame[8] [2]), 
            .I3(GND_net), .O(n52130));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1567.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1568 (.I0(\data_out_frame[14] [5]), .I1(n1655), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n57528));
    defparam i2_3_lut_adj_1568.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26310));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1570 (.I0(n58024), .I1(n58042), .I2(n68629), 
            .I3(GND_net), .O(n57744));
    defparam i2_3_lut_adj_1570.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1571 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(n57528), .I3(n52130), .O(n57908));
    defparam i3_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1572 (.I0(\data_out_frame[15] [1]), .I1(n57750), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[17] [2]), 
            .O(n57574));
    defparam i3_4_lut_adj_1572.LUT_INIT = 16'h6996;
    SB_LUT4 i24049_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6]_c [7]), 
            .I2(n22792), .I3(GND_net), .O(n29719));
    defparam i24049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1573 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[3]_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5572));
    defparam i1_2_lut_adj_1573.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1574 (.I0(n52188), .I1(n57812), .I2(GND_net), 
            .I3(GND_net), .O(n58069));
    defparam i1_2_lut_adj_1574.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1575 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[4] [2]), .I3(n6_adj_5572), .O(n57519));
    defparam i4_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1576 (.I0(\data_out_frame[19][3] ), .I1(n57574), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5573));
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1577 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n57156));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1577.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1578 (.I0(\data_in_frame[5] [4]), .I1(n57725), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n25784));
    defparam i2_3_lut_adj_1578.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1579 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[3][0] ), 
            .I2(\data_in_frame[0] [6]), .I3(n35692), .O(n58014));
    defparam i3_4_lut_adj_1579.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1580 (.I0(\data_in_frame[3][2] ), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [0]), .O(n57725));
    defparam i1_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53871 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n69619));
    defparam byte_transmit_counter_0__bdd_4_lut_53871.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1581 (.I0(\data_in_frame[5] [2]), .I1(n58014), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5574));
    defparam i1_2_lut_adj_1581.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1582 (.I0(\data_out_frame[21] [4]), .I1(n26664), 
            .I2(n26896), .I3(n6_adj_5573), .O(n53093));
    defparam i4_4_lut_adj_1582.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1583 (.I0(\data_in_frame[7][4] ), .I1(n26231), 
            .I2(n57725), .I3(n6_adj_5574), .O(n57631));
    defparam i4_4_lut_adj_1583.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1584 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n57157));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1584.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1585 (.I0(\data_out_frame[21][3] ), .I1(n57908), 
            .I2(n57744), .I3(n26310), .O(n52390));
    defparam i3_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1586 (.I0(\data_in_frame[7] [6]), .I1(n57669), 
            .I2(GND_net), .I3(GND_net), .O(n24009));
    defparam i1_2_lut_adj_1586.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n57691));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1588 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n57158));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1588.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1589 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n57159));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1589.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1590 (.I0(\data_in_frame[3][6] ), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26428));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1590.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1591 (.I0(n26428), .I1(n57694), .I2(n57551), 
            .I3(\data_in_frame[1] [4]), .O(n26853));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1591.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1592 (.I0(\data_in_frame[6]_c [6]), .I1(\data_in_frame[7] [0]), 
            .I2(\data_in_frame[4] [6]), .I3(GND_net), .O(n57697));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1592.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1593 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22][3] ), 
            .O(n57160));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1593.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1594 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n57161));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1594.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1595 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(n35692), .I3(GND_net), .O(n26231));
    defparam i2_3_lut_adj_1595.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1596 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57873));
    defparam i1_2_lut_adj_1596.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1597 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[3][1] ), 
            .I2(\data_in_frame[5] [2]), .I3(GND_net), .O(n57678));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1597.LUT_INIT = 16'h9696;
    SB_LUT4 n69619_bdd_4_lut (.I0(n69619), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n69622));
    defparam n69619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1598 (.I0(\data_out_frame[21] [2]), .I1(n60087), 
            .I2(GND_net), .I3(GND_net), .O(n53176));
    defparam i1_2_lut_adj_1598.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53862 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n69613));
    defparam byte_transmit_counter_0__bdd_4_lut_53862.LUT_INIT = 16'he4aa;
    SB_LUT4 n69613_bdd_4_lut (.I0(n69613), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n69616));
    defparam n69613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1599 (.I0(n52011), .I1(\data_out_frame[23] [2]), 
            .I2(\data_out_frame[23][3] ), .I3(n53176), .O(n58136));
    defparam i1_2_lut_3_lut_4_lut_adj_1599.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1600 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n57162));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1600.LUT_INIT = 16'h4500;
    SB_LUT4 i24050_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6]_c [6]), 
            .I2(n22792), .I3(GND_net), .O(n29720));
    defparam i24050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_208_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n8_adj_5575), .I3(n57873), 
            .O(n3_adj_5548));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i4_4_lut_adj_1601 (.I0(n57580), .I1(n26690), .I2(n57678), 
            .I3(\data_in_frame[4] [7]), .O(n10_adj_5576));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1601.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1602 (.I0(n57959), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[5] [1]), .O(n14_adj_5577));
    defparam i6_4_lut_adj_1602.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1603 (.I0(\data_in_frame[7][2] ), .I1(n14_adj_5577), 
            .I2(n10_adj_5578), .I3(\data_in_frame[3][0] ), .O(n26496));
    defparam i7_4_lut_adj_1603.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1604 (.I0(n12_adj_5579), .I1(n57697), .I2(n26373), 
            .I3(n26370), .O(n26336));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1604.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1605 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n57163));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1605.LUT_INIT = 16'h4500;
    SB_LUT4 i52895_2_lut (.I0(n60278), .I1(\data_in_frame[7][3] ), .I2(GND_net), 
            .I3(GND_net), .O(n68623));   // verilog/coms.v(99[12:25])
    defparam i52895_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1606 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n57164));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1606.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1607 (.I0(\data_in_frame[8] [2]), .I1(n26853), 
            .I2(n25962), .I3(GND_net), .O(n3));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1607.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1608 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n57165));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1608.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1609 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n57166));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1609.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1610 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n57167));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1610.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1611 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n57293));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1611.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [7]), 
            .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5547));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1613 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n57292));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1613.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1614 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n57291));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1614.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1615 (.I0(\data_in_frame[4] [7]), .I1(n26367), 
            .I2(GND_net), .I3(GND_net), .O(n57666));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1615.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1616 (.I0(\data_in_frame[7][1] ), .I1(n58005), 
            .I2(n57666), .I3(\data_in_frame[4] [5]), .O(n26324));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1616.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_772));   // verilog/coms.v(81[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5546));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1617 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n57290));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1617.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1618 (.I0(\data_in_frame[6] [4]), .I1(n26401), 
            .I2(n57619), .I3(\data_in_frame[2] [0]), .O(n57596));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1619 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n57555));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1619.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1620 (.I0(\data_in_frame[8] [5]), .I1(n57596), 
            .I2(\data_in_frame[6] [3]), .I3(Kp_23__N_872), .O(n25891));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1620.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1621 (.I0(n26508), .I1(n57972), .I2(n57555), 
            .I3(Kp_23__N_974), .O(n13));   // verilog/coms.v(77[16:43])
    defparam i5_4_lut_adj_1621.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5545));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1622 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n57289));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1622.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5544));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1623 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n57288));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1623.LUT_INIT = 16'h4500;
    SB_LUT4 i7_4_lut_adj_1624 (.I0(n13), .I1(n11), .I2(n58028), .I3(n25927), 
            .O(n52555));   // verilog/coms.v(77[16:43])
    defparam i7_4_lut_adj_1624.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1625 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n57287));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1625.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1626 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n57286));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1626.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1627 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57446));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1627.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1628 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n57285));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1628.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1629 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n57284));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1629.LUT_INIT = 16'h4500;
    SB_LUT4 i24051_3_lut_4_lut (.I0(\Ki[14] ), .I1(\data_in_frame[4] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29806));
    defparam i24051_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_1630 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57551));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1630.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1631 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25953));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1631.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1632 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3][6] ), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(n57561));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1632.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1633 (.I0(\data_in_frame[1] [5]), .I1(n25953), 
            .I2(\data_in_frame[2] [0]), .I3(n6_adj_5580), .O(Kp_23__N_869));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1633.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1634 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n57283));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1634.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1635 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n57282));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1635.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5540));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1636 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n57281));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1636.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1637 (.I0(n25962), .I1(Kp_23__N_869), .I2(\data_in_frame[6] [2]), 
            .I3(\data_in_frame[8] [3]), .O(n4_c));   // verilog/coms.v(239[9:81])
    defparam i3_4_lut_adj_1637.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1638 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n57280));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1638.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1639 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n57279));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1639.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1640 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n57278));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1640.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1641 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n57277));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1641.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1642 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n57276));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1642.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1643 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n57275));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1643.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1644 (.I0(n25941), .I1(Kp_23__N_872), .I2(Kp_23__N_869), 
            .I3(\data_in_frame[8] [4]), .O(n25976));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1645 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n57274));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1645.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1646 (.I0(n25976), .I1(n4_c), .I2(\data_in_frame[10][5] ), 
            .I3(GND_net), .O(n26721));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1646.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1647 (.I0(\data_in_frame[11] [6]), .I1(Kp_23__N_760), 
            .I2(\data_in_frame[2] [6]), .I3(n57631), .O(n58114));
    defparam i1_2_lut_3_lut_4_lut_adj_1647.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1648 (.I0(n26069), .I1(n52034), .I2(GND_net), 
            .I3(GND_net), .O(n57675));
    defparam i1_2_lut_adj_1648.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1649 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n57273));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1649.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1650 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n57272));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1650.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1651 (.I0(\data_in_frame[10]_c [0]), .I1(\data_in_frame[9] [6]), 
            .I2(n68627), .I3(GND_net), .O(n25858));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1651.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1652 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n57271));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1652.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1653 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n57270));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1653.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1654 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n57269));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1654.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1655 (.I0(n25858), .I1(n57675), .I2(n52308), 
            .I3(n26721), .O(n59349));
    defparam i3_4_lut_adj_1655.LUT_INIT = 16'h6996;
    SB_LUT4 i46938_2_lut (.I0(PWMLimit[1]), .I1(PWMLimit[0]), .I2(GND_net), 
            .I3(GND_net), .O(n62656));
    defparam i46938_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1656 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n57268));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1656.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1657 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n57267));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1657.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1658 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n57266));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1658.LUT_INIT = 16'h4500;
    SB_LUT4 i8_4_lut_adj_1659 (.I0(\data_in_frame[7][3] ), .I1(n58056), 
            .I2(\data_in_frame[12] [2]), .I3(n57767), .O(n20_adj_5581));
    defparam i8_4_lut_adj_1659.LUT_INIT = 16'h6996;
    SB_LUT4 i6_2_lut (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5582));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1660 (.I0(n57756), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[11] [3]), .I3(n57852), .O(n19_adj_5583));
    defparam i7_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1661 (.I0(n57752), .I1(n60278), .I2(n59349), 
            .I3(GND_net), .O(n17_adj_5584));
    defparam i5_3_lut_adj_1661.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1662 (.I0(n17_adj_5584), .I1(n19_adj_5583), .I2(n18_adj_5582), 
            .I3(n20_adj_5581), .O(n58141));
    defparam i11_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1663 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n58077));
    defparam i1_2_lut_adj_1663.LUT_INIT = 16'h6666;
    SB_LUT4 i23253_4_lut (.I0(n62656), .I1(n35), .I2(n379), .I3(n380), 
            .O(n4_adj_14));
    defparam i23253_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i6_4_lut_adj_1664 (.I0(n58141), .I1(n52194), .I2(n26304), 
            .I3(n58117), .O(n15_adj_5586));
    defparam i6_4_lut_adj_1664.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1665 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n57265));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1665.LUT_INIT = 16'h4500;
    SB_LUT4 i8_4_lut_adj_1666 (.I0(n15_adj_5586), .I1(n57899), .I2(n14_adj_5587), 
            .I3(n24005), .O(n25266));
    defparam i8_4_lut_adj_1666.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1667 (.I0(\data_out_frame[20]_c [2]), 
            .I1(n52042), .I2(n23735), .I3(\data_out_frame[20][3] ), .O(n52236));
    defparam i1_2_lut_3_lut_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1668 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n57264));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1668.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1669 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n57263));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1669.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25][2] ), 
            .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1671 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n57262));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1671.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5533));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1672 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n57261));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1672.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1673 (.I0(n26517), .I1(n26487), .I2(\data_in_frame[13] [2]), 
            .I3(\data_in_frame[13] [5]), .O(n57761));
    defparam i3_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1674 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[0][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5588));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1674.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1675 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[4] [4]), .I3(n6_adj_5588), .O(n57513));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1675.LUT_INIT = 16'h6996;
    SB_LUT4 i23276_3_lut_4_lut (.I0(deadband[0]), .I1(\data_in_frame[16] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29529));
    defparam i23276_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_777_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1676 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n57260));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1676.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5531));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1677 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n57259));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1677.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1678 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n57258));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1678.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1679 (.I0(\data_in_frame[4] [4]), .I1(n25842), 
            .I2(n26401), .I3(GND_net), .O(n26370));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1679.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1680 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n57257));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1680.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1681 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26304));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1681.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1682 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25745));
    defparam i1_2_lut_adj_1682.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [6]), 
            .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5530));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1684 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n57256));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1684.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1054_i24_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i24_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1685 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n57255));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1685.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1686 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23][3] ), 
            .O(n57168));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1686.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1054_i23_3_lut_4_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i23_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1687 (.I0(\data_in_frame[4] [5]), .I1(n57663), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_993));
    defparam i1_2_lut_adj_1687.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_194_i2_4_lut (.I0(\data_out_frame[24][2] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1688 (.I0(\data_in_frame[11] [1]), .I1(n52555), 
            .I2(\data_in_frame[10][7] ), .I3(n52308), .O(n57752));
    defparam i3_4_lut_adj_1688.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1689 (.I0(\data_in_frame[9] [3]), .I1(n57593), 
            .I2(\data_in_frame[9] [6]), .I3(n25745), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1689.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1690 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57911));
    defparam i1_2_lut_adj_1690.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1691 (.I0(n57761), .I1(n52001), .I2(n52194), 
            .I3(GND_net), .O(n59598));
    defparam i2_3_lut_adj_1691.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1692 (.I0(Kp_23__N_1080), .I1(n57752), .I2(n7_adj_5589), 
            .I3(GND_net), .O(n52107));
    defparam i2_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1054_i22_3_lut_4_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i22_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_adj_1693 (.I0(\data_in_frame[13] [7]), .I1(n52094), 
            .I2(GND_net), .I3(GND_net), .O(n57443));
    defparam i1_2_lut_adj_1693.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1054_i21_3_lut_4_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i21_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1694 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n57169));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1694.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1054_i20_3_lut_4_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i20_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1054_i19_3_lut_4_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i19_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1695 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n57170));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1695.LUT_INIT = 16'h4500;
    SB_LUT4 i47331_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63059));
    defparam i47331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47332_4_lut (.I0(n63059), .I1(n28205), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1] [5]), .O(n63060));
    defparam i47332_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 mux_1054_i18_3_lut_4_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i18_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i52899_2_lut_3_lut_4_lut (.I0(n24005), .I1(\data_in_frame[7] [6]), 
            .I2(n57669), .I3(\data_in_frame[9] [7]), .O(n68627));   // verilog/coms.v(99[12:25])
    defparam i52899_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i47330_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63058));
    defparam i47330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i17_3_lut_4_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[16]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i17_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1696 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n57171));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1696.LUT_INIT = 16'h4500;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [5]), 
            .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1698 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n57172));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1698.LUT_INIT = 16'h4500;
    SB_LUT4 i4_4_lut_adj_1699 (.I0(n52107), .I1(n59598), .I2(n57911), 
            .I3(n6_adj_5327), .O(n53022));
    defparam i4_4_lut_adj_1699.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53857 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n69607));
    defparam byte_transmit_counter_0__bdd_4_lut_53857.LUT_INIT = 16'he4aa;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1054_i16_3_lut_4_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i16_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1700 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n57173));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1700.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_adj_1701 (.I0(\data_in_frame[18] [1]), .I1(n53022), 
            .I2(GND_net), .I3(GND_net), .O(n57525));
    defparam i1_2_lut_adj_1701.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1702 (.I0(n60454), .I1(n58021), .I2(n57685), 
            .I3(n6_adj_5590), .O(n57809));
    defparam i4_4_lut_adj_1702.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [4]), 
            .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1704 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n57174));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1704.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_187_i2_4_lut (.I0(\data_out_frame[23][3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1705 (.I0(\data_in_frame[20] [1]), .I1(\data_in_frame[22] [3]), 
            .I2(n57809), .I3(n57525), .O(n10_adj_5591));
    defparam i4_4_lut_adj_1705.LUT_INIT = 16'h6996;
    SB_LUT4 i46958_4_lut (.I0(n22911), .I1(\data_in_frame[19]_c [7]), .I2(n10_adj_5591), 
            .I3(n57830), .O(n62676));
    defparam i46958_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1706 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24][2] ), 
            .O(n57175));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1706.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut_adj_1707 (.I0(n51954), .I1(\data_in_frame[20] [5]), 
            .I2(n52147), .I3(n57792), .O(n8_adj_5592));
    defparam i3_4_lut_adj_1707.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1708 (.I0(\data_in_frame[23] [5]), .I1(n57564), 
            .I2(n57615), .I3(GND_net), .O(n52504));
    defparam i1_3_lut_adj_1708.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1709 (.I0(\data_in_frame[19] [5]), .I1(n59240), 
            .I2(n59871), .I3(n59287), .O(n53032));
    defparam i2_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 i52096_3_lut (.I0(n69610), .I1(n69568), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n67824));
    defparam i52096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_adj_1710 (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[18] [2]), 
            .I2(n57809), .I3(GND_net), .O(n8_adj_5593));
    defparam i3_3_lut_adj_1710.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1711 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n57176));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1711.LUT_INIT = 16'h4500;
    SB_LUT4 i14072_3_lut (.I0(\data_out_frame[1] [6]), .I1(\data_out_frame[3] [6]), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28147));   // verilog/coms.v(109[34:55])
    defparam i14072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47322_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63050));
    defparam i47322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1712 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n57177));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1712.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1054_i15_3_lut_4_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i15_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i14_3_lut_4_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i14_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1713 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n57178));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1713.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_1714 (.I0(n52036), .I1(n57792), .I2(\data_in_frame[23] [1]), 
            .I3(GND_net), .O(n59453));
    defparam i2_3_lut_adj_1714.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1715 (.I0(n52036), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[23] [3]), .I3(n57634), .O(n60320));
    defparam i2_4_lut_adj_1715.LUT_INIT = 16'h6996;
    SB_LUT4 i1_rep_204_2_lut (.I0(\data_in_frame[20] [1]), .I1(\data_in_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n70027));
    defparam i1_rep_204_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1716 (.I0(\data_in_frame[17] [6]), .I1(n70027), 
            .I2(n25808), .I3(\data_in_frame[22] [2]), .O(n12_adj_5594));
    defparam i5_4_lut_adj_1716.LUT_INIT = 16'h6996;
    SB_LUT4 i47323_4_lut (.I0(n63050), .I1(n28147), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63051));
    defparam i47323_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i4_4_lut_adj_1717 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[22] [0]), .I3(\data_in_frame[21] [6]), .O(n10_adj_5595));
    defparam i4_4_lut_adj_1717.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1718 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[23] [2]), 
            .I2(n52147), .I3(GND_net), .O(n60373));
    defparam i2_3_lut_adj_1718.LUT_INIT = 16'h9696;
    SB_LUT4 i47321_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63049));
    defparam i47321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1719 (.I0(\data_in_frame[20] [0]), .I1(n12_adj_5594), 
            .I2(n57830), .I3(n59287), .O(n59724));
    defparam i6_4_lut_adj_1719.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1720 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n57112));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1720.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1721 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n57120));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1721.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1054_i13_3_lut_4_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i13_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i46964_4_lut (.I0(\data_in_frame[22] [6]), .I1(n62676), .I2(n57816), 
            .I3(\data_in_frame[20] [4]), .O(n62682));
    defparam i46964_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1722 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n57179));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1722.LUT_INIT = 16'h4500;
    SB_LUT4 i7_4_lut_adj_1723 (.I0(\data_in_frame[22] [7]), .I1(n52504), 
            .I2(n8_adj_5592), .I3(n58061), .O(n24_adj_5596));
    defparam i7_4_lut_adj_1723.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19][3] ), 
            .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'ha088;
    SB_LUT4 i46966_4_lut (.I0(n57615), .I1(n59724), .I2(n57984), .I3(\data_in_frame[23] [6]), 
            .O(n62684));
    defparam i46966_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1725 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n57180));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1725.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1726 (.I0(n60373), .I1(Kp_23__N_1551), .I2(n10_adj_5595), 
            .I3(n59871), .O(n23_adj_5597));
    defparam i6_4_lut_adj_1726.LUT_INIT = 16'h2882;
    SB_LUT4 i3_3_lut_adj_1727 (.I0(\data_in_frame[22] [1]), .I1(\data_in_frame[17] [6]), 
            .I2(n57956), .I3(GND_net), .O(n8_adj_5598));
    defparam i3_3_lut_adj_1727.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1728 (.I0(n57564), .I1(n57634), .I2(\data_in_frame[23] [4]), 
            .I3(GND_net), .O(n60421));
    defparam i2_3_lut_adj_1728.LUT_INIT = 16'h9696;
    SB_LUT4 i47414_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63142));
    defparam i47414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1729 (.I0(\data_in_frame[23] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(n53032), .I3(n57984), .O(n59645));
    defparam i2_4_lut_adj_1729.LUT_INIT = 16'h6996;
    SB_LUT4 i47415_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63143));
    defparam i47415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47412_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63140));
    defparam i47412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i12_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i12_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1730 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25][2] ), 
            .O(n57181));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1730.LUT_INIT = 16'h4500;
    SB_LUT4 i47411_3_lut (.I0(\data_out_frame[20]_c [0]), .I1(\data_out_frame[21][0] ), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63139));
    defparam i47411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i11_3_lut_4_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i11_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_3_lut_adj_1731 (.I0(\data_out_frame[19] [6]), .I1(n52663), 
            .I2(\data_out_frame[22] [0]), .I3(GND_net), .O(n53137));
    defparam i1_2_lut_3_lut_adj_1731.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1732 (.I0(\data_in_frame[21] [7]), .I1(n60421), 
            .I2(n8_adj_5598), .I3(n57541), .O(n19_adj_5599));
    defparam i2_4_lut_adj_1732.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1733 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n57254));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1733.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47285_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63013));
    defparam i47285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1734 (.I0(n59679), .I1(n59453), .I2(n8_adj_5593), 
            .I3(\data_in_frame[22] [4]), .O(n22_adj_5600));
    defparam i5_4_lut_adj_1734.LUT_INIT = 16'h1221;
    SB_LUT4 mux_1054_i10_3_lut_4_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i10_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i46968_4_lut (.I0(\data_in_frame[23] [0]), .I1(n60320), .I2(n52147), 
            .I3(n57792), .O(n62686));
    defparam i46968_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i15_4_lut_adj_1735 (.I0(n23_adj_5597), .I1(n62684), .I2(n24_adj_5596), 
            .I3(n62682), .O(n32_adj_5601));
    defparam i15_4_lut_adj_1735.LUT_INIT = 16'h0020;
    SB_LUT4 i10_4_lut_adj_1736 (.I0(n19_adj_5599), .I1(n59645), .I2(\data_in_frame[22] [5]), 
            .I3(n57706), .O(n27_c));
    defparam i10_4_lut_adj_1736.LUT_INIT = 16'h2002;
    SB_LUT4 i16_4_lut (.I0(n27_c), .I1(n32_adj_5601), .I2(n62686), .I3(n22_adj_5600), 
            .O(n33793));
    defparam i16_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i47286_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63014));
    defparam i47286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47289_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63017));
    defparam i47289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47288_3_lut (.I0(\data_out_frame[20]_c [1]), .I1(\data_out_frame[21] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63016));
    defparam i47288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i9_3_lut_4_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i9_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1737 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n57253));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1737.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5484));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i21833_3_lut_4_lut (.I0(\data_in_frame[19]_c [7]), .I1(\data_in_frame[3]_c [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[7]));
    defparam i21833_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1738 (.I0(\data_out_frame[19] [6]), .I1(n52663), 
            .I2(\data_out_frame[17] [6]), .I3(GND_net), .O(n6_adj_5403));
    defparam i1_2_lut_3_lut_adj_1738.LUT_INIT = 16'h9696;
    SB_LUT4 i47423_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63151));
    defparam i47423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1739 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n57252));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1739.LUT_INIT = 16'h4500;
    SB_LUT4 i47424_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63152));
    defparam i47424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47268_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62996));
    defparam i47268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5482));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1054_i7_3_lut_4_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3][6] ), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i7_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i47267_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62995));
    defparam i47267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i6_3_lut_4_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i6_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5481));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47399_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63127));
    defparam i47399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1740 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n57251));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1740.LUT_INIT = 16'h4500;
    SB_LUT4 i47400_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63128));
    defparam i47400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5480));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1741 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n57182));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1741.LUT_INIT = 16'h4500;
    SB_LUT4 i47274_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63002));
    defparam i47274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i5_3_lut_4_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3][4] ), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i5_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1742 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n57183));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1742.LUT_INIT = 16'h4500;
    SB_LUT4 i47273_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63001));
    defparam i47273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50571_2_lut (.I0(n69616), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65734));
    defparam i50571_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1743 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n57184));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1743.LUT_INIT = 16'h4500;
    SB_LUT4 i14070_3_lut (.I0(\data_out_frame[1] [7]), .I1(\data_out_frame[3] [7]), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28145));   // verilog/coms.v(109[34:55])
    defparam i14070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1744 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(n57631), .O(n24005));
    defparam i1_2_lut_3_lut_4_lut_adj_1744.LUT_INIT = 16'h6996;
    SB_LUT4 i47316_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63044));
    defparam i47316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5479));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47317_4_lut (.I0(n63044), .I1(n28145), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63045));
    defparam i47317_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 mux_1054_i4_3_lut_4_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3][3] ), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i4_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1745 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n57185));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1745.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1746 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n57110));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1746.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1747 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n57250));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1747.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1054_i3_3_lut_4_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3][2] ), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i3_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i47315_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63043));
    defparam i47315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i2_3_lut_4_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3][1] ), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i2_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5478));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1748 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n57249));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1748.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1749 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n57248));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1749.LUT_INIT = 16'h4500;
    SB_LUT4 select_777_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i50376_2_lut (.I0(n69622), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65735));
    defparam i50376_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1750 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n57247));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1750.LUT_INIT = 16'h4500;
    SB_LUT4 i47387_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63115));
    defparam i47387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1751 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n57246));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1751.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_4_lut_adj_1752 (.I0(n1954), .I1(n1951), .I2(n1957), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n59892));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1752.LUT_INIT = 16'h8000;
    SB_LUT4 select_777_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47388_3_lut (.I0(\data_out_frame[18][4] ), .I1(\data_out_frame[19] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63116));
    defparam i47388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47337_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63065));
    defparam i47337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47336_3_lut (.I0(\data_out_frame[20]_c [4]), .I1(\data_out_frame[21] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63064));
    defparam i47336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1753 (.I0(n25842), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0][2] ), .I3(\data_in_frame[0][1] ), .O(Kp_23__N_799));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1753.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1754 (.I0(\data_in_frame[6]_c [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[0][3] ), .O(n12_adj_5579));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1754.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1755 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(n12_adj_5579), .O(n58005));
    defparam i1_2_lut_3_lut_4_lut_adj_1755.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1756 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(n25621), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_5602));
    defparam i1_3_lut_4_lut_adj_1756.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_3_lut_4_lut_adj_1757 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3545[0]), .I3(n43569), .O(n25545));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1757.LUT_INIT = 16'ha8aa;
    SB_LUT4 i6_4_lut_adj_1758 (.I0(n57822), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[3][6] ), .I3(n57648), .O(n15_adj_5603));
    defparam i6_4_lut_adj_1758.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1759 (.I0(n15_adj_5603), .I1(n26373), .I2(n14_adj_5604), 
            .I3(\data_in_frame[3] [5]), .O(n59699));
    defparam i8_4_lut_adj_1759.LUT_INIT = 16'h6996;
    SB_LUT4 i14080_3_lut (.I0(\data_out_frame[1] [1]), .I1(\data_out_frame[3] [1]), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28155));   // verilog/coms.v(109[34:55])
    defparam i14080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1054_i1_3_lut_4_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3][0] ), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n4762[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i1_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i47095_4_lut (.I0(n59699), .I1(Kp_23__N_974), .I2(n4_c), .I3(\data_in_frame[8] [6]), 
            .O(n62814));
    defparam i47095_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1760 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0][2] ), 
            .I2(\data_in_frame[0][1] ), .I3(n57513), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1760.LUT_INIT = 16'h6996;
    SB_LUT4 i47346_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63074));
    defparam i47346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'ha088;
    SB_LUT4 i47125_4_lut (.I0(n22911), .I1(n62814), .I2(n58028), .I3(\data_in_frame[8] [0]), 
            .O(n62844));
    defparam i47125_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i11_4_lut_adj_1762 (.I0(n24005), .I1(n57461), .I2(n24009), 
            .I3(n26324), .O(n28_adj_5605));
    defparam i11_4_lut_adj_1762.LUT_INIT = 16'h0080;
    SB_LUT4 i47347_4_lut (.I0(n63074), .I1(n28155), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n63075));
    defparam i47347_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 select_777_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47345_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63073));
    defparam i47345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_148_i2_4_lut (.I0(\data_out_frame[18][4] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18][3] ), 
            .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[1] [3]), .I1(n25842), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[5] [7]), .O(n14_adj_5604));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51539_4_lut (.I0(n69538), .I1(n69526), .I2(byte_transmit_counter[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n67267));
    defparam i51539_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_777_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47266_3_lut (.I0(n69556), .I1(n67267), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i47266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47093_4_lut (.I0(n25891), .I1(n25976), .I2(n26336), .I3(n3), 
            .O(n62812));
    defparam i47093_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51691_4_lut (.I0(n69502), .I1(n69550), .I2(byte_transmit_counter[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n67419));
    defparam i51691_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i47194_3_lut (.I0(n69544), .I1(n67419), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[4]));
    defparam i47194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50559_2_lut (.I0(n69532), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65732));
    defparam i50559_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i10_4_lut_adj_1764 (.I0(n26496), .I1(n52693), .I2(n7_adj_5589), 
            .I3(n68623), .O(n27_adj_5606));
    defparam i10_4_lut_adj_1764.LUT_INIT = 16'h0001;
    SB_LUT4 i16_4_lut_adj_1765 (.I0(n27_adj_5606), .I1(n62812), .I2(n28_adj_5605), 
            .I3(n62844), .O(n33801));
    defparam i16_4_lut_adj_1765.LUT_INIT = 16'h0020;
    SB_LUT4 i47294_4_lut (.I0(\data_out_frame[0] [4]), .I1(\data_out_frame[3] [4]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n63022));
    defparam i47294_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0] [3]), 
            .I1(\data_out_frame[1] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5607));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47300_4_lut (.I0(n1_adj_5607), .I1(\data_out_frame[3] [3]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n63028));
    defparam i47300_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i47435_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63163));
    defparam i47435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(n51960), .I3(GND_net), .O(n7_adj_5365));   // verilog/coms.v(79[16:43])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i47436_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63164));
    defparam i47436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47277_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63005));
    defparam i47277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6691_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1951), 
            .I2(n59374), .I3(n4452), .O(n20437));   // verilog/coms.v(148[4] 304[11])
    defparam i6691_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n20437), .I1(n1951), .I2(n22769), .I3(n4_adj_5338), 
            .O(n27049));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hbbba;
    SB_LUT4 i47276_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63004));
    defparam i47276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i456_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2060));   // verilog/coms.v(148[4] 304[11])
    defparam i456_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47282_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63010));
    defparam i47282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1767 (.I0(Kp_23__N_1748), .I1(n33793), .I2(GND_net), 
            .I3(GND_net), .O(n27726));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1767.LUT_INIT = 16'h8888;
    SB_LUT4 i47283_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63011));
    defparam i47283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47292_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63020));
    defparam i47292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47291_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63019));
    defparam i47291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1768 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[17] [6]), .I3(GND_net), .O(n6_adj_5590));
    defparam i1_2_lut_3_lut_adj_1768.LUT_INIT = 16'h9696;
    SB_LUT4 i19732_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(n33801), .I3(n33793), .O(n27767));   // verilog/coms.v(18[27:29])
    defparam i19732_4_lut.LUT_INIT = 16'he420;
    SB_LUT4 i46883_4_lut (.I0(n1951), .I1(n1954), .I2(n3303), .I3(n1957), 
            .O(n62601));   // verilog/coms.v(139[4] 141[7])
    defparam i46883_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1954), 
            .I2(n62601), .I3(n60102), .O(n56292));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hb3a0;
    SB_LUT4 i2_2_lut_3_lut_adj_1770 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[4] [5]), 
            .I2(n57663), .I3(GND_net), .O(n7_adj_5589));
    defparam i2_2_lut_3_lut_adj_1770.LUT_INIT = 16'h9696;
    SB_LUT4 i14130_2_lut (.I0(\byte_transmit_counter[1] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n28205));   // verilog/coms.v(109[34:55])
    defparam i14130_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 select_777_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6696_4_lut (.I0(n1955), .I1(\FRAME_MATCHER.state [3]), .I2(n1957), 
            .I3(n25545), .O(n20442));   // verilog/coms.v(148[4] 304[11])
    defparam i6696_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i445_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2049));   // verilog/coms.v(148[4] 304[11])
    defparam i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1771 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [7]), .I3(GND_net), .O(n57593));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1771.LUT_INIT = 16'h9696;
    SB_LUT4 i47325_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63053));
    defparam i47325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47326_4_lut (.I0(n63053), .I1(n28205), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1] [0]), .O(n63054));
    defparam i47326_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i444_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2048));   // verilog/coms.v(148[4] 304[11])
    defparam i444_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47324_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63052));
    defparam i47324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1772 (.I0(\data_out_frame[20]_c [4]), 
            .I1(n51970), .I2(n52973), .I3(n57905), .O(n53119));
    defparam i1_2_lut_3_lut_4_lut_adj_1772.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1773 (.I0(\data_out_frame[20]_c [4]), 
            .I1(n51970), .I2(n52973), .I3(\data_out_frame[22] [5]), .O(n57805));
    defparam i1_2_lut_3_lut_4_lut_adj_1773.LUT_INIT = 16'h9669;
    SB_LUT4 i28972_4_lut (.I0(n5_adj_5602), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i[3] ), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i28972_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_3_lut_adj_1774 (.I0(n26324), .I1(\data_in_frame[11] [5]), 
            .I2(n51992), .I3(GND_net), .O(n52194));
    defparam i1_2_lut_3_lut_adj_1774.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1775 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[11] [6]), .O(n14_adj_5587));
    defparam i5_3_lut_4_lut_adj_1775.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1776 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3][6] ), .I3(\data_in_frame[1] [4]), .O(n6_adj_5580));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1776.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1777 (.I0(\FRAME_MATCHER.i[4] ), .I1(n25621), .I2(GND_net), 
            .I3(GND_net), .O(n25468));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1777.LUT_INIT = 16'heeee;
    SB_LUT4 i28974_4_lut (.I0(n8_adj_15), .I1(\FRAME_MATCHER.i [31]), .I2(n25468), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i28974_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut_adj_1778 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n22769));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1778.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_4_lut_adj_1779 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[3]_c [7]), .I3(\data_in_frame[6] [1]), .O(n57965));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1779.LUT_INIT = 16'h6996;
    SB_LUT4 i50951_2_lut (.I0(n69634), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65787));
    defparam i50951_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_2_lut (.I0(n25545), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27626));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1780 (.I0(n24005), .I1(\data_in_frame[7] [6]), 
            .I2(n57669), .I3(GND_net), .O(n26508));
    defparam i1_2_lut_3_lut_adj_1780.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1781 (.I0(n4452), .I1(n27626), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n22769), .O(n59773));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1781.LUT_INIT = 16'hffdc;
    SB_LUT4 i2_3_lut_4_lut_adj_1782 (.I0(n26373), .I1(n57513), .I2(n57596), 
            .I3(\data_in_frame[6] [5]), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1782.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1783 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [6]), .O(n57619));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1783.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_139_i2_4_lut (.I0(\data_out_frame[17][3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n25550), .I1(n1957), .I2(n1955), .I3(n59773), 
            .O(n27046));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hbaaa;
    SB_LUT4 i47390_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63118));
    defparam i47390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1785 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n57396), .I3(LED_c), .O(n27315));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1785.LUT_INIT = 16'hfe00;
    SB_LUT4 i2_2_lut_adj_1786 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5609));
    defparam i2_2_lut_adj_1786.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1787 (.I0(\data_in_frame[5] [0]), .I1(n25842), 
            .I2(\data_in_frame[2] [3]), .I3(n57728), .O(n26367));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1787.LUT_INIT = 16'h6996;
    SB_LUT4 i47391_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63119));
    defparam i47391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1788 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5610));
    defparam i6_4_lut_adj_1788.LUT_INIT = 16'hfeff;
    SB_LUT4 select_777_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1789 (.I0(\data_in[3] [6]), .I1(n14_adj_5610), 
            .I2(n10_adj_5609), .I3(\data_in[2] [1]), .O(n25618));
    defparam i7_4_lut_adj_1789.LUT_INIT = 16'hfffd;
    SB_LUT4 i47310_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63038));
    defparam i47310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1790 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n25618), .I3(\data_in[0] [5]), .O(n20_adj_5611));
    defparam i8_4_lut_adj_1790.LUT_INIT = 16'hfbff;
    SB_LUT4 i47309_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63037));
    defparam i47309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47393_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63121));
    defparam i47393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1791 (.I0(n25492), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_5612));
    defparam i7_4_lut_adj_1791.LUT_INIT = 16'hfeff;
    SB_LUT4 i47083_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [3]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n62802));
    defparam i47083_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i47394_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63122));
    defparam i47394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_adj_1792 (.I0(n62802), .I1(n19_adj_5612), .I2(n20_adj_5611), 
            .I3(GND_net), .O(n1951));
    defparam i11_3_lut_adj_1792.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1793 (.I0(\data_in[2] [4]), .I1(n25618), .I2(\data_in[1] [5]), 
            .I3(n25676), .O(n18_adj_5613));
    defparam i7_4_lut_adj_1793.LUT_INIT = 16'hfffd;
    SB_LUT4 i47298_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63026));
    defparam i47298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1794 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3470));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1794.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut_adj_1795 (.I0(\data_in[0] [6]), .I1(n18_adj_5613), 
            .I2(\data_in[3] [0]), .I3(n25572), .O(n20_adj_5614));
    defparam i9_4_lut_adj_1795.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5615));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 select_777_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1796 (.I0(\data_in_frame[0] [4]), .I1(n57506), 
            .I2(n10_adj_5576), .I3(n58099), .O(n60278));   // verilog/coms.v(73[16:69])
    defparam i5_3_lut_4_lut_adj_1796.LUT_INIT = 16'h6996;
    SB_LUT4 i47297_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63025));
    defparam i47297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1797 (.I0(n15_adj_5615), .I1(n20_adj_5614), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1954));
    defparam i10_4_lut_adj_1797.LUT_INIT = 16'hfeff;
    SB_LUT4 select_777_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1798 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n33795));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1798.LUT_INIT = 16'heeee;
    SB_LUT4 i47189_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62917));
    defparam i47189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1799 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5616));
    defparam i4_4_lut_adj_1799.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1800 (.I0(\data_in[3] [4]), .I1(n10_adj_5616), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n25676));
    defparam i5_3_lut_adj_1800.LUT_INIT = 16'hdfdf;
    SB_LUT4 i47190_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62918));
    defparam i47190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1801 (.I0(\data_in[1] [0]), .I1(\data_in[2] [4]), 
            .I2(\data_in[3] [0]), .I3(GND_net), .O(n14_adj_5617));
    defparam i5_3_lut_adj_1801.LUT_INIT = 16'hdfdf;
    SB_LUT4 i47445_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63173));
    defparam i47445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1802 (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), 
            .I2(n25676), .I3(\data_in[1] [5]), .O(n15_adj_5618));
    defparam i6_4_lut_adj_1802.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1803 (.I0(n15_adj_5618), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5617), .I3(\data_in[0] [3]), .O(n25492));
    defparam i8_4_lut_adj_1803.LUT_INIT = 16'hfbff;
    SB_LUT4 i47444_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n63172));
    defparam i47444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1804 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5619));
    defparam i6_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1805 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_5620));
    defparam i7_4_lut_adj_1805.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1806 (.I0(n17_adj_5620), .I1(\data_in[1] [6]), 
            .I2(n16_adj_5619), .I3(\data_in[3] [7]), .O(n25572));
    defparam i9_4_lut_adj_1806.LUT_INIT = 16'hfbff;
    SB_LUT4 i3_4_lut_adj_1807 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[2] [3]), .I3(\data_in[3] [1]), .O(n60447));
    defparam i3_4_lut_adj_1807.LUT_INIT = 16'h8000;
    SB_LUT4 i3_3_lut_4_lut_adj_1808 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[21] [2]), 
            .I2(n60087), .I3(n58090), .O(n8_adj_5575));
    defparam i3_3_lut_4_lut_adj_1808.LUT_INIT = 16'h6996;
    SB_LUT4 i23275_3_lut_4_lut (.I0(n380), .I1(n460), .I2(n459), .I3(n379), 
            .O(n4_adj_16));
    defparam i23275_3_lut_4_lut.LUT_INIT = 16'h40f4;
    SB_LUT4 select_777_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1809 (.I0(\data_in[0] [7]), .I1(n25572), .I2(n25492), 
            .I3(n60447), .O(n12_adj_5622));
    defparam i5_4_lut_adj_1809.LUT_INIT = 16'hfeff;
    SB_LUT4 select_777_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18_4_lut_adj_1810 (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [20]), .I3(\FRAME_MATCHER.i [18]), .O(n44));
    defparam i18_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1811 (.I0(\data_in[3] [3]), .I1(n12_adj_5622), 
            .I2(\data_in[3] [6]), .I3(\data_in[2] [1]), .O(n1957));
    defparam i6_4_lut_adj_1811.LUT_INIT = 16'hfdff;
    SB_LUT4 i362_2_lut (.I0(n1954), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n1955));   // verilog/coms.v(142[4] 144[7])
    defparam i362_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1812 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(n62562), .I3(n57599), .O(n62566));   // verilog/coms.v(79[16:43])
    defparam i1_3_lut_4_lut_adj_1812.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1813 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [9]), .O(n42));
    defparam i16_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1814 (.I0(n43569), .I1(n59892), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(n42760), .O(n6_adj_5623));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1814.LUT_INIT = 16'hccec;
    SB_LUT4 i3_4_lut_adj_1815 (.I0(n33795), .I1(n6_adj_5623), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n69866));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1815.LUT_INIT = 16'hefee;
    SB_LUT4 i17_4_lut_adj_1816 (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [16]), .O(n43_adj_5624));
    defparam i17_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1817 (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [19]), .I3(\FRAME_MATCHER.i [8]), .O(n41));
    defparam i15_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_4_lut_adj_1818 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[16] [1]), .I3(n10_adj_5363), .O(n52973));
    defparam i5_3_lut_4_lut_adj_1818.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1819 (.I0(n52390), .I1(n53093), .I2(n52188), 
            .I3(n57812), .O(n58090));
    defparam i1_3_lut_4_lut_adj_1819.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14_4_lut_adj_1820 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [26]), .O(n40));
    defparam i14_4_lut_adj_1820.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1821 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(n35692), .I3(n57914), .O(n58099));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_4_lut_adj_1821.LUT_INIT = 16'h6996;
    SB_LUT4 i13_2_lut_adj_1822 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut_adj_1822.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43_adj_5624), .I2(n42), .I3(n44), 
            .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1823 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[18] [5]), .I3(\data_out_frame[14] [4]), 
            .O(n60035));
    defparam i2_3_lut_4_lut_adj_1823.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n57303));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h5100;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [29]), 
            .I2(\FRAME_MATCHER.i [17]), .I3(\FRAME_MATCHER.i [24]), .O(n45_adj_5625));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 select_777_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1825 (.I0(\data_in_frame[1] [5]), .I1(n4_adj_5538), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[1] [3]), .O(n57568));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1825.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n57304));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26][2] ), 
            .O(n57305));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1828 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n25709));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1828.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_131_i2_4_lut (.I0(\data_out_frame[16][3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1829 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n25751));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1829.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(n45_adj_5625), .I1(n50), .I2(n39), .I3(n40), 
            .O(n25621));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28975_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25621), .I3(\FRAME_MATCHER.i[4] ), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i28975_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i464_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2068));   // verilog/coms.v(148[4] 304[11])
    defparam i464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1830 (.I0(\data_out_frame[16][3] ), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n58024));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1830.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1831 (.I0(n57722), .I1(\data_out_frame[17] [5]), 
            .I2(n57604), .I3(\data_out_frame[21] [6]), .O(n57741));
    defparam i1_2_lut_4_lut_adj_1831.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n57301));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_adj_1833 (.I0(n57722), .I1(\data_out_frame[17] [5]), 
            .I2(n57604), .I3(\data_out_frame[19][3] ), .O(n57608));
    defparam i1_2_lut_4_lut_adj_1833.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1834 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[10][1] ), 
            .I2(n58011), .I3(\data_in_frame[12] [5]), .O(n57756));
    defparam i2_3_lut_4_lut_adj_1834.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1835 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[16] [4]), .I3(n59803), .O(n57836));
    defparam i2_3_lut_4_lut_adj_1835.LUT_INIT = 16'h9669;
    SB_LUT4 i12_2_lut_4_lut (.I0(n26279), .I1(n1516), .I2(\data_out_frame[12] [4]), 
            .I3(\data_out_frame[14] [5]), .O(n26931));   // verilog/coms.v(100[12:26])
    defparam i12_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1836 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[7] [7]), 
            .I2(n58108), .I3(n52198), .O(n26899));
    defparam i1_2_lut_4_lut_adj_1836.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1837 (.I0(n57893), .I1(\data_out_frame[16] [0]), 
            .I2(n51946), .I3(GND_net), .O(n53199));
    defparam i1_2_lut_3_lut_adj_1837.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1838 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n57306));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1838.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1839 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n57299));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1839.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n57307));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n57308));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1842 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [6]), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'ha088;
    SB_LUT4 i1_3_lut_4_lut_adj_1843 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[15] [1]), .I3(\data_out_frame[15] [7]), 
            .O(n62292));
    defparam i1_3_lut_4_lut_adj_1843.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1844 (.I0(\data_out_frame[7] [1]), .I1(n26461), 
            .I2(\data_out_frame[9] [2]), .I3(\data_out_frame[6] [6]), .O(n14_adj_5543));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_4_lut_adj_1844.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1845 (.I0(\data_out_frame[4] [1]), .I1(n57577), 
            .I2(n57538), .I3(\data_out_frame[8] [5]), .O(n26461));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1845.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1846 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n60278), .I3(\data_in_frame[7][3] ), .O(n51992));
    defparam i2_3_lut_4_lut_adj_1846.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1847 (.I0(\data_in_frame[13] [0]), .I1(n26069), 
            .I2(n57657), .I3(GND_net), .O(n26517));
    defparam i1_2_lut_3_lut_adj_1847.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n57309));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h5100;
    SB_LUT4 select_777_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1849 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[18] [5]), .I3(n58093), .O(n59475));
    defparam i1_3_lut_4_lut_adj_1849.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1850 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[6] [6]), 
            .I2(n57496), .I3(GND_net), .O(n58105));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1850.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1851 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [5]), .I3(n1168), .O(n57496));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1851.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1852 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n57310));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1852.LUT_INIT = 16'h5100;
    SB_LUT4 select_777_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5457));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1853 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n57962));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_3_lut_adj_1853.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1854 (.I0(\data_out_frame[20]_c [2]), .I1(n52042), 
            .I2(n53027), .I3(\data_out_frame[22][3] ), .O(n52026));
    defparam i2_3_lut_4_lut_adj_1854.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1855 (.I0(n26645), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[11] [4]), .O(n57473));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1855.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[9] [0]), .I3(Kp_23__N_974), .O(n20_adj_5516));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27][2] ), 
            .O(n57311));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h5100;
    SB_LUT4 i20_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_17), .O(n19));
    defparam i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 select_777_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1857 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n57302));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1857.LUT_INIT = 16'h5100;
    SB_LUT4 i23283_3_lut_4_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10]_c [0]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29665));
    defparam i23283_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n57312));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h5100;
    SB_LUT4 i11_3_lut_4_lut (.I0(n52693), .I1(n52308), .I2(n22_adj_5506), 
            .I3(\data_in_frame[6] [0]), .O(n25_adj_5509));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1859 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[7][1] ), .I3(\data_in_frame[4] [7]), .O(n57479));
    defparam i2_3_lut_4_lut_adj_1859.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1860 (.I0(\data_in_frame[9] [7]), .I1(n52693), 
            .I2(n26853), .I3(n25927), .O(n53024));
    defparam i1_2_lut_4_lut_adj_1860.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1861 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n57300));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1861.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_adj_1862 (.I0(n26623), .I1(n57625), .I2(\data_in_frame[16] [3]), 
            .I3(n59679), .O(n26738));
    defparam i1_2_lut_4_lut_adj_1862.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1863 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[16] [0]), .I3(\data_in_frame[13] [1]), .O(n14_adj_5502));
    defparam i5_3_lut_4_lut_adj_1863.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1864 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(n26496), .O(n57975));
    defparam i2_3_lut_4_lut_adj_1864.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1865 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n57298));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1865.LUT_INIT = 16'h5100;
    SB_LUT4 select_777_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1866 (.I0(n26731), .I1(n52024), .I2(\data_out_frame[13] [5]), 
            .I3(n25162), .O(n52173));
    defparam i2_3_lut_4_lut_adj_1866.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1867 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[5] [1]), .O(n8_adj_5498));   // verilog/coms.v(88[17:70])
    defparam i2_2_lut_4_lut_adj_1867.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n57313));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1869 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n6_adj_5496));
    defparam i1_2_lut_3_lut_adj_1869.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1870 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[10] [0]), 
            .I2(n26104), .I3(GND_net), .O(n6_adj_5494));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_3_lut_adj_1870.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1871 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(n58053), .I3(GND_net), .O(n6_adj_5493));
    defparam i1_2_lut_3_lut_adj_1871.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1872 (.I0(n3470), .I1(\FRAME_MATCHER.i [0]), .I2(GND_net), 
            .I3(GND_net), .O(n57399));
    defparam i1_2_lut_adj_1872.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_4_lut_adj_1873 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[13] [6]), .I3(n25266), .O(n57737));
    defparam i1_2_lut_4_lut_adj_1873.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1874 (.I0(n52011), .I1(n58049), .I2(n52390), 
            .I3(n52143), .O(n8_c));
    defparam i3_3_lut_4_lut_adj_1874.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1875 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [2]), .O(n26121));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1875.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_2_lut_4_lut (.I0(n21_c), .I1(n19_c), .I2(n20_adj_5492), 
            .I3(\data_in_frame[21] [7]), .O(n22_adj_5486));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1876 (.I0(\data_in_frame[15] [6]), .I1(n25990), 
            .I2(n26009), .I3(\data_in_frame[13] [5]), .O(n57685));
    defparam i1_2_lut_4_lut_adj_1876.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1877 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(n10_adj_5469), .I3(\data_out_frame[12] [2]), .O(n58108));   // verilog/coms.v(77[16:27])
    defparam i5_3_lut_4_lut_adj_1877.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1878 (.I0(n59287), .I1(n60454), .I2(n53215), 
            .I3(\data_in_frame[17] [5]), .O(Kp_23__N_1551));
    defparam i1_2_lut_4_lut_adj_1878.LUT_INIT = 16'h6996;
    SB_LUT4 i26952_4_lut (.I0(n28413), .I1(n106), .I2(rx_data[2]), .I3(\data_in_frame[20] [2]), 
            .O(n40952));   // verilog/coms.v(94[13:20])
    defparam i26952_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i26953_3_lut (.I0(n40952), .I1(\data_in_frame[20] [2]), .I2(reset), 
            .I3(GND_net), .O(n30222));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1879 (.I0(n10_adj_5304), .I1(n145), .I2(GND_net), 
            .I3(GND_net), .O(n106));
    defparam i1_2_lut_adj_1879.LUT_INIT = 16'h4444;
    SB_LUT4 i26997_4_lut (.I0(n28413), .I1(n106), .I2(rx_data[1]), .I3(\data_in_frame[20] [1]), 
            .O(n40997));   // verilog/coms.v(94[13:20])
    defparam i26997_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i26998_3_lut (.I0(n40997), .I1(\data_in_frame[20] [1]), .I2(reset), 
            .I3(GND_net), .O(n30229));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1880 (.I0(n52338), .I1(n26623), .I2(\data_in_frame[16] [3]), 
            .I3(n58120), .O(n6_adj_5465));
    defparam i1_2_lut_4_lut_adj_1880.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1881 (.I0(n57476), .I1(n57930), .I2(n10_adj_5461), 
            .I3(\data_out_frame[9] [3]), .O(n26432));
    defparam i5_3_lut_4_lut_adj_1881.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1882 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[13] [5]), 
            .I2(n25162), .I3(GND_net), .O(n57891));
    defparam i1_2_lut_3_lut_adj_1882.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1883 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n62300));
    defparam i1_2_lut_3_lut_adj_1883.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1884 (.I0(n26795), .I1(n57574), .I2(n57908), 
            .I3(n57608), .O(n6_adj_5362));
    defparam i1_2_lut_3_lut_4_lut_adj_1884.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1885 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[7] [3]), .O(n62466));
    defparam i1_2_lut_4_lut_adj_1885.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[11] [7]), 
            .O(n10_adj_5379));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1886 (.I0(n57918), .I1(n10_adj_5571), .I2(\data_out_frame[8] [2]), 
            .I3(n26291), .O(n6_adj_5449));
    defparam i1_2_lut_4_lut_adj_1886.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1887 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[4] [3]), .O(n36));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1887.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1888 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n26664));
    defparam i1_2_lut_3_lut_adj_1888.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1889 (.I0(\data_in_frame[19]_c [7]), .I1(n28409), 
            .I2(n28464), .I3(rx_data[7]), .O(n56554));
    defparam i12_4_lut_adj_1889.LUT_INIT = 16'h3a0a;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1890 (.I0(n59684), .I1(\data_in_frame[16] [6]), 
            .I2(n52413), .I3(n57833), .O(n10_adj_5491));
    defparam i2_2_lut_3_lut_4_lut_adj_1890.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1891 (.I0(\data_out_frame[16] [0]), .I1(n51946), 
            .I2(n57893), .I3(n2076), .O(n57747));
    defparam i1_3_lut_4_lut_adj_1891.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1892 (.I0(n23735), .I1(\data_out_frame[20]_c [1]), 
            .I2(\data_out_frame[20][3] ), .I3(n59292), .O(n52991));
    defparam i2_3_lut_4_lut_adj_1892.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1893 (.I0(\data_out_frame[17] [5]), .I1(n57604), 
            .I2(n57848), .I3(GND_net), .O(n6_adj_5409));
    defparam i1_2_lut_3_lut_adj_1893.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1894 (.I0(\data_in_frame[16] [4]), .I1(n26623), 
            .I2(n57996), .I3(n57833), .O(n53052));
    defparam i1_2_lut_3_lut_4_lut_adj_1894.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1895 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[5] [0]), 
            .I2(n10_adj_5463), .I3(\data_out_frame[6] [7]), .O(n6_adj_5407));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1895.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1896 (.I0(n59803), .I1(n51920), .I2(\data_out_frame[18][4] ), 
            .I3(\data_out_frame[18][3] ), .O(n59944));
    defparam i2_3_lut_4_lut_adj_1896.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1897 (.I0(\data_in_frame[10] [6]), .I1(n25976), 
            .I2(n58056), .I3(\data_in_frame[13] [1]), .O(n6_adj_5520));
    defparam i2_2_lut_3_lut_4_lut_adj_1897.LUT_INIT = 16'h6996;
    SB_LUT4 select_779_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5557));
    defparam select_779_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i16308_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30384));   // verilog/coms.v(130[12] 305[6])
    defparam i16308_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15603_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29679));   // verilog/coms.v(130[12] 305[6])
    defparam i15603_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_779_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(byte_transmit_counter[7]), 
            .I3(GND_net), .O(n1_adj_5556));
    defparam select_779_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i16338_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30414));   // verilog/coms.v(130[12] 305[6])
    defparam i16338_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_779_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(byte_transmit_counter[6]), 
            .I3(GND_net), .O(n1_adj_5555));
    defparam select_779_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut_adj_1898 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5262));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1898.LUT_INIT = 16'ha088;
    SB_LUT4 select_779_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(byte_transmit_counter[5]), 
            .I3(GND_net), .O(n1_adj_5554));
    defparam select_779_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i16337_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30413));   // verilog/coms.v(130[12] 305[6])
    defparam i16337_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1899 (.I0(\data_out_frame[16][3] ), .I1(n60167), 
            .I2(n57709), .I3(GND_net), .O(n53178));
    defparam i1_2_lut_3_lut_adj_1899.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1900 (.I0(\FRAME_MATCHER.i[5] ), .I1(n31), .I2(n91), 
            .I3(reset), .O(n28464));
    defparam i3_4_lut_adj_1900.LUT_INIT = 16'h0010;
    SB_LUT4 i16336_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30412));   // verilog/coms.v(130[12] 305[6])
    defparam i16336_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1901 (.I0(\data_out_frame[15] [7]), .I1(n57839), 
            .I2(n57470), .I3(n26138), .O(n51920));
    defparam i2_3_lut_4_lut_adj_1901.LUT_INIT = 16'h6996;
    SB_LUT4 select_779_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n1_adj_5553));
    defparam select_779_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_4_lut_adj_1902 (.I0(\data_out_frame[13] [7]), .I1(n26731), 
            .I2(n52024), .I3(n26818), .O(n57839));
    defparam i1_2_lut_4_lut_adj_1902.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1903 (.I0(\data_out_frame[20]_c [5]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n4_adj_5398));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1903.LUT_INIT = 16'h9696;
    SB_LUT4 select_779_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n1_adj_5552));
    defparam select_779_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_779_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n1_adj_5551));
    defparam select_779_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1904 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n57396));
    defparam i1_2_lut_3_lut_adj_1904.LUT_INIT = 16'hfefe;
    SB_LUT4 select_779_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state [3]), .I2(\byte_transmit_counter[1] ), 
            .I3(GND_net), .O(n1_adj_5550));
    defparam select_779_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1905 (.I0(\data_out_frame[13] [6]), .I1(n26432), 
            .I2(n52024), .I3(GND_net), .O(n57876));
    defparam i1_2_lut_3_lut_adj_1905.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1906 (.I0(\data_out_frame[18][3] ), .I1(n53042), 
            .I2(n57470), .I3(n26138), .O(n51970));
    defparam i1_2_lut_4_lut_adj_1906.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1907 (.I0(reset), .I1(n3470), .I2(rx_data_ready), 
            .I3(\FRAME_MATCHER.rx_data_ready_prev ), .O(n56993));   // verilog/coms.v(94[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_1907.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_1908 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[20]_c [2]), 
            .I2(n52042), .I3(n26539), .O(n57885));
    defparam i1_2_lut_4_lut_adj_1908.LUT_INIT = 16'h6996;
    SB_LUT4 i16335_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30411));   // verilog/coms.v(130[12] 305[6])
    defparam i16335_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16334_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30410));   // verilog/coms.v(130[12] 305[6])
    defparam i16334_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n52026), .I2(\FRAME_MATCHER.state [3]), .I3(n57902), .O(n3_adj_5549));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i1_2_lut_4_lut_adj_1909 (.I0(\data_out_frame[24] [5]), .I1(n23735), 
            .I2(n57571), .I3(n59292), .O(n57902));
    defparam i1_2_lut_4_lut_adj_1909.LUT_INIT = 16'h9669;
    SB_LUT4 i16333_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30409));   // verilog/coms.v(130[12] 305[6])
    defparam i16333_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5261));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16332_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30408));   // verilog/coms.v(130[12] 305[6])
    defparam i16332_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1910 (.I0(n23735), .I1(\data_out_frame[20][3] ), 
            .I2(n57805), .I3(GND_net), .O(n53077));
    defparam i1_2_lut_3_lut_adj_1910.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1911 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5629));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1911.LUT_INIT = 16'heeee;
    SB_LUT4 i16331_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30407));   // verilog/coms.v(130[12] 305[6])
    defparam i16331_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5260));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(byte_transmit_counter[4]), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\byte_transmit_counter[1] ), 
            .O(n4_adj_5630));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'ha8a0;
    SB_LUT4 i29595_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[7]), 
            .I2(n4_adj_5630), .I3(n4_adj_5629), .O(n43569));
    defparam i29595_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i28792_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42760));
    defparam i28792_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16330_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30406));   // verilog/coms.v(130[12] 305[6])
    defparam i16330_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16329_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30405));   // verilog/coms.v(130[12] 305[6])
    defparam i16329_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15818_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29894));
    defparam i15818_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1913 (.I0(n10), .I1(n56993), .I2(GND_net), .I3(GND_net), 
            .O(n57430));
    defparam i1_2_lut_adj_1913.LUT_INIT = 16'heeee;
    SB_LUT4 i16328_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30404));   // verilog/coms.v(130[12] 305[6])
    defparam i16328_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16327_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30403));   // verilog/coms.v(130[12] 305[6])
    defparam i16327_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1914 (.I0(n4_adj_5398), .I1(\data_out_frame[22] [7]), 
            .I2(\data_out_frame[25][2] ), .I3(GND_net), .O(n8_adj_5331));
    defparam i1_2_lut_3_lut_adj_1914.LUT_INIT = 16'h9696;
    SB_LUT4 i14866_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28942));   // verilog/coms.v(130[12] 305[6])
    defparam i14866_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut_adj_1915 (.I0(\FRAME_MATCHER.i [0]), .I1(n58272), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i [1]), .O(n145));
    defparam i3_4_lut_adj_1915.LUT_INIT = 16'h0040;
    SB_LUT4 i2_2_lut_3_lut_adj_1916 (.I0(\data_out_frame[25] [5]), .I1(n26545), 
            .I2(\data_out_frame[23][3] ), .I3(GND_net), .O(n6_adj_5325));
    defparam i2_2_lut_3_lut_adj_1916.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1917 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(n33795), .O(n6_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut_adj_1917.LUT_INIT = 16'hfffe;
    SB_LUT4 i14855_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28931));   // verilog/coms.v(130[12] 305[6])
    defparam i14855_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1918 (.I0(n10_adj_5323), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5631));
    defparam i1_2_lut_adj_1918.LUT_INIT = 16'heeee;
    SB_LUT4 i15821_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29897));
    defparam i15821_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15825_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29901));
    defparam i15825_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14402_4_lut (.I0(n5_adj_5631), .I1(reset), .I2(n57399), .I3(n43390), 
            .O(n58278));
    defparam i14402_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i15829_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29905));
    defparam i15829_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1919 (.I0(n10), .I1(n145), .I2(GND_net), .I3(GND_net), 
            .O(n107));
    defparam i1_2_lut_adj_1919.LUT_INIT = 16'h4444;
    SB_LUT4 i15833_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29909));
    defparam i15833_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14404_3_lut (.I0(n31), .I1(reset), .I2(n57437), .I3(GND_net), 
            .O(n7_adj_18));
    defparam i14404_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1920 (.I0(current_limit[14]), .I1(current_limit[15]), 
            .I2(n26), .I3(current_limit[13]), .O(n21));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i1_4_lut_adj_1920.LUT_INIT = 16'h3332;
    SB_LUT4 n69607_bdd_4_lut (.I0(n69607), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n69610));
    defparam n69607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15837_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29913));
    defparam i15837_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15840_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29916));
    defparam i15840_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16052_3_lut (.I0(\data_in_frame[10]_c [0]), .I1(rx_data[0]), 
            .I2(n57424), .I3(GND_net), .O(n30128));   // verilog/coms.v(130[12] 305[6])
    defparam i16052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16326_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30402));   // verilog/coms.v(130[12] 305[6])
    defparam i16326_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15844_3_lut_4_lut (.I0(n8_adj_12), .I1(n57430), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29920));
    defparam i15844_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16325_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30401));   // verilog/coms.v(130[12] 305[6])
    defparam i16325_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i50405_3_lut (.I0(current_limit[14]), .I1(n26), .I2(current_limit[13]), 
            .I3(GND_net), .O(n65697));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i50405_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21706_4_lut (.I0(n21), .I1(n65697), .I2(\current[15] ), .I3(current_limit[15]), 
            .O(n260));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i21706_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i1_2_lut_3_lut_adj_1921 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[0][1] ), .I3(GND_net), .O(n26401));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1921.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1922 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[4] [6]), .I3(GND_net), .O(n14_adj_5564));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1922.LUT_INIT = 16'h9696;
    SB_LUT4 i16324_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30400));   // verilog/coms.v(130[12] 305[6])
    defparam i16324_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_31_i2_3_lut (.I0(\data_out_frame[3] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1923 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n57959));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_adj_1923.LUT_INIT = 16'h9696;
    SB_LUT4 i47019_3_lut_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[0] [5]), .I3(n26373), .O(n62738));   // verilog/coms.v(80[16:27])
    defparam i47019_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i2_2_lut_3_lut_adj_1924 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0][2] ), 
            .I2(\data_in_frame[5] [0]), .I3(GND_net), .O(n10_adj_5578));   // verilog/coms.v(169[9:87])
    defparam i2_2_lut_3_lut_adj_1924.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1925 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0][2] ), 
            .I2(\data_in_frame[0][3] ), .I3(GND_net), .O(n25842));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1925.LUT_INIT = 16'h9696;
    SB_LUT4 i16323_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30399));   // verilog/coms.v(130[12] 305[6])
    defparam i16323_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16322_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30398));   // verilog/coms.v(130[12] 305[6])
    defparam i16322_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i26982_4_lut (.I0(n172), .I1(n107), .I2(rx_data[6]), .I3(\data_in_frame[4] [6]), 
            .O(n40982));   // verilog/coms.v(94[13:20])
    defparam i26982_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i26983_3_lut (.I0(n40982), .I1(\data_in_frame[4] [6]), .I2(reset), 
            .I3(GND_net), .O(n29997));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16321_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30397));   // verilog/coms.v(130[12] 305[6])
    defparam i16321_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i52882_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[7] [7]), .I2(n7_adj_10), 
            .I3(GND_net), .O(n56518));   // verilog/coms.v(94[13:20])
    defparam i52882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15428_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29504));
    defparam i15428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i52883_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[7] [6]), .I2(n7_adj_10), 
            .I3(GND_net), .O(n56520));   // verilog/coms.v(94[13:20])
    defparam i52883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n56504));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15874_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[3][0] ), .O(n29950));
    defparam i15874_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15877_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[3][1] ), .O(n29953));
    defparam i15877_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15881_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[3][2] ), .O(n29957));
    defparam i15881_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15884_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[3][3] ), .O(n29960));
    defparam i15884_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15887_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[3][4] ), .O(n29963));
    defparam i15887_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15890_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29966));
    defparam i15890_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15893_3_lut_4_lut (.I0(n28439), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[3][6] ), .O(n29969));
    defparam i15893_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15422_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29498));
    defparam i15422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut_adj_1926 (.I0(n28439), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[3]_c [7]), .O(n56700));
    defparam i11_4_lut_4_lut_adj_1926.LUT_INIT = 16'hfe10;
    SB_LUT4 i52881_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[7] [0]), .I2(n7_adj_10), 
            .I3(GND_net), .O(n56514));   // verilog/coms.v(94[13:20])
    defparam i52881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14378_3_lut_4_lut (.I0(n10), .I1(n58272), .I2(reset), .I3(n8_adj_15), 
            .O(n7));
    defparam i14378_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i16320_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30396));   // verilog/coms.v(130[12] 305[6])
    defparam i16320_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16318_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30394));   // verilog/coms.v(130[12] 305[6])
    defparam i16318_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 equal_307_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_13));   // verilog/coms.v(158[12:15])
    defparam equal_307_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1927 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n31));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1927.LUT_INIT = 16'hbfbf;
    SB_LUT4 i15419_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29495));
    defparam i15419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16317_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30393));   // verilog/coms.v(130[12] 305[6])
    defparam i16317_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16316_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30392));   // verilog/coms.v(130[12] 305[6])
    defparam i16316_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i29420_2_lut_3_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n43390));
    defparam i29420_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i16315_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30391));   // verilog/coms.v(130[12] 305[6])
    defparam i16315_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16314_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30390));   // verilog/coms.v(130[12] 305[6])
    defparam i16314_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n69841));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69841_bdd_4_lut (.I0(n69841), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n63105));
    defparam n69841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54044 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n69835));
    defparam byte_transmit_counter_0__bdd_4_lut_54044.LUT_INIT = 16'he4aa;
    SB_LUT4 n69835_bdd_4_lut (.I0(n69835), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n63111));
    defparam n69835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50512_2_lut_3_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(n8_adj_15), 
            .I2(n91), .I3(GND_net), .O(n65728));   // verilog/coms.v(158[12:15])
    defparam i50512_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1928 (.I0(\FRAME_MATCHER.i[5] ), .I1(n8_adj_15), 
            .I2(n57410), .I3(GND_net), .O(n105));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1928.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n63172), .I2(n63173), .I3(\byte_transmit_counter[2] ), 
            .O(n69595));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i15973_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[7]), 
            .I3(\data_in_frame[6]_c [7]), .O(n30049));
    defparam i15973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15970_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[6]), 
            .I3(\data_in_frame[6]_c [6]), .O(n30046));
    defparam i15970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_30_i2_3_lut (.I0(\data_out_frame[3] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5452));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15967_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n30043));
    defparam i15967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15964_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n30040));
    defparam i15964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15961_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n30037));
    defparam i15961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15958_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n30034));
    defparam i15958_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15955_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n30031));
    defparam i15955_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69595_bdd_4_lut (.I0(n69595), .I1(n62918), .I2(n62917), .I3(\byte_transmit_counter[2] ), 
            .O(n69598));
    defparam n69595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15952_3_lut_4_lut (.I0(n8), .I1(n57430), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n30028));
    defparam i15952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16313_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30389));   // verilog/coms.v(130[12] 305[6])
    defparam i16313_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15416_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29492));
    defparam i15416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_293_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_15));   // verilog/coms.v(158[12:15])
    defparam equal_293_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n41114), .I3(\FRAME_MATCHER.i [0]), .O(n59370));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut_adj_1929.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_300_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_12));   // verilog/coms.v(158[12:15])
    defparam equal_300_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i15847_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29923));
    defparam i15847_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15850_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29926));
    defparam i15850_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15854_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29930));
    defparam i15854_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53843 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63025), .I2(n63026), .I3(\byte_transmit_counter[2] ), 
            .O(n69589));
    defparam byte_transmit_counter_1__bdd_4_lut_53843.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54039 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n69829));
    defparam byte_transmit_counter_0__bdd_4_lut_54039.LUT_INIT = 16'he4aa;
    SB_LUT4 n69829_bdd_4_lut (.I0(n69829), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n63114));
    defparam n69829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15857_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29933));
    defparam i15857_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15861_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29937));
    defparam i15861_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15864_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29940));
    defparam i15864_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15867_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29943));
    defparam i15867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15871_3_lut_4_lut (.I0(n8_adj_13), .I1(n57430), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29947));
    defparam i15871_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i27132_4_lut (.I0(n105), .I1(n65728), .I2(rx_data[1]), .I3(\data_in_frame[16] [1]), 
            .O(n41131));   // verilog/coms.v(94[13:20])
    defparam i27132_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i27133_3_lut (.I0(n41131), .I1(\data_in_frame[16] [1]), .I2(reset), 
            .I3(GND_net), .O(n30370));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16184_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n30260));
    defparam i16184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16312_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30388));   // verilog/coms.v(130[12] 305[6])
    defparam i16312_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16150_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n30226));
    defparam i16150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16147_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n30223));
    defparam i16147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69589_bdd_4_lut (.I0(n69589), .I1(n63122), .I2(n63121), .I3(\byte_transmit_counter[2] ), 
            .O(n69592));
    defparam n69589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16311_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30387));   // verilog/coms.v(130[12] 305[6])
    defparam i16311_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16310_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30386));   // verilog/coms.v(130[12] 305[6])
    defparam i16310_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16143_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n30219));
    defparam i16143_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16140_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n30216));
    defparam i16140_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16309_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30385));   // verilog/coms.v(130[12] 305[6])
    defparam i16309_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16137_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n30213));
    defparam i16137_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15413_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29489));
    defparam i15413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16133_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n30209));
    defparam i16133_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20980_3_lut_4_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n30466));
    defparam i20980_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16130_3_lut_4_lut (.I0(n10_adj_5323), .I1(n57434), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n30206));
    defparam i16130_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15410_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29486));
    defparam i15410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16319_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30395));   // verilog/coms.v(130[12] 305[6])
    defparam i16319_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1930 (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(GND_net), .O(n10_adj_5304));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1930.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1931 (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(GND_net), .O(n10));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1931.LUT_INIT = 16'hfefe;
    SB_LUT4 select_777_Select_28_i2_3_lut (.I0(\data_out_frame[3] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15407_3_lut_4_lut (.I0(n28421), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29483));
    defparam i15407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53838 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63037), .I2(n63038), .I3(\byte_transmit_counter[2] ), 
            .O(n69583));
    defparam byte_transmit_counter_1__bdd_4_lut_53838.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_4_lut (.I0(n40928), .I1(reset), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n3470), .O(n57434));   // verilog/coms.v(158[12:15])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 n69583_bdd_4_lut (.I0(n69583), .I1(n63119), .I2(n63118), .I3(\byte_transmit_counter[2] ), 
            .O(n69586));
    defparam n69583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54034 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n69823));
    defparam byte_transmit_counter_0__bdd_4_lut_54034.LUT_INIT = 16'he4aa;
    SB_LUT4 n69823_bdd_4_lut (.I0(n69823), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n63126));
    defparam n69823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1932 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3][4] ), .I3(\data_in_frame[3][3] ), .O(n6_adj_5560));   // verilog/coms.v(79[16:43])
    defparam i2_2_lut_3_lut_4_lut_adj_1932.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1933 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3][4] ), .I3(n25784), .O(n57669));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1933.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n69466), .I2(n65787), .I3(byte_transmit_counter[4]), .O(n69817));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1934 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3][4] ), .I3(\data_in_frame[5] [6]), .O(n57694));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1934.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_27_i2_3_lut (.I0(\data_out_frame[3] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 n69817_bdd_4_lut (.I0(n69817), .I1(n69580), .I2(n7_adj_5635), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n69817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53833 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63019), .I2(n63020), .I3(\byte_transmit_counter[2] ), 
            .O(n69577));
    defparam byte_transmit_counter_1__bdd_4_lut_53833.LUT_INIT = 16'he4aa;
    SB_LUT4 i15716_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[7]), .I3(\data_in_frame[23] [7]), .O(n29792));
    defparam i15716_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15713_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[6]), .I3(\data_in_frame[23] [6]), .O(n29789));
    defparam i15713_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15710_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[5]), .I3(\data_in_frame[23] [5]), .O(n29786));
    defparam i15710_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15707_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[4]), .I3(\data_in_frame[23] [4]), .O(n29783));
    defparam i15707_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1935 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(n57446), .O(n57914));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1935.LUT_INIT = 16'h6996;
    SB_LUT4 i15695_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[3]), .I3(\data_in_frame[23] [3]), .O(n29771));
    defparam i15695_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n69577_bdd_4_lut (.I0(n69577), .I1(n63011), .I2(n63010), .I3(\byte_transmit_counter[2] ), 
            .O(n69580));
    defparam n69577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1936 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(n57519), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1936.LUT_INIT = 16'h6996;
    SB_LUT4 i15692_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[2]), .I3(\data_in_frame[23] [2]), .O(n29768));
    defparam i15692_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15685_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[1]), .I3(\data_in_frame[23] [1]), .O(n29761));
    defparam i15685_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53828 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63004), .I2(n63005), .I3(\byte_transmit_counter[2] ), 
            .O(n69571));
    defparam byte_transmit_counter_1__bdd_4_lut_53828.LUT_INIT = 16'he4aa;
    SB_LUT4 n69571_bdd_4_lut (.I0(n69571), .I1(n63164), .I2(n63163), .I3(\byte_transmit_counter[2] ), 
            .O(n69574));
    defparam n69571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15650_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[0]), .I3(\data_in_frame[23] [0]), .O(n29726));
    defparam i15650_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1937 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(n58024), .I3(n53095), .O(n62546));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1937.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53823 (.I0(\byte_transmit_counter[1] ), 
            .I1(\data_out_frame[21] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(\byte_transmit_counter[0] ), .O(n69565));
    defparam byte_transmit_counter_1__bdd_4_lut_53823.LUT_INIT = 16'he4aa;
    SB_LUT4 i26967_4_lut (.I0(n172), .I1(n107), .I2(rx_data[5]), .I3(\data_in_frame[4] [5]), 
            .O(n40967));   // verilog/coms.v(94[13:20])
    defparam i26967_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i26968_3_lut (.I0(n40967), .I1(\data_in_frame[4] [5]), .I2(reset), 
            .I3(GND_net), .O(n29994));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5259));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1938 (.I0(ID[6]), .I1(\data_in_frame[0][7] ), .I2(\data_in_frame[0] [6]), 
            .I3(ID[7]), .O(n12_adj_5636));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1938.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1939 (.I0(\data_in_frame[0][1] ), .I1(\data_in_frame[0][2] ), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_5637));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1939.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1940 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0][3] ), 
            .I2(ID[4]), .I3(ID[3]), .O(n11_adj_5638));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1940.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1941 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[0] [5]), 
            .I2(ID[0]), .I3(ID[5]), .O(n9_adj_5639));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1941.LUT_INIT = 16'h7bde;
    SB_LUT4 n69565_bdd_4_lut (.I0(n69565), .I1(\data_out_frame[22] [5]), 
            .I2(\data_out_frame[20]_c [5]), .I3(\byte_transmit_counter[0] ), 
            .O(n69568));
    defparam n69565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1942 (.I0(n9_adj_5639), .I1(n11_adj_5638), .I2(n10_adj_5637), 
            .I3(n12_adj_5636), .O(n22911));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1942.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1943 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n57506));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1943.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1944 (.I0(\data_in_frame[0][0] ), .I1(Kp_23__N_748), 
            .I2(GND_net), .I3(GND_net), .O(n57651));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1944.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53852 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n69559));
    defparam byte_transmit_counter_0__bdd_4_lut_53852.LUT_INIT = 16'he4aa;
    SB_LUT4 i15608_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[7]), .I3(\data_in_frame[21] [7]), .O(n29684));
    defparam i15608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1945 (.I0(\data_in_frame[0][7] ), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57638));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1945.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1946 (.I0(\data_in_frame[0][2] ), .I1(\data_in_frame[0][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n57728));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1946.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_760));   // verilog/coms.v(99[12:25])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1947 (.I0(Kp_23__N_760), .I1(n57728), .I2(n57638), 
            .I3(\data_in_frame[0][3] ), .O(Kp_23__N_748));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1947.LUT_INIT = 16'h6996;
    SB_LUT4 i46956_3_lut (.I0(\data_in_frame[0][7] ), .I1(n26401), .I2(\data_in_frame[1] [1]), 
            .I3(GND_net), .O(n62674));
    defparam i46956_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i15604_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[6]), .I3(\data_in_frame[21] [6]), .O(n29680));
    defparam i15604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1948 (.I0(n25842), .I1(n14_adj_5342), .I2(Kp_23__N_748), 
            .I3(\data_in_frame[2] [1]), .O(n18_adj_5640));
    defparam i7_4_lut_adj_1948.LUT_INIT = 16'h0440;
    SB_LUT4 n69559_bdd_4_lut (.I0(n69559), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20]_c [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n69562));
    defparam n69559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15590_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[5]), .I3(\data_in_frame[21] [5]), .O(n29666));
    defparam i15590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15581_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[4]), .I3(\data_in_frame[21] [4]), .O(n29657));
    defparam i15581_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1949 (.I0(\data_in_frame[2] [0]), .I1(n18_adj_5640), 
            .I2(n62674), .I3(n57651), .O(n20_adj_5641));
    defparam i9_4_lut_adj_1949.LUT_INIT = 16'h0804;
    SB_LUT4 i15573_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[3]), .I3(\data_in_frame[21] [3]), .O(n29649));
    defparam i15573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1950 (.I0(n52588), .I1(n20_adj_5641), .I2(n62738), 
            .I3(n25835), .O(n60517));
    defparam i10_4_lut_adj_1950.LUT_INIT = 16'h0008;
    SB_LUT4 i5_4_lut_adj_1951 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [6]), .O(n12_adj_5642));
    defparam i5_4_lut_adj_1951.LUT_INIT = 16'h8000;
    SB_LUT4 i15570_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[2]), .I3(\data_in_frame[21] [2]), .O(n29646));
    defparam i15570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1952 (.I0(n22911), .I1(n12_adj_5642), .I2(n60517), 
            .I3(\data_in_frame[1] [5]), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i6_4_lut_adj_1952.LUT_INIT = 16'h4000;
    SB_LUT4 i15565_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[1]), .I3(\data_in_frame[21] [1]), .O(n29641));
    defparam i15565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15562_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57427), 
            .I2(rx_data[0]), .I3(\data_in_frame[21] [0]), .O(n29638));
    defparam i15562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_1_lut (.I0(reset), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2873));   // verilog/coms.v(94[13:20])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 select_777_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(n63105), .I2(n63126), .I3(byte_transmit_counter[3]), .O(n69553));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69553_bdd_4_lut (.I0(n69553), .I1(n63029), .I2(n63028), .I3(byte_transmit_counter[3]), 
            .O(n69556));
    defparam n69553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53813 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n69547));
    defparam byte_transmit_counter_0__bdd_4_lut_53813.LUT_INIT = 16'he4aa;
    SB_LUT4 n69547_bdd_4_lut (.I0(n69547), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n69550));
    defparam n69547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54029 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n69805));
    defparam byte_transmit_counter_0__bdd_4_lut_54029.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_53808 (.I0(\byte_transmit_counter[2] ), 
            .I1(n63114), .I2(n63111), .I3(byte_transmit_counter[3]), .O(n69541));
    defparam byte_transmit_counter_2__bdd_4_lut_53808.LUT_INIT = 16'he4aa;
    SB_LUT4 n69805_bdd_4_lut (.I0(n69805), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n69808));
    defparam n69805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69541_bdd_4_lut (.I0(n69541), .I1(n63023), .I2(n63022), .I3(byte_transmit_counter[3]), 
            .O(n69544));
    defparam n69541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53818 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63007), .I2(n63008), .I3(\byte_transmit_counter[2] ), 
            .O(n69535));
    defparam byte_transmit_counter_1__bdd_4_lut_53818.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54024 (.I0(byte_transmit_counter[3]), 
            .I1(n69472), .I2(n65732), .I3(byte_transmit_counter[4]), .O(n69799));
    defparam byte_transmit_counter_3__bdd_4_lut_54024.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_4_lut_adj_1953 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1951), .I3(n1954), .O(n25550));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1953.LUT_INIT = 16'h4000;
    SB_LUT4 i2_3_lut_4_lut_adj_1954 (.I0(n1951), .I1(n4452), .I2(n1954), 
            .I3(n1957), .O(n59374));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1954.LUT_INIT = 16'h2000;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1951), .I1(n4452), .I2(n4_adj_5338), 
            .I3(\FRAME_MATCHER.i_31__N_2514 ), .O(n60102));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 n69535_bdd_4_lut (.I0(n69535), .I1(n63155), .I2(n63154), .I3(\byte_transmit_counter[2] ), 
            .O(n69538));
    defparam n69535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69799_bdd_4_lut (.I0(n69799), .I1(n69574), .I2(n7_adj_5643), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n69799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1955 (.I0(n58272), .I1(\FRAME_MATCHER.i[4] ), .I2(\FRAME_MATCHER.i[3] ), 
            .I3(GND_net), .O(n57410));
    defparam i2_3_lut_adj_1955.LUT_INIT = 16'hf7f7;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53803 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n69529));
    defparam byte_transmit_counter_0__bdd_4_lut_53803.LUT_INIT = 16'he4aa;
    SB_LUT4 n69529_bdd_4_lut (.I0(n69529), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n69532));
    defparam n69529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53789 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n69523));
    defparam byte_transmit_counter_0__bdd_4_lut_53789.LUT_INIT = 16'he4aa;
    SB_LUT4 n69523_bdd_4_lut (.I0(n69523), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n69526));
    defparam n69523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53784 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n69517));
    defparam byte_transmit_counter_0__bdd_4_lut_53784.LUT_INIT = 16'he4aa;
    SB_LUT4 n69517_bdd_4_lut (.I0(n69517), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n69520));
    defparam n69517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53779 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n69511));
    defparam byte_transmit_counter_0__bdd_4_lut_53779.LUT_INIT = 16'he4aa;
    SB_LUT4 n69511_bdd_4_lut (.I0(n69511), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n69514));
    defparam n69511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53794 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63064), .I2(n63065), .I3(\byte_transmit_counter[2] ), 
            .O(n69499));
    defparam byte_transmit_counter_1__bdd_4_lut_53794.LUT_INIT = 16'he4aa;
    SB_LUT4 n69499_bdd_4_lut (.I0(n69499), .I1(n63116), .I2(n63115), .I3(\byte_transmit_counter[2] ), 
            .O(n69502));
    defparam n69499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54009 (.I0(byte_transmit_counter[3]), 
            .I1(n69478), .I2(n65735), .I3(byte_transmit_counter[4]), .O(n69793));
    defparam byte_transmit_counter_3__bdd_4_lut_54009.LUT_INIT = 16'he4aa;
    SB_LUT4 n69793_bdd_4_lut (.I0(n69793), .I1(n69598), .I2(n7_adj_5644), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n69793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1956 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [4]), .I3(n58072), .O(n58027));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1956.LUT_INIT = 16'h9669;
    SB_LUT4 i23282_3_lut_4_lut (.I0(deadband[1]), .I1(\data_in_frame[16] [1]), 
            .I2(Kp_23__N_1748), .I3(n33793), .O(n29880));
    defparam i23282_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i20985_3_lut (.I0(n30), .I1(PWMLimit[15]), .I2(n365), .I3(GND_net), 
            .O(n32));
    defparam i20985_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n63060), .I3(n63058), 
            .O(n7_adj_5647));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1957 (.I0(\FRAME_MATCHER.i[5] ), .I1(n57410), .I2(GND_net), 
            .I3(GND_net), .O(n41114));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_adj_1957.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53774 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n69487));
    defparam byte_transmit_counter_0__bdd_4_lut_53774.LUT_INIT = 16'he4aa;
    SB_LUT4 n69487_bdd_4_lut (.I0(n69487), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n69490));
    defparam n69487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1958 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));
    defparam i2_3_lut_adj_1958.LUT_INIT = 16'hf7f7;
    SB_LUT4 i4_3_lut_4_lut_adj_1959 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[20] [1]), .O(n23_adj_5489));
    defparam i4_3_lut_4_lut_adj_1959.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54004 (.I0(byte_transmit_counter[3]), 
            .I1(n69484), .I2(n65734), .I3(byte_transmit_counter[4]), .O(n69787));
    defparam byte_transmit_counter_3__bdd_4_lut_54004.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53764 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63001), .I2(n63002), .I3(\byte_transmit_counter[2] ), 
            .O(n69481));
    defparam byte_transmit_counter_1__bdd_4_lut_53764.LUT_INIT = 16'he4aa;
    SB_LUT4 n69481_bdd_4_lut (.I0(n69481), .I1(n63128), .I2(n63127), .I3(\byte_transmit_counter[2] ), 
            .O(n69484));
    defparam n69481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n63051), .I3(n63049), 
            .O(n7_adj_5648));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1960 (.I0(\data_in_frame[6]_c [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n58144), .I3(GND_net), .O(n57648));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_3_lut_adj_1960.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53750 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62995), .I2(n62996), .I3(\byte_transmit_counter[2] ), 
            .O(n69475));
    defparam byte_transmit_counter_1__bdd_4_lut_53750.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1961 (.I0(\data_in_frame[6]_c [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n26370), .I3(Kp_23__N_878), .O(n57663));   // verilog/coms.v(80[16:43])
    defparam i2_3_lut_4_lut_adj_1961.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n63045), .I3(n63043), 
            .O(n7_adj_5644));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 n69475_bdd_4_lut (.I0(n69475), .I1(n63152), .I2(n63151), .I3(\byte_transmit_counter[2] ), 
            .O(n69478));
    defparam n69475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1962 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n58114), .I3(GND_net), .O(n57587));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1962.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53745 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63016), .I2(n63017), .I3(\byte_transmit_counter[2] ), 
            .O(n69469));
    defparam byte_transmit_counter_1__bdd_4_lut_53745.LUT_INIT = 16'he4aa;
    SB_LUT4 n69469_bdd_4_lut (.I0(n69469), .I1(n63014), .I2(n63013), .I3(\byte_transmit_counter[2] ), 
            .O(n69472));
    defparam n69469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n63075), .I3(n63073), 
            .O(n7_adj_5643));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53740 (.I0(\byte_transmit_counter[1] ), 
            .I1(n63139), .I2(n63140), .I3(\byte_transmit_counter[2] ), 
            .O(n69463));
    defparam byte_transmit_counter_1__bdd_4_lut_53740.LUT_INIT = 16'he4aa;
    SB_LUT4 n69463_bdd_4_lut (.I0(n69463), .I1(n63143), .I2(n63142), .I3(\byte_transmit_counter[2] ), 
            .O(n69466));
    defparam n69463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69787_bdd_4_lut (.I0(n69787), .I1(n69592), .I2(n7_adj_5648), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n69787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n63069), .I3(n63067), 
            .O(n7_adj_5330));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1963 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n25266), .I3(GND_net), .O(n52001));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1963.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53999 (.I0(byte_transmit_counter[3]), 
            .I1(n67824), .I2(n65564), .I3(byte_transmit_counter[4]), .O(n69781));
    defparam byte_transmit_counter_3__bdd_4_lut_53999.LUT_INIT = 16'he4aa;
    SB_LUT4 n69781_bdd_4_lut (.I0(n69781), .I1(n69586), .I2(n7_adj_5647), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n69781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n63054), .I3(n63052), 
            .O(n7_adj_5635));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i15949_3_lut_4_lut (.I0(n10), .I1(n57434), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n30025));
    defparam i15949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.tx_o(tx_o), .clk16MHz(clk16MHz), .tx_data({tx_data}), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
            .n29690(n29690), .tx_active(tx_active), .GND_net(GND_net), 
            .n58304(n58304), .r_Clock_Count({r_Clock_Count}), .VCC_net(VCC_net), 
            .n58925(n58925), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n6(n6_adj_19), .n4940(n4940), .n29(n29), .n23(n23_adj_5650), 
            .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
            .n27(n27), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .baudrate({baudrate}), .clk16MHz(clk16MHz), 
            .\r_SM_Main[2] (\r_SM_Main[2]_adj_20 ), .r_Rx_Data(r_Rx_Data), 
            .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
            .n4937(n4937), .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
            .n29(n29), .n23(n23_adj_5650), .n61106(n61106), .n29912(n29912), 
            .rx_data({rx_data}), .n61058(n61058), .n57317(n57317), .\r_SM_Main[1] (\r_SM_Main[1]_adj_21 ), 
            .n27(n27), .n27754(n27754), .n61138(n61138), .n29900(n29900), 
            .VCC_net(VCC_net), .n25593(n25593), .n29798(n29798), .n29797(n29797), 
            .n29796(n29796), .\r_Bit_Index[0] (\r_Bit_Index[0] ), .r_Clock_Count({r_Clock_Count_adj_30}), 
            .n27996(n27996), .n58373(n58373), .n30533(n30533), .n53222(n53222), 
            .rx_data_ready(rx_data_ready), .n30529(n30529), .n30231(n30231), 
            .n30230(n30230), .n4940(n4940), .\r_SM_Main[0] (r_SM_Main[0]), 
            .n58925(n58925), .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), 
            .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), 
            .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), 
            .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), 
            .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), .n61170(n61170), 
            .n61154(n61154), .n61090(n61090), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
            .n61074(n61074), .n61122(n61122)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (tx_o, clk16MHz, tx_data, r_SM_Main, \r_SM_Main_2__N_3536[1] , 
            n29690, tx_active, GND_net, n58304, r_Clock_Count, VCC_net, 
            n58925, \r_SM_Main_2__N_3545[0] , n6, n4940, n29, n23, 
            \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , n27, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    input n29690;
    output tx_active;
    input GND_net;
    input n58304;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input n58925;
    input \r_SM_Main_2__N_3545[0] ;
    output n6;
    input n4940;
    input n29;
    input n23;
    input \o_Rx_DV_N_3488[12] ;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n3, n40736, n25100;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n53254, n65613, n58401;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n58896, n53252, n40708;
    wire [2:0]n460;
    
    wire n57295, n29222;
    wire [8:0]n41;
    
    wire n50928, n50927, n50926, n50925, n50924, n50923, n50922, 
        n50921, n69865, n3_adj_5258, n60888, n60894, n63133, n63134, 
        n63167, n63166, n65598, n65595, n9, n69604, n14, n15, 
        n69601;
    
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n40736), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n53254), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i12_4_lut (.I0(n65613), .I1(n58401), .I2(r_Bit_Index[0]), 
            .I3(n58896), .O(n53252));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i53656_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n40708));
    defparam i53656_4_lut.LUT_INIT = 16'h1113;
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29690));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i26725_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i26725_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i42480_rep_29_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n58896));
    defparam i42480_rep_29_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n58304), .I1(n58896), .I2(r_SM_Main[1]), .I3(n57295), 
            .O(n29222));
    defparam i1_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i16_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Clock_Count_1953_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n50928), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1953_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n50927), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_9 (.CI(n50927), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n50928));
    SB_LUT4 r_Clock_Count_1953_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n50926), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_8 (.CI(n50926), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n50927));
    SB_LUT4 r_Clock_Count_1953_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n50925), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_7 (.CI(n50925), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n50926));
    SB_LUT4 r_Clock_Count_1953_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n50924), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_6 (.CI(n50924), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n50925));
    SB_LUT4 r_Clock_Count_1953_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n50923), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_5 (.CI(n50923), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n50924));
    SB_LUT4 r_Clock_Count_1953_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n50922), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_4 (.CI(n50922), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n50923));
    SB_LUT4 r_Clock_Count_1953_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n50921), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_3 (.CI(n50921), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n50922));
    SB_LUT4 r_Clock_Count_1953_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n50921));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n58401), 
            .D(n460[1]), .R(n29222));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n58401), 
            .D(n460[2]), .R(n29222));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Clock_Count_1953__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n40736), .D(n41[1]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n40736), .D(n41[2]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n40736), .D(n41[3]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n40736), .D(n41[4]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n40736), .D(n41[5]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n40736), .D(n41[6]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n40736), .D(n41[7]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n40736), .D(n41[8]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n40736), .D(n41[0]), .R(n40708));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n53252));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n69865));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5258), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25100), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n58925), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n25100));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut (.I0(n4940), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n60888));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1102 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n60888), .O(n60894));
    defparam i1_4_lut_adj_1102.LUT_INIT = 16'h0100;
    SB_LUT4 i10_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n60894), .O(n3_adj_5258));   // verilog/uart_tx.v(32[16:25])
    defparam i10_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i47405_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63133));
    defparam i47405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47406_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63134));
    defparam i47406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47439_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63167));
    defparam i47439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47438_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n63166));
    defparam i47438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n57295));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i50914_3_lut (.I0(n57295), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4940), 
            .I3(GND_net), .O(n65598));   // verilog/uart_tx.v(32[16:25])
    defparam i50914_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i50911_4_lut (.I0(n65598), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65595));   // verilog/uart_tx.v(32[16:25])
    defparam i50911_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i23_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n65595), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n9));   // verilog/uart_tx.v(32[16:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut (.I0(n9), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n53254));   // verilog/uart_tx.v(32[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40736));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(n69604), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i53704_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n58401));
    defparam i53704_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4940), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n40736), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n69865));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i50949_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n65613));   // verilog/uart_tx.v(32[16:25])
    defparam i50949_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(n63166), 
            .I2(n63167), .I3(r_Bit_Index[1]), .O(n69601));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69601_bdd_4_lut (.I0(n69601), .I1(n63134), .I2(n63133), .I3(r_Bit_Index[1]), 
            .O(n69604));
    defparam n69601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, baudrate, clk16MHz, \r_SM_Main[2] , r_Rx_Data, 
            RX_N_2, \o_Rx_DV_N_3488[12] , n4937, \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[24] , n29, n23, n61106, n29912, rx_data, 
            n61058, n57317, \r_SM_Main[1] , n27, n27754, n61138, 
            n29900, VCC_net, n25593, n29798, n29797, n29796, \r_Bit_Index[0] , 
            r_Clock_Count, n27996, n58373, n30533, n53222, rx_data_ready, 
            n30529, n30231, n30230, n4940, \r_SM_Main[0] , n58925, 
            \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , n61170, n61154, 
            n61090, \r_SM_Main_2__N_3536[1] , n61074, n61122) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [31:0]baudrate;
    input clk16MHz;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[12] ;
    input n4937;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    output n61106;
    input n29912;
    output [7:0]rx_data;
    output n61058;
    input n57317;
    output \r_SM_Main[1] ;
    output n27;
    output n27754;
    output n61138;
    input n29900;
    input VCC_net;
    output n25593;
    input n29798;
    input n29797;
    input n29796;
    output \r_Bit_Index[0] ;
    output [7:0]r_Clock_Count;
    output n27996;
    output n58373;
    input n30533;
    input n53222;
    output rx_data_ready;
    input n30529;
    input n30231;
    input n30230;
    input n4940;
    input \r_SM_Main[0] ;
    output n58925;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n61170;
    output n61154;
    output n61090;
    output \r_SM_Main_2__N_3536[1] ;
    output n61074;
    output n61122;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n2239;
    wire [23:0]n8217;
    wire [23:0]n294;
    
    wire n2365, n2099;
    wire [23:0]n8191;
    
    wire n2228, n2236, n2362, n29_c, n2098, n2227, n2100, n2229, 
        n14, n37, n32, n43, n68123, n31, n68124, n35, n33, 
        n65973, n65967, n12, n65958, n68462, n68034, n2101, n2230, 
        n41, n2102, n2231, n39, n2103, n2232, n37_adj_4987, n25645, 
        n48, n2240, n2105, n2234, n8, n23_c, n68125, n25, n68126, 
        n21, n65993, n66898, n10, n67678, n2106, n2235, n2104, 
        n2233, n31_adj_4988, n33_adj_4989, n35_adj_4990, n27_c, n68032, 
        n1966;
    wire [23:0]n8165;
    
    wire n65980, n67892, n1968, n68580, n68119, n68602, n3155, 
        n68603, n1967, n1971, n3154, n68599, n37_adj_4991, n1972, 
        n3153, n68394, n3152, n68395, n35_adj_4992, n1977, n2109, 
        n1969, n3151, n48_adj_4993, n41_adj_4994, n1970, n39_adj_4995, 
        n1973, n1974, n2107, n29_adj_4996, n31_adj_4997, n33_adj_4998, 
        n62168, n62116, n62166, n61214, n62176, n62172, n62174, 
        n2108, n27_adj_4999, n66371, n30, n38, n58472, n26, n67894, 
        n67895, n66365, n28, n66363, n68371, n67083, n68545, n68546, 
        n68483, n1975, n1831;
    wire [23:0]n8139;
    
    wire n1839, n1832, n1833, n1836, n1837, n35_adj_5000, n37_adj_5001, 
        n1834, n41_adj_5002, n1835, n39_adj_5003, n1693;
    wire [23:0]n8113;
    
    wire n1694, n1697, n39_adj_5004, n1698, n37_adj_5005, n25636, 
        n48_adj_5006, n1841, n1695, n43_adj_5007, n1696, n41_adj_5008, 
        n1699, n1701, n31_adj_5009, n1838, n33_adj_5010, n35_adj_5011, 
        n1702, n1840, n29_adj_5012, n66408, n32_adj_5013, n40, n28_adj_5014, 
        n67916, n67917, n66400, n30_adj_5015, n66398, n68347, n67071, 
        n68533, n68534, n1700, n29_adj_5016, n31_adj_5017, n33_adj_5018, 
        n1976, n27_adj_5019, n66390, n30_adj_5020, n38_adj_5021, n26_adj_5022, 
        n67912, n67913, n66383, n28_adj_5023, n66381, n68369, n67075, 
        n68543, n68544, n68485, n48_adj_5024, n2237, n2238, n25_adj_5025, 
        n27_adj_5026, n29_adj_5027, n2110, n23_adj_5028, n66353, n66348, 
        n22, n28_adj_5029, n30_adj_5030, n26_adj_5031, n34, n24, 
        n66346, n68373, n68374, n68190, n68079, n66350, n68147, 
        n67093, n68345, n68346, n2364, n23_adj_5032, n25_adj_5033, 
        n2363, n27_adj_5034, n2366, n21_adj_5035, n66332, n33_adj_5036, 
        n31_adj_5037, n66325, n2367, n20, n26_adj_5038, n28_adj_5039, 
        n24_adj_5040, n35_adj_5041, n32_adj_5042, n22_adj_5043, n66323, 
        n68375, n37_adj_5044, n68376, n39_adj_5045, n68186, n68077, 
        n66329, n68452, n41_adj_5046, n67099, n68519, n2355, n68520, 
        n2354, n68447;
    wire [23:0]n8243;
    
    wire n2486, n2487, n25_adj_5047, n27_adj_5048, n2480, n39_adj_5049, 
        n2490, n19, n23_adj_5050, n21_adj_5051, n66309, n31_adj_5052, 
        n29_adj_5053, n66305, n37_adj_5054, n35_adj_5055, n33_adj_5056, 
        n68075, n2491, n18, n41_adj_5057, n67880, n43_adj_5058, 
        n67881, n66307, n67202, n24_adj_5059, n26_adj_5060, n45, 
        n67105, n22_adj_5061, n30_adj_5062, n20_adj_5063, n66303, 
        n68377, n68378, n68184, n67204, n68006, n67103, n68008, 
        n2488;
    wire [23:0]n8269;
    
    wire n2608, n23_adj_5064, n2607, n25_adj_5065, n2611, n17, n21_adj_5066, 
        n19_adj_5067, n66279, n29_adj_5068, n27_adj_5069, n66273, 
        n35_adj_5070, n33_adj_5071, n31_adj_5072, n68069, n2612, n16, 
        n39_adj_5073, n67874, n41_adj_5074, n67875, n66275, n67174, 
        n22_adj_5075, n68009, n43_adj_5076, n67111, n20_adj_5077, 
        n28_adj_5078, n18_adj_5079, n66269, n68379, n68380, n68182, 
        n37_adj_5080, n67178, n68177, n67109, n68478, n2597, n68479, 
        n2730;
    wire [23:0]n8321;
    
    wire n2844, n2843, n15, n2842, n17_adj_5081, n35_adj_5082, n23_adj_5083, 
        n21_adj_5084, n19_adj_5085, n66164, n67130, n67672, n29_adj_5086, 
        n27_adj_5087, n25_adj_5088, n67658, n33_adj_5089, n31_adj_5090, 
        n66166, n2845, n12_adj_5091, n68141, n20_adj_5092, n43_adj_5093, 
        n38_adj_5094, n37_adj_5095, n68142, n41_adj_5096, n39_adj_5097, 
        n66159, n18_adj_5098, n66157, n68139, n68016, n16_adj_5099, 
        n24_adj_5100, n14_adj_5101, n66178, n68454, n68455, n68342, 
        n67978, n68444, n68270, n68586, n2828, n68587, n2728;
    wire [23:0]n8347;
    
    wire n2953, n17_adj_5102, n2952, n19_adj_5103, n2951, n21_adj_5104, 
        n2945, n33_adj_5105, n66123, n15_adj_5106, n13, n2956, n67032, 
        n67646, n27_adj_5107, n25_adj_5108, n23_adj_5109, n67644, 
        n31_adj_5110, n29_adj_5111, n66125, n2957, n10_adj_5112, n68137, 
        n35_adj_5113, n68138, n18_adj_5114, n41_adj_5115, n36, n39_adj_5116, 
        n37_adj_5117, n66108, n16_adj_5118, n66105, n68458, n68022, 
        n14_adj_5119, n22_adj_5120, n12_adj_5121, n66138, n68456, 
        n68457, n68338, n67952, n68576, n68274, n68606, n2940, 
        n68607, n2939, n68601, n2954;
    wire [23:0]n8373;
    
    wire n3062, n3061, n15_adj_5122, n17_adj_5123, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n3060, n19_adj_5124, n3054, n31_adj_5125, r_Rx_Data_R, n66053, 
        n13_adj_5126, n11, n3065, n66972, n67622, n25_adj_5127, 
        n23_adj_5128, n21_adj_5129, n67616, n29_adj_5130, n27_adj_5131, 
        n66055, n3066, n8_adj_5132, n68131, n33_adj_5133, n68132, 
        n16_adj_5134, n39_adj_5135, n34_adj_5136, n37_adj_5137, n35_adj_5138, 
        n66043, n14_adj_5139, n66032, n68460, n68028, n10_adj_5140, 
        n68133, n68134, n66065, n66956, n12_adj_5141, n20_adj_5142, 
        n25657, n58469, n26_adj_5143, n67938, n68578, n67674, n68604, 
        n3049, n68605, n3048, n68595, n3047, n67676, n2938, n3046, 
        n3186;
    wire [23:0]n8399;
    
    wire n61094, n61100, n62276, n62278, n62114, n62274, n58437, 
        n6, n61046, n61052, n62864, n58487, n65654, n65651, n61126, 
        n61132, n3165, n3169, n16_adj_5147, n49674, n49673, n60642, 
        n2723, n2727, n66219, n18_adj_5148, n62906, n49672, n60742, 
        n2725, n20_adj_5149, n2715, n2724, n66196, n49671;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n22_adj_5150, n49670, n60740, n62840, n48_adj_5151, n62870, 
        n48_adj_5152, n1552;
    wire [23:0]n8087;
    
    wire n1553, n1554, n43_adj_5153, n1557, n37_adj_5154, n1556, 
        n39_adj_5155, n1555, n41_adj_5156, n1560, n1558, n1559, 
        n62158, n62144, n62146, n62134, n61998, n58481, n32_adj_5157, 
        n67918, n67919, n66423, n67320, n49669, n60738, n34_adj_5158, 
        n67996, n58495, n67066, n68219, n68220, n49668, n49667, 
        n60736, n69846, n57075, n65670, n65667, n65664;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n29178, n60766, n60772, n27797, n62030, n62806, n49666, 
        n60734, n60700, n3172, n49665, n60640, n62748, n25666, 
        n49664, n60732, n60660, n62752, n61332, n25682, n65705, 
        n48_adj_5159, n65985, n60698;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]n479;
    
    wire n62010, n62012;
    wire [7:0]n1;
    
    wire n50920, n50919, n50918, n50917, n50916, n50915, n50914, 
        n62868, n49663;
    wire [23:0]n8425;
    
    wire n50760, n3082, n50759, n3188, n50758, n3084, n50757, 
        n2977, n50756, n3156, n2867, n50755, n3157, n2754, n50754, 
        n3158, n2638, n50753, n3159, n2519, n50752, n3160, n2397, 
        n50751, n3161, n2272, n50750, n3162, n2144, n50749, n3163, 
        n2013, n50748, n3164, n1879, n50747, n1742, n50746, n3166, 
        n1602, n50745, n3167, n1459, n50744, n3168, n1460, n50743, 
        n1011, n50742, n3170, n856, n50741, n3171, n698, n50740, 
        n858, n50739, n60702, n538, n50738, n50737, n50736, n50735, 
        n50734, n3050, n50733, n3051, n50732, n3052, n50731, n3053, 
        n50730, n50729, n3055, n50728, n3056, n50727, n3057, n50726, 
        n3058, n50725, n3059, n50724, n50723, n50722, n50721, 
        n3063, n50720, n3064, n50719, n50718, n50717, n58441, 
        n50716, n50715, n50714, n2941, n50713, n2942, n50712, 
        n2943, n50711, n2944, n50710, n50709, n2946, n50708, n2947, 
        n50707, n2948, n50706, n2949, n50705, n2950, n50704, n50703, 
        n50702, n50701, n50700, n2955, n50699, n50698, n50697, 
        n58445, n2827, n50696, n50695, n2829, n50694, n2830, n50693, 
        n2831, n50692, n2832, n50691, n2833, n50690, n2834, n50689, 
        n49662, n2835, n50688, n2836, n50687, n2837, n50686, n2838, 
        n50685, n2839, n50684, n2840, n50683, n2841, n50682, n50681, 
        n50680, n50679, n50678, n49661, n60696, n58449, n2713, 
        n50677, n2714, n50676, n50675, n2716, n50674, n2717, n50673, 
        n2718, n50672, n2719, n50671, n2720, n50670, n2721, n50669, 
        n2722, n50668, n50667, n50666, n50665, n2726, n50664, 
        n50663, n50662, n2729, n50661, n50660, n60694, n58453;
    wire [23:0]n8295;
    
    wire n2596, n50659, n50658, n2598, n50657, n2599, n50656, 
        n2600, n50655, n2601, n50654, n2602, n50653, n49660, n2603, 
        n50652, n2604, n50651, n2605, n50650, n2606, n50649, n50648, 
        n50647, n3_adj_5166, n2609, n50646, n2610, n50645, n50644, 
        n50643, n60692, n58457, n2476, n50642, n2477, n50641, 
        n2478, n50640, n2479, n50639, n50638, n2481, n50637, n2482, 
        n50636, n2483, n50635, n2484, n50634, n2485, n50633, n50632, 
        n50631, n50630, n2489, n50629, n50628, n50627, n60690, 
        n58461, n2353, n50626, n50625, n50624, n2356, n50623, 
        n2357, n50622, n2358, n50621, n2359, n50620, n2360, n50619, 
        n2361, n50618, n50617, n50616, n50615, n50614, n50613, 
        n50612, n60688, n58465, n50611, n50610, n50609, n50608, 
        n50607, n50606, n50605, n50604, n50603, n50602, n50601, 
        n50600, n50599, n50598, n60686, n50597, n50596, n50595, 
        n50594, n50593, n50592, n50591, n50590, n50589, n50588, 
        n50587, n50586, n50585, n50584, n50583, n50582, n50581, 
        n50580, n50579, n50578, n50577, n50576, n50575, n50574, 
        n50573, n50572, n50571, n50570, n50569, n50568, n50567, 
        n50566, n50565, n50564, n50563, n60684, n58478, n50562, 
        n50561, n50560, n50559, n50558, n50557, n49659, n50556, 
        n50555, n50554, n50553, n50552, n50551, n50550, n50549, 
        n50548, n50547, n50546, n50545, n25663;
    wire [23:0]n8061;
    
    wire n1408, n50544, n1409, n50543, n1410, n50542, n1411, n50541, 
        n1412, n50540, n1413, n50539, n1414, n50538, n1415, n50537, 
        n60682;
    wire [23:0]n8035;
    
    wire n1261, n50536, n1262, n50535, n60748, n1263, n50534, 
        n1264, n50533, n49658, n1265, n50532, n1266, n50531, n1267, 
        n50530, n60680, n58491;
    wire [23:0]n8009;
    
    wire n1111, n50529, n1112, n50528, n1113, n50527, n1114, n50526, 
        n1115, n50525, n1116, n50524, n60678, n49657, n49656, 
        n49655, n49654, n49653, n49652, n49651, n59626, n62648, 
        n60115, n48_adj_5168, n25692, n65987, n44_adj_5169, n62602, 
        n805, n42_adj_5170, n20994, n43_adj_5171, n37_adj_5172, n41_adj_5173, 
        n39_adj_5174, n962, n48_adj_5175, n25605, n961, n42_adj_5176, 
        n32_adj_5177, n67920, n67921, n66435, n67330, n34_adj_5178, 
        n67994, n67063, n11428, n68221, n68222, n43_adj_5179, n45_adj_5180, 
        n41_adj_5181, n39_adj_5182, n34_adj_5183, n67924, n67925, 
        n66445, n67338, n36_adj_5184, n38_adj_5185, n67059, n67988, 
        n65682, n65688, n65679, n65685, n41_adj_5186, n36_adj_5187, 
        n38_adj_5188, n40_adj_5189, n66452, n68361, n68362, n68224, 
        n68428, n25660, n14_adj_5190, n15_adj_5191, n61158, n61164, 
        n61142, n61148, n61078, n61084, n60714, n959, n58926, 
        n44_adj_5192, n46, n58193, n40_adj_5193, n960, n21004, n21006, 
        n43_adj_5194, n38_adj_5195, n40_adj_5196, n42_adj_5197, n66458, 
        n68349, n68350, n803, n58972, n44_adj_5198, n46_adj_5199, 
        n58191, n804, n42960, n20996, n62162, n62164, n62160, 
        n62020, n58498, n42_adj_5200, n67928, n67929, n25670, n60672, 
        n61774, n3_adj_5201, n61778, n61062, n61068, n5, n61110, 
        n61116, n58189, n61782, n8_adj_5202, n68641, n62866, n42_adj_5203, 
        n67930, n67931, n60806, n60812, n62782, n62888, n2, n11645, 
        n61274, n58984, n59856, n65628, n58258, n61328, n65629, 
        n62272, n61008, n62826, n61036, n62586, n62896, n62884, 
        n61356, n62004, n62002, n62000, n61340, n46_adj_5204, n62762, 
        n42962, n60658, n62788, n60618, n62838, n60952, n60970, 
        n62832, n62898, n4, n62112, n62808, n62584, n61192, n61188, 
        n61190, n61186, n62902, n41_adj_5205, n39_adj_5206, n35_adj_5207, 
        n37_adj_5208, n29_adj_5209, n31_adj_5210, n23_adj_5211, n25_adj_5212, 
        n33_adj_5213, n7, n43_adj_5214, n45_adj_5215, n9, n17_adj_5216, 
        n19_adj_5217, n21_adj_5218, n11_adj_5219, n61196, n13_adj_5220, 
        n15_adj_5221, n27_adj_5222, n62118, n65923, n61234, n62650, 
        n65931, n16_adj_5223, n61194, n61208, n61210, n65892, n8_adj_5224, 
        n24_adj_5225, n3274, n65945, n66819, n66815, n68179, n67558, 
        n68398, n12_adj_5226, n4_adj_5227, n68113, n68114, n65913, 
        n10_adj_5228, n30_adj_5229, n65915, n41_adj_5230, n45_adj_5231, 
        n68464, n39_adj_5232, n43_adj_5233, n68044, n68582, n68583, 
        n33_adj_5234, n35_adj_5235, n6_adj_5236, n27_adj_5237, n29_adj_5238, 
        n31_adj_5239, n68117, n68118, n17_adj_5240, n19_adj_5241, 
        n65897, n67680, n21_adj_5242, n23_adj_5243, n25_adj_5244, 
        n37_adj_5245, n68042, n66204, n67164, n68524, n65899, n67702, 
        n67698, n66206, n68283, n14_adj_5246, n67868, n40_adj_5247, 
        n67869, n40_adj_5248, n66200, n68011, n60630, n67123, n3253, 
        n26_adj_5249, n68285, n68381, n68382, n68176, n60638, n68053, 
        n68426, n67121, n9_adj_5250, n11_adj_5251, n19_adj_5252, n13_adj_5253, 
        n15_adj_5254, n17_adj_5255, n29_adj_5256, n66910, n67594, 
        n67592, n6_adj_5257;
    
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8217[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8191[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8217[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8191[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8191[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14), .I1(baudrate[17]), 
            .I2(n37), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52396_3_lut (.I0(n68123), .I1(baudrate[14]), .I2(n31), .I3(GND_net), 
            .O(n68124));   // verilog/uart_rx.v(119[33:55])
    defparam i52396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50239_4_lut (.I0(n35), .I1(n33), .I2(n31), .I3(n65973), 
            .O(n65967));
    defparam i50239_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52734_4_lut (.I0(n32), .I1(n12), .I2(n37), .I3(n65958), 
            .O(n68462));   // verilog/uart_rx.v(119[33:55])
    defparam i52734_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52306_3_lut (.I0(n68124), .I1(baudrate[15]), .I2(n33), .I3(GND_net), 
            .O(n68034));   // verilog/uart_rx.v(119[33:55])
    defparam i52306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8191[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8191[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8191[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4987));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(n25645), .I1(n48), .I2(baudrate[0]), .I3(GND_net), 
            .O(n2240));
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8191[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52397_3_lut (.I0(n8), .I1(baudrate[10]), .I2(n23_c), .I3(GND_net), 
            .O(n68125));   // verilog/uart_rx.v(119[33:55])
    defparam i52397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52398_3_lut (.I0(n68125), .I1(baudrate[11]), .I2(n25), .I3(GND_net), 
            .O(n68126));   // verilog/uart_rx.v(119[33:55])
    defparam i52398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51170_4_lut (.I0(n25), .I1(n23_c), .I2(n21), .I3(n65993), 
            .O(n66898));
    defparam i51170_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51950_3_lut (.I0(n10), .I1(baudrate[9]), .I2(n21), .I3(GND_net), 
            .O(n67678));   // verilog/uart_rx.v(119[33:55])
    defparam i51950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8191[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8191[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4988));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4989));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4990));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52304_3_lut (.I0(n68126), .I1(baudrate[12]), .I2(n27_c), 
            .I3(GND_net), .O(n68032));   // verilog/uart_rx.v(119[33:55])
    defparam i52304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8165[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52164_4_lut (.I0(n35), .I1(n33), .I2(n31), .I3(n65980), 
            .O(n67892));
    defparam i52164_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8165[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52852_4_lut (.I0(n68034), .I1(n68462), .I2(n37), .I3(n65967), 
            .O(n68580));   // verilog/uart_rx.v(119[33:55])
    defparam i52852_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52391_4_lut (.I0(n68032), .I1(n67678), .I2(n27_c), .I3(n66898), 
            .O(n68119));   // verilog/uart_rx.v(119[33:55])
    defparam i52391_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52874_4_lut (.I0(n68119), .I1(n68580), .I2(n37), .I3(n67892), 
            .O(n68602));   // verilog/uart_rx.v(119[33:55])
    defparam i52874_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52875_3_lut (.I0(n68602), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n68603));   // verilog/uart_rx.v(119[33:55])
    defparam i52875_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8165[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8165[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52871_3_lut (.I0(n68603), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n68599));   // verilog/uart_rx.v(119[33:55])
    defparam i52871_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4991));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8165[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52666_3_lut (.I0(n68599), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n68394));   // verilog/uart_rx.v(119[33:55])
    defparam i52666_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52667_3_lut (.I0(n68394), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n68395));   // verilog/uart_rx.v(119[33:55])
    defparam i52667_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4992));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8165[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8165[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52312_3_lut (.I0(n68395), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_4993));   // verilog/uart_rx.v(119[33:55])
    defparam i52312_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4994));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8165[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4995));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8165[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8165[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4996));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4997));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4998));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n62168));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_983 (.I0(n62116), .I1(n62166), .I2(n61214), .I3(GND_net), 
            .O(n62176));
    defparam i1_3_lut_adj_983.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_984 (.I0(n62176), .I1(n62172), .I2(n62174), .I3(n62168), 
            .O(n25645));
    defparam i1_4_lut_adj_984.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4999));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50643_4_lut (.I0(n33_adj_4998), .I1(n31_adj_4997), .I2(n29_adj_4996), 
            .I3(n27_adj_4999), .O(n66371));
    defparam i50643_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30), .I1(baudrate[10]), 
            .I2(n41_adj_4994), .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29021_rep_4_2_lut (.I0(n8165[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n58472));   // verilog/uart_rx.v(119[33:55])
    defparam i29021_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n58472), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52166_3_lut (.I0(n26), .I1(baudrate[6]), .I2(n33_adj_4998), 
            .I3(GND_net), .O(n67894));   // verilog/uart_rx.v(119[33:55])
    defparam i52166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52167_3_lut (.I0(n67894), .I1(baudrate[7]), .I2(n35_adj_4992), 
            .I3(GND_net), .O(n67895));   // verilog/uart_rx.v(119[33:55])
    defparam i52167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50637_4_lut (.I0(n39_adj_4995), .I1(n37_adj_4991), .I2(n35_adj_4992), 
            .I3(n66371), .O(n66365));
    defparam i50637_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52643_4_lut (.I0(n38), .I1(n28), .I2(n41_adj_4994), .I3(n66363), 
            .O(n68371));   // verilog/uart_rx.v(119[33:55])
    defparam i52643_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51355_3_lut (.I0(n67895), .I1(baudrate[8]), .I2(n37_adj_4991), 
            .I3(GND_net), .O(n67083));   // verilog/uart_rx.v(119[33:55])
    defparam i51355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52817_4_lut (.I0(n67083), .I1(n68371), .I2(n41_adj_4994), 
            .I3(n66365), .O(n68545));   // verilog/uart_rx.v(119[33:55])
    defparam i52817_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52818_3_lut (.I0(n68545), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n68546));   // verilog/uart_rx.v(119[33:55])
    defparam i52818_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52755_3_lut (.I0(n68546), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n68483));   // verilog/uart_rx.v(119[33:55])
    defparam i52755_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51361_3_lut (.I0(n68483), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i51361_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8165[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8191[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8139[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8139[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8139[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8139[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8139[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8139[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5000));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5001));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8139[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5002));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8139[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5003));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8113[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8113[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8113[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5004));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8113[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5005));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_985 (.I0(n25636), .I1(n48_adj_5006), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_985.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8113[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5007));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8113[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5008));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8113[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8113[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5009));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5010));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8113[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5012));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50680_4_lut (.I0(n35_adj_5011), .I1(n33_adj_5010), .I2(n31_adj_5009), 
            .I3(n29_adj_5012), .O(n66408));
    defparam i50680_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5013), .I1(baudrate[9]), 
            .I2(n43_adj_5007), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5014));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52188_3_lut (.I0(n28_adj_5014), .I1(baudrate[5]), .I2(n35_adj_5011), 
            .I3(GND_net), .O(n67916));   // verilog/uart_rx.v(119[33:55])
    defparam i52188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52189_3_lut (.I0(n67916), .I1(baudrate[6]), .I2(n37_adj_5005), 
            .I3(GND_net), .O(n67917));   // verilog/uart_rx.v(119[33:55])
    defparam i52189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50672_4_lut (.I0(n41_adj_5008), .I1(n39_adj_5004), .I2(n37_adj_5005), 
            .I3(n66408), .O(n66400));
    defparam i50672_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52619_4_lut (.I0(n40), .I1(n30_adj_5015), .I2(n43_adj_5007), 
            .I3(n66398), .O(n68347));   // verilog/uart_rx.v(119[33:55])
    defparam i52619_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51343_3_lut (.I0(n67917), .I1(baudrate[7]), .I2(n39_adj_5004), 
            .I3(GND_net), .O(n67071));   // verilog/uart_rx.v(119[33:55])
    defparam i51343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52805_4_lut (.I0(n67071), .I1(n68347), .I2(n43_adj_5007), 
            .I3(n66400), .O(n68533));   // verilog/uart_rx.v(119[33:55])
    defparam i52805_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52806_3_lut (.I0(n68533), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n68534));   // verilog/uart_rx.v(119[33:55])
    defparam i52806_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8113[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8139[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8139[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5016));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5017));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5018));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5019));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50662_4_lut (.I0(n33_adj_5018), .I1(n31_adj_5017), .I2(n29_adj_5016), 
            .I3(n27_adj_5019), .O(n66390));
    defparam i50662_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5020), .I1(baudrate[9]), 
            .I2(n41_adj_5002), .I3(GND_net), .O(n38_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52184_3_lut (.I0(n26_adj_5022), .I1(baudrate[5]), .I2(n33_adj_5018), 
            .I3(GND_net), .O(n67912));   // verilog/uart_rx.v(119[33:55])
    defparam i52184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52185_3_lut (.I0(n67912), .I1(baudrate[6]), .I2(n35_adj_5000), 
            .I3(GND_net), .O(n67913));   // verilog/uart_rx.v(119[33:55])
    defparam i52185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50655_4_lut (.I0(n39_adj_5003), .I1(n37_adj_5001), .I2(n35_adj_5000), 
            .I3(n66390), .O(n66383));
    defparam i50655_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52641_4_lut (.I0(n38_adj_5021), .I1(n28_adj_5023), .I2(n41_adj_5002), 
            .I3(n66381), .O(n68369));   // verilog/uart_rx.v(119[33:55])
    defparam i52641_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51347_3_lut (.I0(n67913), .I1(baudrate[7]), .I2(n37_adj_5001), 
            .I3(GND_net), .O(n67075));   // verilog/uart_rx.v(119[33:55])
    defparam i51347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52815_4_lut (.I0(n67075), .I1(n68369), .I2(n41_adj_5002), 
            .I3(n66383), .O(n68543));   // verilog/uart_rx.v(119[33:55])
    defparam i52815_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52816_3_lut (.I0(n68543), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n68544));   // verilog/uart_rx.v(119[33:55])
    defparam i52816_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52757_3_lut (.I0(n68544), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n68485));   // verilog/uart_rx.v(119[33:55])
    defparam i52757_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51353_3_lut (.I0(n68485), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam i51353_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8139[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8165[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8191[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8191[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50625_4_lut (.I0(n29_adj_5027), .I1(n27_adj_5026), .I2(n25_adj_5025), 
            .I3(n23_adj_5028), .O(n66353));
    defparam i50625_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50620_4_lut (.I0(n35_adj_4990), .I1(n33_adj_4989), .I2(n31_adj_4988), 
            .I3(n66353), .O(n66348));
    defparam i50620_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5029), .I1(baudrate[7]), 
            .I2(n33_adj_4989), .I3(GND_net), .O(n30_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5031), .I1(baudrate[9]), 
            .I2(n37_adj_4987), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52645_4_lut (.I0(n34), .I1(n24), .I2(n37_adj_4987), .I3(n66346), 
            .O(n68373));   // verilog/uart_rx.v(119[33:55])
    defparam i52645_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52646_3_lut (.I0(n68373), .I1(baudrate[10]), .I2(n39), .I3(GND_net), 
            .O(n68374));   // verilog/uart_rx.v(119[33:55])
    defparam i52646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52462_3_lut (.I0(n68374), .I1(baudrate[11]), .I2(n41), .I3(GND_net), 
            .O(n68190));   // verilog/uart_rx.v(119[33:55])
    defparam i52462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52351_4_lut (.I0(n41), .I1(n39), .I2(n37_adj_4987), .I3(n66348), 
            .O(n68079));
    defparam i52351_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52419_4_lut (.I0(n30_adj_5030), .I1(n22), .I2(n33_adj_4989), 
            .I3(n66350), .O(n68147));   // verilog/uart_rx.v(119[33:55])
    defparam i52419_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51365_3_lut (.I0(n68190), .I1(baudrate[12]), .I2(n43), .I3(GND_net), 
            .O(n67093));   // verilog/uart_rx.v(119[33:55])
    defparam i51365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52617_4_lut (.I0(n67093), .I1(n68147), .I2(n43), .I3(n68079), 
            .O(n68345));   // verilog/uart_rx.v(119[33:55])
    defparam i52617_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52618_3_lut (.I0(n68345), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n68346));   // verilog/uart_rx.v(119[33:55])
    defparam i52618_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8191[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8217[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8217[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50604_4_lut (.I0(n27_adj_5034), .I1(n25_adj_5033), .I2(n23_adj_5032), 
            .I3(n21_adj_5035), .O(n66332));
    defparam i50604_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50597_4_lut (.I0(n33_adj_5036), .I1(n31_adj_5037), .I2(n29_c), 
            .I3(n66332), .O(n66325));
    defparam i50597_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5038), .I1(baudrate[7]), 
            .I2(n31_adj_5037), .I3(GND_net), .O(n28_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5040), .I1(baudrate[9]), 
            .I2(n35_adj_5041), .I3(GND_net), .O(n32_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52647_4_lut (.I0(n32_adj_5042), .I1(n22_adj_5043), .I2(n35_adj_5041), 
            .I3(n66323), .O(n68375));   // verilog/uart_rx.v(119[33:55])
    defparam i52647_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52648_3_lut (.I0(n68375), .I1(baudrate[10]), .I2(n37_adj_5044), 
            .I3(GND_net), .O(n68376));   // verilog/uart_rx.v(119[33:55])
    defparam i52648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52458_3_lut (.I0(n68376), .I1(baudrate[11]), .I2(n39_adj_5045), 
            .I3(GND_net), .O(n68186));   // verilog/uart_rx.v(119[33:55])
    defparam i52458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52349_4_lut (.I0(n39_adj_5045), .I1(n37_adj_5044), .I2(n35_adj_5041), 
            .I3(n66325), .O(n68077));
    defparam i52349_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52724_4_lut (.I0(n28_adj_5039), .I1(n20), .I2(n31_adj_5037), 
            .I3(n66329), .O(n68452));   // verilog/uart_rx.v(119[33:55])
    defparam i52724_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51371_3_lut (.I0(n68186), .I1(baudrate[12]), .I2(n41_adj_5046), 
            .I3(GND_net), .O(n67099));   // verilog/uart_rx.v(119[33:55])
    defparam i51371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52791_4_lut (.I0(n67099), .I1(n68452), .I2(n41_adj_5046), 
            .I3(n68077), .O(n68519));   // verilog/uart_rx.v(119[33:55])
    defparam i52791_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52792_3_lut (.I0(n68519), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n68520));   // verilog/uart_rx.v(119[33:55])
    defparam i52792_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52719_3_lut (.I0(n68520), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n68447));   // verilog/uart_rx.v(119[33:55])
    defparam i52719_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8217[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8243[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8243[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50581_4_lut (.I0(n25_adj_5047), .I1(n23_adj_5050), .I2(n21_adj_5051), 
            .I3(n19), .O(n66309));
    defparam i50581_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50577_4_lut (.I0(n31_adj_5052), .I1(n29_adj_5053), .I2(n27_adj_5048), 
            .I3(n66309), .O(n66305));
    defparam i50577_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52347_4_lut (.I0(n37_adj_5054), .I1(n35_adj_5055), .I2(n33_adj_5056), 
            .I3(n66305), .O(n68075));
    defparam i52347_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52152_3_lut (.I0(n18), .I1(baudrate[13]), .I2(n41_adj_5057), 
            .I3(GND_net), .O(n67880));   // verilog/uart_rx.v(119[33:55])
    defparam i52152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52153_3_lut (.I0(n67880), .I1(baudrate[14]), .I2(n43_adj_5058), 
            .I3(GND_net), .O(n67881));   // verilog/uart_rx.v(119[33:55])
    defparam i52153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51474_4_lut (.I0(n43_adj_5058), .I1(n41_adj_5057), .I2(n29_adj_5053), 
            .I3(n66307), .O(n67202));
    defparam i51474_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5059), .I1(baudrate[7]), 
            .I2(n29_adj_5053), .I3(GND_net), .O(n26_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51377_3_lut (.I0(n67881), .I1(baudrate[15]), .I2(n45), .I3(GND_net), 
            .O(n67105));   // verilog/uart_rx.v(119[33:55])
    defparam i51377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5061), .I1(baudrate[9]), 
            .I2(n33_adj_5056), .I3(GND_net), .O(n30_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52649_4_lut (.I0(n30_adj_5062), .I1(n20_adj_5063), .I2(n33_adj_5056), 
            .I3(n66303), .O(n68377));   // verilog/uart_rx.v(119[33:55])
    defparam i52649_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52650_3_lut (.I0(n68377), .I1(baudrate[10]), .I2(n35_adj_5055), 
            .I3(GND_net), .O(n68378));   // verilog/uart_rx.v(119[33:55])
    defparam i52650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52456_3_lut (.I0(n68378), .I1(baudrate[11]), .I2(n37_adj_5054), 
            .I3(GND_net), .O(n68184));   // verilog/uart_rx.v(119[33:55])
    defparam i52456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51476_4_lut (.I0(n43_adj_5058), .I1(n41_adj_5057), .I2(n39_adj_5049), 
            .I3(n68075), .O(n67204));
    defparam i51476_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52278_4_lut (.I0(n67105), .I1(n26_adj_5060), .I2(n45), .I3(n67202), 
            .O(n68006));   // verilog/uart_rx.v(119[33:55])
    defparam i52278_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51375_3_lut (.I0(n68184), .I1(baudrate[12]), .I2(n39_adj_5049), 
            .I3(GND_net), .O(n67103));   // verilog/uart_rx.v(119[33:55])
    defparam i51375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52280_4_lut (.I0(n67103), .I1(n68006), .I2(n45), .I3(n67204), 
            .O(n68008));   // verilog/uart_rx.v(119[33:55])
    defparam i52280_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8243[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8269[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50551_4_lut (.I0(n23_adj_5064), .I1(n21_adj_5066), .I2(n19_adj_5067), 
            .I3(n17), .O(n66279));
    defparam i50551_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50545_4_lut (.I0(n29_adj_5068), .I1(n27_adj_5069), .I2(n25_adj_5065), 
            .I3(n66279), .O(n66273));
    defparam i50545_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52341_4_lut (.I0(n35_adj_5070), .I1(n33_adj_5071), .I2(n31_adj_5072), 
            .I3(n66273), .O(n68069));
    defparam i52341_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52146_3_lut (.I0(n16), .I1(baudrate[13]), .I2(n39_adj_5073), 
            .I3(GND_net), .O(n67874));   // verilog/uart_rx.v(119[33:55])
    defparam i52146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52147_3_lut (.I0(n67874), .I1(baudrate[14]), .I2(n41_adj_5074), 
            .I3(GND_net), .O(n67875));   // verilog/uart_rx.v(119[33:55])
    defparam i52147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51446_4_lut (.I0(n41_adj_5074), .I1(n39_adj_5073), .I2(n27_adj_5069), 
            .I3(n66275), .O(n67174));
    defparam i51446_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52281_3_lut (.I0(n22_adj_5075), .I1(baudrate[7]), .I2(n27_adj_5069), 
            .I3(GND_net), .O(n68009));   // verilog/uart_rx.v(119[33:55])
    defparam i52281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51383_3_lut (.I0(n67875), .I1(baudrate[15]), .I2(n43_adj_5076), 
            .I3(GND_net), .O(n67111));   // verilog/uart_rx.v(119[33:55])
    defparam i51383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5077), .I1(baudrate[9]), 
            .I2(n31_adj_5072), .I3(GND_net), .O(n28_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52651_4_lut (.I0(n28_adj_5078), .I1(n18_adj_5079), .I2(n31_adj_5072), 
            .I3(n66269), .O(n68379));   // verilog/uart_rx.v(119[33:55])
    defparam i52651_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52652_3_lut (.I0(n68379), .I1(baudrate[10]), .I2(n33_adj_5071), 
            .I3(GND_net), .O(n68380));   // verilog/uart_rx.v(119[33:55])
    defparam i52652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52454_3_lut (.I0(n68380), .I1(baudrate[11]), .I2(n35_adj_5070), 
            .I3(GND_net), .O(n68182));   // verilog/uart_rx.v(119[33:55])
    defparam i52454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51450_4_lut (.I0(n41_adj_5074), .I1(n39_adj_5073), .I2(n37_adj_5080), 
            .I3(n68069), .O(n67178));
    defparam i51450_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52449_4_lut (.I0(n67111), .I1(n68009), .I2(n43_adj_5076), 
            .I3(n67174), .O(n68177));   // verilog/uart_rx.v(119[33:55])
    defparam i52449_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51381_3_lut (.I0(n68182), .I1(baudrate[12]), .I2(n37_adj_5080), 
            .I3(GND_net), .O(n67109));   // verilog/uart_rx.v(119[33:55])
    defparam i51381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52750_4_lut (.I0(n67109), .I1(n68177), .I2(n43_adj_5076), 
            .I3(n67178), .O(n68478));   // verilog/uart_rx.v(119[33:55])
    defparam i52750_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52751_3_lut (.I0(n68478), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n68479));   // verilog/uart_rx.v(119[33:55])
    defparam i52751_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8321[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50436_4_lut (.I0(n35_adj_5082), .I1(n23_adj_5083), .I2(n21_adj_5084), 
            .I3(n19_adj_5085), .O(n66164));
    defparam i50436_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51402_4_lut (.I0(n17_adj_5081), .I1(n15), .I2(n2844), .I3(baudrate[2]), 
            .O(n67130));
    defparam i51402_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51944_4_lut (.I0(n23_adj_5083), .I1(n21_adj_5084), .I2(n19_adj_5085), 
            .I3(n67130), .O(n67672));
    defparam i51944_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51930_4_lut (.I0(n29_adj_5086), .I1(n27_adj_5087), .I2(n25_adj_5088), 
            .I3(n67672), .O(n67658));
    defparam i51930_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50438_4_lut (.I0(n35_adj_5082), .I1(n33_adj_5089), .I2(n31_adj_5090), 
            .I3(n67658), .O(n66166));
    defparam i50438_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52413_3_lut (.I0(n12_adj_5091), .I1(baudrate[13]), .I2(n35_adj_5082), 
            .I3(GND_net), .O(n68141));   // verilog/uart_rx.v(119[33:55])
    defparam i52413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5092), .I1(baudrate[17]), 
            .I2(n43_adj_5093), .I3(GND_net), .O(n38_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52414_3_lut (.I0(n68141), .I1(baudrate[14]), .I2(n37_adj_5095), 
            .I3(GND_net), .O(n68142));   // verilog/uart_rx.v(119[33:55])
    defparam i52414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50431_4_lut (.I0(n41_adj_5096), .I1(n39_adj_5097), .I2(n37_adj_5095), 
            .I3(n66164), .O(n66159));
    defparam i50431_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52411_4_lut (.I0(n38_adj_5094), .I1(n18_adj_5098), .I2(n43_adj_5093), 
            .I3(n66157), .O(n68139));   // verilog/uart_rx.v(119[33:55])
    defparam i52411_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52288_3_lut (.I0(n68142), .I1(baudrate[15]), .I2(n39_adj_5097), 
            .I3(GND_net), .O(n68016));   // verilog/uart_rx.v(119[33:55])
    defparam i52288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5099), .I1(baudrate[9]), 
            .I2(n27_adj_5087), .I3(GND_net), .O(n24_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52726_4_lut (.I0(n24_adj_5100), .I1(n14_adj_5101), .I2(n27_adj_5087), 
            .I3(n66178), .O(n68454));   // verilog/uart_rx.v(119[33:55])
    defparam i52726_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52727_3_lut (.I0(n68454), .I1(baudrate[10]), .I2(n29_adj_5086), 
            .I3(GND_net), .O(n68455));   // verilog/uart_rx.v(119[33:55])
    defparam i52727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52614_3_lut (.I0(n68455), .I1(baudrate[11]), .I2(n31_adj_5090), 
            .I3(GND_net), .O(n68342));   // verilog/uart_rx.v(119[33:55])
    defparam i52614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52250_4_lut (.I0(n41_adj_5096), .I1(n39_adj_5097), .I2(n37_adj_5095), 
            .I3(n66166), .O(n67978));
    defparam i52250_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52716_4_lut (.I0(n68016), .I1(n68139), .I2(n43_adj_5093), 
            .I3(n66159), .O(n68444));   // verilog/uart_rx.v(119[33:55])
    defparam i52716_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52542_3_lut (.I0(n68342), .I1(baudrate[12]), .I2(n33_adj_5089), 
            .I3(GND_net), .O(n68270));   // verilog/uart_rx.v(119[33:55])
    defparam i52542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52858_4_lut (.I0(n68270), .I1(n68444), .I2(n43_adj_5093), 
            .I3(n67978), .O(n68586));   // verilog/uart_rx.v(119[33:55])
    defparam i52858_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52859_3_lut (.I0(n68586), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n68587));   // verilog/uart_rx.v(119[33:55])
    defparam i52859_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8321[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8347[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50395_4_lut (.I0(n33_adj_5105), .I1(n21_adj_5104), .I2(n19_adj_5103), 
            .I3(n17_adj_5102), .O(n66123));
    defparam i50395_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51304_4_lut (.I0(n15_adj_5106), .I1(n13), .I2(n2956), .I3(baudrate[2]), 
            .O(n67032));
    defparam i51304_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51918_4_lut (.I0(n21_adj_5104), .I1(n19_adj_5103), .I2(n17_adj_5102), 
            .I3(n67032), .O(n67646));
    defparam i51918_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51916_4_lut (.I0(n27_adj_5107), .I1(n25_adj_5108), .I2(n23_adj_5109), 
            .I3(n67646), .O(n67644));
    defparam i51916_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50397_4_lut (.I0(n33_adj_5105), .I1(n31_adj_5110), .I2(n29_adj_5111), 
            .I3(n67644), .O(n66125));
    defparam i50397_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52409_3_lut (.I0(n10_adj_5112), .I1(baudrate[13]), .I2(n33_adj_5105), 
            .I3(GND_net), .O(n68137));   // verilog/uart_rx.v(119[33:55])
    defparam i52409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52410_3_lut (.I0(n68137), .I1(baudrate[14]), .I2(n35_adj_5113), 
            .I3(GND_net), .O(n68138));   // verilog/uart_rx.v(119[33:55])
    defparam i52410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5114), .I1(baudrate[17]), 
            .I2(n41_adj_5115), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50380_4_lut (.I0(n39_adj_5116), .I1(n37_adj_5117), .I2(n35_adj_5113), 
            .I3(n66123), .O(n66108));
    defparam i50380_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52730_4_lut (.I0(n36), .I1(n16_adj_5118), .I2(n41_adj_5115), 
            .I3(n66105), .O(n68458));   // verilog/uart_rx.v(119[33:55])
    defparam i52730_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52294_3_lut (.I0(n68138), .I1(baudrate[15]), .I2(n37_adj_5117), 
            .I3(GND_net), .O(n68022));   // verilog/uart_rx.v(119[33:55])
    defparam i52294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5119), .I1(baudrate[9]), 
            .I2(n25_adj_5108), .I3(GND_net), .O(n22_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52728_4_lut (.I0(n22_adj_5120), .I1(n12_adj_5121), .I2(n25_adj_5108), 
            .I3(n66138), .O(n68456));   // verilog/uart_rx.v(119[33:55])
    defparam i52728_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52729_3_lut (.I0(n68456), .I1(baudrate[10]), .I2(n27_adj_5107), 
            .I3(GND_net), .O(n68457));   // verilog/uart_rx.v(119[33:55])
    defparam i52729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52610_3_lut (.I0(n68457), .I1(baudrate[11]), .I2(n29_adj_5111), 
            .I3(GND_net), .O(n68338));   // verilog/uart_rx.v(119[33:55])
    defparam i52610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52224_4_lut (.I0(n39_adj_5116), .I1(n37_adj_5117), .I2(n35_adj_5113), 
            .I3(n66125), .O(n67952));
    defparam i52224_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52848_4_lut (.I0(n68022), .I1(n68458), .I2(n41_adj_5115), 
            .I3(n66108), .O(n68576));   // verilog/uart_rx.v(119[33:55])
    defparam i52848_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52546_3_lut (.I0(n68338), .I1(baudrate[12]), .I2(n31_adj_5110), 
            .I3(GND_net), .O(n68274));   // verilog/uart_rx.v(119[33:55])
    defparam i52546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52878_4_lut (.I0(n68274), .I1(n68576), .I2(n41_adj_5115), 
            .I3(n67952), .O(n68606));   // verilog/uart_rx.v(119[33:55])
    defparam i52878_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52879_3_lut (.I0(n68606), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n68607));   // verilog/uart_rx.v(119[33:55])
    defparam i52879_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52873_3_lut (.I0(n68607), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n68601));   // verilog/uart_rx.v(119[33:55])
    defparam i52873_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8347[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8373[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8373[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 i50325_4_lut (.I0(n31_adj_5125), .I1(n19_adj_5124), .I2(n17_adj_5123), 
            .I3(n15_adj_5122), .O(n66053));
    defparam i50325_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51244_4_lut (.I0(n13_adj_5126), .I1(n11), .I2(n3065), .I3(baudrate[2]), 
            .O(n66972));
    defparam i51244_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51894_4_lut (.I0(n19_adj_5124), .I1(n17_adj_5123), .I2(n15_adj_5122), 
            .I3(n66972), .O(n67622));
    defparam i51894_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51888_4_lut (.I0(n25_adj_5127), .I1(n23_adj_5128), .I2(n21_adj_5129), 
            .I3(n67622), .O(n67616));
    defparam i51888_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50327_4_lut (.I0(n31_adj_5125), .I1(n29_adj_5130), .I2(n27_adj_5131), 
            .I3(n67616), .O(n66055));
    defparam i50327_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52403_3_lut (.I0(n8_adj_5132), .I1(baudrate[13]), .I2(n31_adj_5125), 
            .I3(GND_net), .O(n68131));   // verilog/uart_rx.v(119[33:55])
    defparam i52403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52404_3_lut (.I0(n68131), .I1(baudrate[14]), .I2(n33_adj_5133), 
            .I3(GND_net), .O(n68132));   // verilog/uart_rx.v(119[33:55])
    defparam i52404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5134), .I1(baudrate[17]), 
            .I2(n39_adj_5135), .I3(GND_net), .O(n34_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50315_4_lut (.I0(n37_adj_5137), .I1(n35_adj_5138), .I2(n33_adj_5133), 
            .I3(n66053), .O(n66043));
    defparam i50315_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52732_4_lut (.I0(n34_adj_5136), .I1(n14_adj_5139), .I2(n39_adj_5135), 
            .I3(n66032), .O(n68460));   // verilog/uart_rx.v(119[33:55])
    defparam i52732_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52300_3_lut (.I0(n68132), .I1(baudrate[15]), .I2(n35_adj_5138), 
            .I3(GND_net), .O(n68028));   // verilog/uart_rx.v(119[33:55])
    defparam i52300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52405_3_lut (.I0(n10_adj_5140), .I1(baudrate[10]), .I2(n25_adj_5127), 
            .I3(GND_net), .O(n68133));   // verilog/uart_rx.v(119[33:55])
    defparam i52405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52406_3_lut (.I0(n68133), .I1(baudrate[11]), .I2(n27_adj_5131), 
            .I3(GND_net), .O(n68134));   // verilog/uart_rx.v(119[33:55])
    defparam i52406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51228_4_lut (.I0(n27_adj_5131), .I1(n25_adj_5127), .I2(n23_adj_5128), 
            .I3(n66065), .O(n66956));
    defparam i51228_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5141), .I1(baudrate[9]), 
            .I2(n23_adj_5128), .I3(GND_net), .O(n20_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46933_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[15]), .I1(baudrate[16]), 
            .I2(baudrate[17]), .I3(n25657), .O(n58469));
    defparam i46933_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i52298_3_lut (.I0(n68134), .I1(baudrate[12]), .I2(n29_adj_5130), 
            .I3(GND_net), .O(n26_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam i52298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52210_4_lut (.I0(n37_adj_5137), .I1(n35_adj_5138), .I2(n33_adj_5133), 
            .I3(n66055), .O(n67938));
    defparam i52210_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52850_4_lut (.I0(n68028), .I1(n68460), .I2(n39_adj_5135), 
            .I3(n66043), .O(n68578));   // verilog/uart_rx.v(119[33:55])
    defparam i52850_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51946_4_lut (.I0(n26_adj_5143), .I1(n20_adj_5142), .I2(n29_adj_5130), 
            .I3(n66956), .O(n67674));   // verilog/uart_rx.v(119[33:55])
    defparam i51946_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52876_4_lut (.I0(n67674), .I1(n68578), .I2(n39_adj_5135), 
            .I3(n67938), .O(n68604));   // verilog/uart_rx.v(119[33:55])
    defparam i52876_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52877_3_lut (.I0(n68604), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n68605));   // verilog/uart_rx.v(119[33:55])
    defparam i52877_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52867_3_lut (.I0(n68605), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n68595));   // verilog/uart_rx.v(119[33:55])
    defparam i52867_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51948_3_lut (.I0(n68595), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n67676));   // verilog/uart_rx.v(119[33:55])
    defparam i51948_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8373[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8399[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_986 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61094), .O(n61100));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_986.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_987 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61100), .O(n61106));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_987.LUT_INIT = 16'hfffe;
    SB_LUT4 i42751_1_lut_4_lut (.I0(n62276), .I1(n62278), .I2(n62114), 
            .I3(n62274), .O(n58437));
    defparam i42751_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29912));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i1_4_lut_adj_988 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61046), .O(n61052));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_988.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_989 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61052), .O(n61058));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 i47146_1_lut (.I0(n62864), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58487));
    defparam i47146_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50903_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4937), .I3(n57317), .O(n65654));
    defparam i50903_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i50900_4_lut (.I0(n65654), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65651));
    defparam i50900_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n65651), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27754));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i1_4_lut_adj_990 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61126), .O(n61132));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_991 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61132), .O(n61138));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_991.LUT_INIT = 16'hfffe;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29900));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50265_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n65993));
    defparam i50265_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n49674), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n60642), .I1(n25593), .I2(VCC_net), 
            .I3(n49673), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i50491_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n66219));
    defparam i50491_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY sub_38_add_2_25 (.CI(n49673), .I0(n25593), .I1(VCC_net), 
            .CO(n49674));
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n60742), .I1(n62906), .I2(VCC_net), 
            .I3(n49672), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50468_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n66196));
    defparam i50468_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY sub_38_add_2_24 (.CI(n49672), .I0(n62906), .I1(VCC_net), 
            .CO(n49673));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n49671), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_38_add_2_23 (.CI(n49671), .I0(n294[21]), .I1(VCC_net), 
            .CO(n49672));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n60740), .I1(n294[20]), .I2(VCC_net), 
            .I3(n49670), .O(n60742)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i47145_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n62840), .I3(baudrate[9]), .O(n62864));
    defparam i47145_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53676_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n62840), .I3(n48_adj_5151), .O(n294[14]));
    defparam i53676_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i53661_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n62870), .I3(n48_adj_5152), .O(n294[19]));
    defparam i53661_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8087[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8087[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8087[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8087[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8087[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8087[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_22 (.CI(n49670), .I0(n294[20]), .I1(VCC_net), 
            .CO(n49671));
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8087[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8087[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8087[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n62114));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_992 (.I0(n62158), .I1(n62114), .I2(n62116), .I3(baudrate[11]), 
            .O(n62144));
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_993 (.I0(n62144), .I1(n62146), .I2(n62134), .I3(n61998), 
            .O(n25636));
    defparam i1_4_lut_adj_993.LUT_INIT = 16'hfffe;
    SB_LUT4 i29014_rep_5_2_lut (.I0(n8087[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n58481));   // verilog/uart_rx.v(119[33:55])
    defparam i29014_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n58481), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52190_3_lut (.I0(n32_adj_5157), .I1(baudrate[6]), .I2(n39_adj_5155), 
            .I3(GND_net), .O(n67918));   // verilog/uart_rx.v(119[33:55])
    defparam i52190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52191_3_lut (.I0(n67918), .I1(baudrate[7]), .I2(n41_adj_5156), 
            .I3(GND_net), .O(n67919));   // verilog/uart_rx.v(119[33:55])
    defparam i52191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51592_4_lut (.I0(n41_adj_5156), .I1(n39_adj_5155), .I2(n37_adj_5154), 
            .I3(n66423), .O(n67320));
    defparam i51592_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n60738), .I1(n294[19]), .I2(VCC_net), 
            .I3(n49669), .O(n60740)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i52268_3_lut (.I0(n34_adj_5158), .I1(baudrate[5]), .I2(n37_adj_5154), 
            .I3(GND_net), .O(n67996));   // verilog/uart_rx.v(119[33:55])
    defparam i52268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47152_1_lut_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), 
            .I2(n62864), .I3(GND_net), .O(n58495));
    defparam i47152_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i51338_3_lut (.I0(n67919), .I1(baudrate[8]), .I2(n43_adj_5153), 
            .I3(GND_net), .O(n67066));   // verilog/uart_rx.v(119[33:55])
    defparam i51338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52491_4_lut (.I0(n67066), .I1(n67996), .I2(n43_adj_5153), 
            .I3(n67320), .O(n68219));   // verilog/uart_rx.v(119[33:55])
    defparam i52491_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_38_add_2_21 (.CI(n49669), .I0(n294[19]), .I1(VCC_net), 
            .CO(n49670));
    SB_LUT4 i52492_3_lut (.I0(n68219), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n68220));   // verilog/uart_rx.v(119[33:55])
    defparam i52492_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n68220), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5006));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n49668), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n49668), .I0(n294[18]), .I1(VCC_net), 
            .CO(n49669));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n60736), .I1(n294[17]), .I2(VCC_net), 
            .I3(n49667), .O(n60738)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29798));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29797));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29796));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n69846));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i50947_2_lut (.I0(n57075), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n65670));
    defparam i50947_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50944_4_lut (.I0(n65670), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n65667));
    defparam i50944_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50314_4_lut (.I0(n65667), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n65664));
    defparam i50314_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i53341_4_lut (.I0(\r_SM_Main[2] ), .I1(n65664), .I2(r_SM_Main_2__N_3446[1]), 
            .I3(\r_SM_Main[1] ), .O(n29178));
    defparam i53341_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_994 (.I0(n57075), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n60766));
    defparam i1_4_lut_adj_994.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_995 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n60766), .O(n60772));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'h0100;
    SB_LUT4 i52928_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n60772), .O(n27797));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52928_4_lut.LUT_INIT = 16'h5455;
    SB_CARRY sub_38_add_2_19 (.CI(n49667), .I0(n294[17]), .I1(VCC_net), 
            .CO(n49668));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n62030));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47087_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n62806));
    defparam i47087_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_38_add_2_18_lut (.I0(n60734), .I1(n294[16]), .I2(VCC_net), 
            .I3(n49666), .O(n60736)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_18 (.CI(n49666), .I0(n294[16]), .I1(VCC_net), 
            .CO(n49667));
    SB_LUT4 i1_2_lut_4_lut (.I0(n67676), .I1(baudrate[21]), .I2(n3046), 
            .I3(n60700), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n60640), .I1(n294[15]), .I2(VCC_net), 
            .I3(n49665), .O(n60642)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i47029_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n62748));
    defparam i47029_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53722_2_lut_4_lut (.I0(n67676), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25666), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i53722_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY sub_38_add_2_17 (.CI(n49665), .I0(n294[15]), .I1(VCC_net), 
            .CO(n49666));
    SB_LUT4 sub_38_add_2_16_lut (.I0(n60732), .I1(n294[14]), .I2(VCC_net), 
            .I3(n49664), .O(n60734)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[25]), .I2(baudrate[26]), 
            .I3(baudrate[29]), .O(n60660));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47033_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n62752));
    defparam i47033_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_996 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n61332));
    defparam i1_2_lut_4_lut_adj_996.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_997 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n62172));
    defparam i1_2_lut_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_LUT4 i50891_2_lut_3_lut (.I0(n25682), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n65705));   // verilog/uart_rx.v(119[33:55])
    defparam i50891_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_4_lut_adj_998 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n62174));
    defparam i1_2_lut_4_lut_adj_998.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_999 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n62134));
    defparam i1_2_lut_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 i50257_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5159), .I2(n25682), 
            .I3(GND_net), .O(n65985));   // verilog/uart_rx.v(119[33:55])
    defparam i50257_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_4_lut_adj_1000 (.I0(n68601), .I1(baudrate[20]), .I2(n2938), 
            .I3(n60698), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1000.LUT_INIT = 16'h7100;
    SB_CARRY sub_38_add_2_16 (.CI(n49664), .I0(n294[14]), .I1(VCC_net), 
            .CO(n49665));
    SB_LUT4 i2162_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2162_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2155_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2155_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1001 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n62010));
    defparam i1_2_lut_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1002 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n62012));
    defparam i1_2_lut_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 r_Clock_Count_1951_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n50920), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27996), 
            .D(n479[1]), .R(n58373));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27996), 
            .D(n479[2]), .R(n58373));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Clock_Count_1951__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27797), .D(n1[1]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27797), .D(n1[2]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27797), .D(n1[3]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27797), .D(n1[4]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27797), .D(n1[5]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27797), .D(n1[6]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27797), .D(n1[7]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27797), .D(n1[0]), .R(n29178));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 r_Clock_Count_1951_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n50919), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_8 (.CI(n50919), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n50920));
    SB_LUT4 r_Clock_Count_1951_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n50918), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_7 (.CI(n50918), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n50919));
    SB_LUT4 r_Clock_Count_1951_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n50917), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_6 (.CI(n50917), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n50918));
    SB_LUT4 r_Clock_Count_1951_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n50916), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_5 (.CI(n50916), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n50917));
    SB_LUT4 r_Clock_Count_1951_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n50915), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_4 (.CI(n50915), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n50916));
    SB_LUT4 r_Clock_Count_1951_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n50914), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_3 (.CI(n50914), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n50915));
    SB_LUT4 r_Clock_Count_1951_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n50914));
    SB_LUT4 i53717_2_lut_4_lut (.I0(n68601), .I1(baudrate[20]), .I2(n2938), 
            .I3(n62868), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i53717_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n49663), .O(n60732)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30533));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n53222));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30529));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2802_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n50760), 
            .O(n8425[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2802_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n50759), 
            .O(n8425[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_24 (.CI(n50759), .I0(n3152), .I1(n3082), .CO(n50760));
    SB_LUT4 add_2802_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n50758), 
            .O(n8425[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_23 (.CI(n50758), .I0(n3153), .I1(n3188), .CO(n50759));
    SB_LUT4 add_2802_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n50757), 
            .O(n8425[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_22 (.CI(n50757), .I0(n3154), .I1(n3084), .CO(n50758));
    SB_LUT4 add_2802_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n50756), 
            .O(n8425[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_21 (.CI(n50756), .I0(n3155), .I1(n2977), .CO(n50757));
    SB_LUT4 add_2802_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n50755), 
            .O(n8425[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_20 (.CI(n50755), .I0(n3156), .I1(n2867), .CO(n50756));
    SB_LUT4 add_2802_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n50754), 
            .O(n8425[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_19 (.CI(n50754), .I0(n3157), .I1(n2754), .CO(n50755));
    SB_LUT4 add_2802_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n50753), 
            .O(n8425[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_18 (.CI(n50753), .I0(n3158), .I1(n2638), .CO(n50754));
    SB_LUT4 add_2802_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n50752), 
            .O(n8425[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_17 (.CI(n50752), .I0(n3159), .I1(n2519), .CO(n50753));
    SB_LUT4 add_2802_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n50751), 
            .O(n8425[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_16 (.CI(n50751), .I0(n3160), .I1(n2397), .CO(n50752));
    SB_LUT4 add_2802_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n50750), 
            .O(n8425[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_15 (.CI(n50750), .I0(n3161), .I1(n2272), .CO(n50751));
    SB_LUT4 add_2802_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n50749), 
            .O(n8425[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_14 (.CI(n50749), .I0(n3162), .I1(n2144), .CO(n50750));
    SB_LUT4 add_2802_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n50748), 
            .O(n8425[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_13 (.CI(n50748), .I0(n3163), .I1(n2013), .CO(n50749));
    SB_LUT4 add_2802_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n50747), 
            .O(n8425[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_12 (.CI(n50747), .I0(n3164), .I1(n1879), .CO(n50748));
    SB_LUT4 add_2802_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n50746), 
            .O(n8425[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_11 (.CI(n50746), .I0(n3165), .I1(n1742), .CO(n50747));
    SB_LUT4 add_2802_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n50745), 
            .O(n8425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_10 (.CI(n50745), .I0(n3166), .I1(n1602), .CO(n50746));
    SB_LUT4 add_2802_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n50744), 
            .O(n8425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_9 (.CI(n50744), .I0(n3167), .I1(n1459), .CO(n50745));
    SB_LUT4 add_2802_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n50743), 
            .O(n8425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_8 (.CI(n50743), .I0(n3168), .I1(n1460), .CO(n50744));
    SB_LUT4 add_2802_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n50742), 
            .O(n8425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_7 (.CI(n50742), .I0(n3169), .I1(n1011), .CO(n50743));
    SB_LUT4 add_2802_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n50741), 
            .O(n8425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_6 (.CI(n50741), .I0(n3170), .I1(n856), .CO(n50742));
    SB_LUT4 add_2802_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n50740), 
            .O(n8425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_5 (.CI(n50740), .I0(n3171), .I1(n698), .CO(n50741));
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n30231));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n30230));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2802_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n50739), 
            .O(n8425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_4 (.CI(n50739), .I0(n3172), .I1(n858), .CO(n50740));
    SB_LUT4 add_2802_3_lut (.I0(n58437), .I1(GND_net), .I2(n538), .I3(n50738), 
            .O(n60702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2802_3 (.CI(n50738), .I0(GND_net), .I1(n538), .CO(n50739));
    SB_CARRY add_2802_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n50738));
    SB_LUT4 add_2801_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n50737), 
            .O(n8399[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2801_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n50736), 
            .O(n8399[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_22 (.CI(n50736), .I0(n3047), .I1(n3188), .CO(n50737));
    SB_LUT4 add_2801_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n50735), 
            .O(n8399[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_21 (.CI(n50735), .I0(n3048), .I1(n3084), .CO(n50736));
    SB_LUT4 add_2801_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n50734), 
            .O(n8399[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_20 (.CI(n50734), .I0(n3049), .I1(n2977), .CO(n50735));
    SB_LUT4 add_2801_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n50733), 
            .O(n8399[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_19 (.CI(n50733), .I0(n3050), .I1(n2867), .CO(n50734));
    SB_LUT4 add_2801_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n50732), 
            .O(n8399[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_18 (.CI(n50732), .I0(n3051), .I1(n2754), .CO(n50733));
    SB_LUT4 add_2801_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n50731), 
            .O(n8399[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_17 (.CI(n50731), .I0(n3052), .I1(n2638), .CO(n50732));
    SB_LUT4 add_2801_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n50730), 
            .O(n8399[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_16 (.CI(n50730), .I0(n3053), .I1(n2519), .CO(n50731));
    SB_LUT4 add_2801_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n50729), 
            .O(n8399[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_15 (.CI(n50729), .I0(n3054), .I1(n2397), .CO(n50730));
    SB_LUT4 add_2801_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n50728), 
            .O(n8399[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_14 (.CI(n50728), .I0(n3055), .I1(n2272), .CO(n50729));
    SB_LUT4 add_2801_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n50727), 
            .O(n8399[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_13 (.CI(n50727), .I0(n3056), .I1(n2144), .CO(n50728));
    SB_LUT4 add_2801_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n50726), 
            .O(n8399[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_12 (.CI(n50726), .I0(n3057), .I1(n2013), .CO(n50727));
    SB_LUT4 add_2801_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n50725), 
            .O(n8399[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_11 (.CI(n50725), .I0(n3058), .I1(n1879), .CO(n50726));
    SB_LUT4 add_2801_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n50724), 
            .O(n8399[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_10 (.CI(n50724), .I0(n3059), .I1(n1742), .CO(n50725));
    SB_LUT4 add_2801_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n50723), 
            .O(n8399[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_9 (.CI(n50723), .I0(n3060), .I1(n1602), .CO(n50724));
    SB_LUT4 add_2801_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n50722), 
            .O(n8399[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_8 (.CI(n50722), .I0(n3061), .I1(n1459), .CO(n50723));
    SB_LUT4 add_2801_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n50721), 
            .O(n8399[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_7 (.CI(n50721), .I0(n3062), .I1(n1460), .CO(n50722));
    SB_LUT4 add_2801_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n50720), 
            .O(n8399[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_6 (.CI(n50720), .I0(n3063), .I1(n1011), .CO(n50721));
    SB_LUT4 add_2801_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n50719), 
            .O(n8399[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_5 (.CI(n50719), .I0(n3064), .I1(n856), .CO(n50720));
    SB_LUT4 add_2801_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n50718), 
            .O(n8399[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_4 (.CI(n50718), .I0(n3065), .I1(n698), .CO(n50719));
    SB_LUT4 add_2801_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n50717), 
            .O(n8399[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_3 (.CI(n50717), .I0(n3066), .I1(n858), .CO(n50718));
    SB_LUT4 add_2801_2_lut (.I0(n58441), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2801_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50717));
    SB_LUT4 add_2800_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n50716), 
            .O(n8373[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2800_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n50715), 
            .O(n8373[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_21 (.CI(n50715), .I0(n2939), .I1(n3084), .CO(n50716));
    SB_LUT4 add_2800_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n50714), 
            .O(n8373[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_20 (.CI(n50714), .I0(n2940), .I1(n2977), .CO(n50715));
    SB_LUT4 add_2800_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n50713), 
            .O(n8373[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_19 (.CI(n50713), .I0(n2941), .I1(n2867), .CO(n50714));
    SB_LUT4 add_2800_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n50712), 
            .O(n8373[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_18 (.CI(n50712), .I0(n2942), .I1(n2754), .CO(n50713));
    SB_LUT4 add_2800_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n50711), 
            .O(n8373[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_17 (.CI(n50711), .I0(n2943), .I1(n2638), .CO(n50712));
    SB_LUT4 add_2800_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n50710), 
            .O(n8373[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_16 (.CI(n50710), .I0(n2944), .I1(n2519), .CO(n50711));
    SB_LUT4 add_2800_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n50709), 
            .O(n8373[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_15 (.CI(n50709), .I0(n2945), .I1(n2397), .CO(n50710));
    SB_LUT4 add_2800_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n50708), 
            .O(n8373[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_14 (.CI(n50708), .I0(n2946), .I1(n2272), .CO(n50709));
    SB_CARRY sub_38_add_2_15 (.CI(n49663), .I0(n294[13]), .I1(VCC_net), 
            .CO(n49664));
    SB_LUT4 add_2800_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n50707), 
            .O(n8373[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_13 (.CI(n50707), .I0(n2947), .I1(n2144), .CO(n50708));
    SB_LUT4 add_2800_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n50706), 
            .O(n8373[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_12 (.CI(n50706), .I0(n2948), .I1(n2013), .CO(n50707));
    SB_LUT4 add_2800_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n50705), 
            .O(n8373[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_11 (.CI(n50705), .I0(n2949), .I1(n1879), .CO(n50706));
    SB_LUT4 add_2800_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n50704), 
            .O(n8373[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_10 (.CI(n50704), .I0(n2950), .I1(n1742), .CO(n50705));
    SB_LUT4 add_2800_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n50703), 
            .O(n8373[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_9 (.CI(n50703), .I0(n2951), .I1(n1602), .CO(n50704));
    SB_LUT4 add_2800_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n50702), 
            .O(n8373[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_8 (.CI(n50702), .I0(n2952), .I1(n1459), .CO(n50703));
    SB_LUT4 add_2800_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n50701), 
            .O(n8373[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_7 (.CI(n50701), .I0(n2953), .I1(n1460), .CO(n50702));
    SB_LUT4 add_2800_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n50700), 
            .O(n8373[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_6 (.CI(n50700), .I0(n2954), .I1(n1011), .CO(n50701));
    SB_LUT4 add_2800_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n50699), 
            .O(n8373[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_5 (.CI(n50699), .I0(n2955), .I1(n856), .CO(n50700));
    SB_LUT4 add_2800_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n50698), 
            .O(n8373[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_4 (.CI(n50698), .I0(n2956), .I1(n698), .CO(n50699));
    SB_LUT4 add_2800_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n50697), 
            .O(n8373[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_3 (.CI(n50697), .I0(n2957), .I1(n858), .CO(n50698));
    SB_LUT4 add_2800_2_lut (.I0(n58445), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2800_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50697));
    SB_LUT4 add_2799_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n50696), 
            .O(n8347[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n50695), 
            .O(n8347[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_20 (.CI(n50695), .I0(n2828), .I1(n2977), .CO(n50696));
    SB_LUT4 add_2799_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n50694), 
            .O(n8347[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_19 (.CI(n50694), .I0(n2829), .I1(n2867), .CO(n50695));
    SB_LUT4 add_2799_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n50693), 
            .O(n8347[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_18 (.CI(n50693), .I0(n2830), .I1(n2754), .CO(n50694));
    SB_LUT4 add_2799_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n50692), 
            .O(n8347[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_17 (.CI(n50692), .I0(n2831), .I1(n2638), .CO(n50693));
    SB_LUT4 add_2799_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n50691), 
            .O(n8347[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_16 (.CI(n50691), .I0(n2832), .I1(n2519), .CO(n50692));
    SB_LUT4 add_2799_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n50690), 
            .O(n8347[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_15 (.CI(n50690), .I0(n2833), .I1(n2397), .CO(n50691));
    SB_LUT4 add_2799_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n50689), 
            .O(n8347[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_14 (.CI(n50689), .I0(n2834), .I1(n2272), .CO(n50690));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n49662), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2799_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n50688), 
            .O(n8347[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_13 (.CI(n50688), .I0(n2835), .I1(n2144), .CO(n50689));
    SB_LUT4 add_2799_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n50687), 
            .O(n8347[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_12 (.CI(n50687), .I0(n2836), .I1(n2013), .CO(n50688));
    SB_LUT4 add_2799_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n50686), 
            .O(n8347[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_11 (.CI(n50686), .I0(n2837), .I1(n1879), .CO(n50687));
    SB_CARRY sub_38_add_2_14 (.CI(n49662), .I0(n294[12]), .I1(VCC_net), 
            .CO(n49663));
    SB_LUT4 add_2799_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n50685), 
            .O(n8347[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_10 (.CI(n50685), .I0(n2838), .I1(n1742), .CO(n50686));
    SB_LUT4 add_2799_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n50684), 
            .O(n8347[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_9 (.CI(n50684), .I0(n2839), .I1(n1602), .CO(n50685));
    SB_LUT4 add_2799_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n50683), 
            .O(n8347[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_8 (.CI(n50683), .I0(n2840), .I1(n1459), .CO(n50684));
    SB_LUT4 add_2799_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n50682), 
            .O(n8347[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_7 (.CI(n50682), .I0(n2841), .I1(n1460), .CO(n50683));
    SB_LUT4 add_2799_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n50681), 
            .O(n8347[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_6 (.CI(n50681), .I0(n2842), .I1(n1011), .CO(n50682));
    SB_LUT4 add_2799_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n50680), 
            .O(n8347[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_5 (.CI(n50680), .I0(n2843), .I1(n856), .CO(n50681));
    SB_LUT4 add_2799_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n50679), 
            .O(n8347[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_4 (.CI(n50679), .I0(n2844), .I1(n698), .CO(n50680));
    SB_LUT4 add_2799_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n50678), 
            .O(n8347[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_3 (.CI(n50678), .I0(n2845), .I1(n858), .CO(n50679));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n49661), .O(n60640)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2799_2_lut (.I0(n58449), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2799_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50678));
    SB_LUT4 add_2798_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n50677), 
            .O(n8321[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2798_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n50676), 
            .O(n8321[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_19 (.CI(n50676), .I0(n2714), .I1(n2867), .CO(n50677));
    SB_LUT4 add_2798_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n50675), 
            .O(n8321[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_18 (.CI(n50675), .I0(n2715), .I1(n2754), .CO(n50676));
    SB_LUT4 add_2798_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n50674), 
            .O(n8321[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_17 (.CI(n50674), .I0(n2716), .I1(n2638), .CO(n50675));
    SB_LUT4 add_2798_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n50673), 
            .O(n8321[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_16 (.CI(n50673), .I0(n2717), .I1(n2519), .CO(n50674));
    SB_LUT4 add_2798_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n50672), 
            .O(n8321[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_15 (.CI(n50672), .I0(n2718), .I1(n2397), .CO(n50673));
    SB_LUT4 add_2798_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n50671), 
            .O(n8321[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_14 (.CI(n50671), .I0(n2719), .I1(n2272), .CO(n50672));
    SB_LUT4 add_2798_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n50670), 
            .O(n8321[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_13 (.CI(n50670), .I0(n2720), .I1(n2144), .CO(n50671));
    SB_LUT4 add_2798_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n50669), 
            .O(n8321[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_12 (.CI(n50669), .I0(n2721), .I1(n2013), .CO(n50670));
    SB_LUT4 add_2798_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n50668), 
            .O(n8321[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_11 (.CI(n50668), .I0(n2722), .I1(n1879), .CO(n50669));
    SB_LUT4 add_2798_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n50667), 
            .O(n8321[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_10 (.CI(n50667), .I0(n2723), .I1(n1742), .CO(n50668));
    SB_LUT4 add_2798_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n50666), 
            .O(n8321[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_9 (.CI(n50666), .I0(n2724), .I1(n1602), .CO(n50667));
    SB_LUT4 add_2798_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n50665), 
            .O(n8321[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_8 (.CI(n50665), .I0(n2725), .I1(n1459), .CO(n50666));
    SB_LUT4 add_2798_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n50664), 
            .O(n8321[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_7 (.CI(n50664), .I0(n2726), .I1(n1460), .CO(n50665));
    SB_LUT4 add_2798_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n50663), 
            .O(n8321[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_6 (.CI(n50663), .I0(n2727), .I1(n1011), .CO(n50664));
    SB_LUT4 add_2798_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n50662), 
            .O(n8321[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_5 (.CI(n50662), .I0(n2728), .I1(n856), .CO(n50663));
    SB_LUT4 add_2798_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n50661), 
            .O(n8321[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_4 (.CI(n50661), .I0(n2729), .I1(n698), .CO(n50662));
    SB_LUT4 add_2798_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n50660), 
            .O(n8321[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_3 (.CI(n50660), .I0(n2730), .I1(n858), .CO(n50661));
    SB_LUT4 add_2798_2_lut (.I0(n58453), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2798_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50660));
    SB_LUT4 add_2797_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n50659), 
            .O(n8295[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n50658), 
            .O(n8295[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_18 (.CI(n50658), .I0(n2597), .I1(n2754), .CO(n50659));
    SB_LUT4 add_2797_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n50657), 
            .O(n8295[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_17 (.CI(n50657), .I0(n2598), .I1(n2638), .CO(n50658));
    SB_LUT4 add_2797_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n50656), 
            .O(n8295[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_16 (.CI(n50656), .I0(n2599), .I1(n2519), .CO(n50657));
    SB_LUT4 add_2797_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n50655), 
            .O(n8295[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_15 (.CI(n50655), .I0(n2600), .I1(n2397), .CO(n50656));
    SB_LUT4 add_2797_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n50654), 
            .O(n8295[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_14 (.CI(n50654), .I0(n2601), .I1(n2272), .CO(n50655));
    SB_LUT4 add_2797_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n50653), 
            .O(n8295[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_13 (.CI(n49661), .I0(n294[11]), .I1(VCC_net), 
            .CO(n49662));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n49660), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_13 (.CI(n50653), .I0(n2602), .I1(n2144), .CO(n50654));
    SB_CARRY sub_38_add_2_12 (.CI(n49660), .I0(n294[10]), .I1(VCC_net), 
            .CO(n49661));
    SB_LUT4 add_2797_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n50652), 
            .O(n8295[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_12 (.CI(n50652), .I0(n2603), .I1(n2013), .CO(n50653));
    SB_LUT4 add_2797_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n50651), 
            .O(n8295[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_11 (.CI(n50651), .I0(n2604), .I1(n1879), .CO(n50652));
    SB_LUT4 add_2797_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n50650), 
            .O(n8295[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_10 (.CI(n50650), .I0(n2605), .I1(n1742), .CO(n50651));
    SB_LUT4 add_2797_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n50649), 
            .O(n8295[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1003 (.I0(n68587), .I1(baudrate[19]), .I2(n2827), 
            .I3(n60696), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1003.LUT_INIT = 16'h7100;
    SB_CARRY add_2797_9 (.CI(n50649), .I0(n2606), .I1(n1602), .CO(n50650));
    SB_LUT4 add_2797_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n50648), 
            .O(n8295[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_8 (.CI(n50648), .I0(n2607), .I1(n1459), .CO(n50649));
    SB_LUT4 add_2797_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n50647), 
            .O(n8295[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_7 (.CI(n50647), .I0(n2608), .I1(n1460), .CO(n50648));
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_5166), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2797_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n50646), 
            .O(n8295[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_6 (.CI(n50646), .I0(n2609), .I1(n1011), .CO(n50647));
    SB_LUT4 add_2797_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n50645), 
            .O(n8295[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_5 (.CI(n50645), .I0(n2610), .I1(n856), .CO(n50646));
    SB_LUT4 add_2797_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n50644), 
            .O(n8295[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_4 (.CI(n50644), .I0(n2611), .I1(n698), .CO(n50645));
    SB_LUT4 add_2797_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n50643), 
            .O(n8295[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_3 (.CI(n50643), .I0(n2612), .I1(n858), .CO(n50644));
    SB_LUT4 add_2797_2_lut (.I0(n58457), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2797_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50643));
    SB_LUT4 add_2796_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n50642), 
            .O(n8269[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2796_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n50641), 
            .O(n8269[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_17 (.CI(n50641), .I0(n2477), .I1(n2638), .CO(n50642));
    SB_LUT4 add_2796_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n50640), 
            .O(n8269[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_16 (.CI(n50640), .I0(n2478), .I1(n2519), .CO(n50641));
    SB_LUT4 add_2796_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n50639), 
            .O(n8269[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_15 (.CI(n50639), .I0(n2479), .I1(n2397), .CO(n50640));
    SB_LUT4 add_2796_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n50638), 
            .O(n8269[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_14 (.CI(n50638), .I0(n2480), .I1(n2272), .CO(n50639));
    SB_LUT4 add_2796_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n50637), 
            .O(n8269[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_13 (.CI(n50637), .I0(n2481), .I1(n2144), .CO(n50638));
    SB_LUT4 add_2796_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n50636), 
            .O(n8269[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_12 (.CI(n50636), .I0(n2482), .I1(n2013), .CO(n50637));
    SB_LUT4 add_2796_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n50635), 
            .O(n8269[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_11 (.CI(n50635), .I0(n2483), .I1(n1879), .CO(n50636));
    SB_LUT4 add_2796_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n50634), 
            .O(n8269[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_10 (.CI(n50634), .I0(n2484), .I1(n1742), .CO(n50635));
    SB_LUT4 add_2796_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n50633), 
            .O(n8269[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_9 (.CI(n50633), .I0(n2485), .I1(n1602), .CO(n50634));
    SB_LUT4 add_2796_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n50632), 
            .O(n8269[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_8 (.CI(n50632), .I0(n2486), .I1(n1459), .CO(n50633));
    SB_LUT4 add_2796_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n50631), 
            .O(n8269[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_7 (.CI(n50631), .I0(n2487), .I1(n1460), .CO(n50632));
    SB_LUT4 add_2796_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n50630), 
            .O(n8269[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_6 (.CI(n50630), .I0(n2488), .I1(n1011), .CO(n50631));
    SB_LUT4 add_2796_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n50629), 
            .O(n8269[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_5 (.CI(n50629), .I0(n2489), .I1(n856), .CO(n50630));
    SB_LUT4 add_2796_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n50628), 
            .O(n8269[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_4 (.CI(n50628), .I0(n2490), .I1(n698), .CO(n50629));
    SB_LUT4 add_2796_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n50627), 
            .O(n8269[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_3 (.CI(n50627), .I0(n2491), .I1(n858), .CO(n50628));
    SB_LUT4 add_2796_2_lut (.I0(n58461), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2796_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50627));
    SB_LUT4 add_2795_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n50626), 
            .O(n8243[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n50625), 
            .O(n8243[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_16 (.CI(n50625), .I0(n2354), .I1(n2519), .CO(n50626));
    SB_LUT4 add_2795_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n50624), 
            .O(n8243[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_15 (.CI(n50624), .I0(n2355), .I1(n2397), .CO(n50625));
    SB_LUT4 add_2795_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n50623), 
            .O(n8243[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_14 (.CI(n50623), .I0(n2356), .I1(n2272), .CO(n50624));
    SB_LUT4 add_2795_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n50622), 
            .O(n8243[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_13 (.CI(n50622), .I0(n2357), .I1(n2144), .CO(n50623));
    SB_LUT4 add_2795_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n50621), 
            .O(n8243[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_12 (.CI(n50621), .I0(n2358), .I1(n2013), .CO(n50622));
    SB_LUT4 add_2795_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n50620), 
            .O(n8243[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_11 (.CI(n50620), .I0(n2359), .I1(n1879), .CO(n50621));
    SB_LUT4 add_2795_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n50619), 
            .O(n8243[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_10 (.CI(n50619), .I0(n2360), .I1(n1742), .CO(n50620));
    SB_LUT4 add_2795_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n50618), 
            .O(n8243[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_9 (.CI(n50618), .I0(n2361), .I1(n1602), .CO(n50619));
    SB_LUT4 add_2795_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n50617), 
            .O(n8243[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_8 (.CI(n50617), .I0(n2362), .I1(n1459), .CO(n50618));
    SB_LUT4 add_2795_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n50616), 
            .O(n8243[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_7 (.CI(n50616), .I0(n2363), .I1(n1460), .CO(n50617));
    SB_LUT4 add_2795_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n50615), 
            .O(n8243[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_6 (.CI(n50615), .I0(n2364), .I1(n1011), .CO(n50616));
    SB_LUT4 add_2795_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n50614), 
            .O(n8243[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_5 (.CI(n50614), .I0(n2365), .I1(n856), .CO(n50615));
    SB_LUT4 add_2795_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n50613), 
            .O(n8243[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_4 (.CI(n50613), .I0(n2366), .I1(n698), .CO(n50614));
    SB_LUT4 add_2795_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n50612), 
            .O(n8243[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_3 (.CI(n50612), .I0(n2367), .I1(n858), .CO(n50613));
    SB_LUT4 add_2795_2_lut (.I0(n58465), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2795_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50612));
    SB_LUT4 add_2794_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n50611), 
            .O(n8217[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n50610), 
            .O(n8217[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_15 (.CI(n50610), .I0(n2228), .I1(n2397), .CO(n50611));
    SB_LUT4 add_2794_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n50609), 
            .O(n8217[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_14 (.CI(n50609), .I0(n2229), .I1(n2272), .CO(n50610));
    SB_LUT4 add_2794_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n50608), 
            .O(n8217[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_13 (.CI(n50608), .I0(n2230), .I1(n2144), .CO(n50609));
    SB_LUT4 add_2794_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n50607), 
            .O(n8217[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_12 (.CI(n50607), .I0(n2231), .I1(n2013), .CO(n50608));
    SB_LUT4 add_2794_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n50606), 
            .O(n8217[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_11 (.CI(n50606), .I0(n2232), .I1(n1879), .CO(n50607));
    SB_LUT4 add_2794_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n50605), 
            .O(n8217[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_10 (.CI(n50605), .I0(n2233), .I1(n1742), .CO(n50606));
    SB_LUT4 add_2794_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n50604), 
            .O(n8217[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_9 (.CI(n50604), .I0(n2234), .I1(n1602), .CO(n50605));
    SB_LUT4 add_2794_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n50603), 
            .O(n8217[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_8 (.CI(n50603), .I0(n2235), .I1(n1459), .CO(n50604));
    SB_LUT4 add_2794_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n50602), 
            .O(n8217[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_7 (.CI(n50602), .I0(n2236), .I1(n1460), .CO(n50603));
    SB_LUT4 add_2794_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n50601), 
            .O(n8217[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_6 (.CI(n50601), .I0(n2237), .I1(n1011), .CO(n50602));
    SB_LUT4 add_2794_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n50600), 
            .O(n8217[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_5 (.CI(n50600), .I0(n2238), .I1(n856), .CO(n50601));
    SB_LUT4 add_2794_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n50599), 
            .O(n8217[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_4 (.CI(n50599), .I0(n2239), .I1(n698), .CO(n50600));
    SB_LUT4 add_2794_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n50598), 
            .O(n8217[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_3 (.CI(n50598), .I0(n2240), .I1(n858), .CO(n50599));
    SB_LUT4 add_2794_2_lut (.I0(n58469), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2794_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50598));
    SB_LUT4 add_2793_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n50597), 
            .O(n8191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n50596), 
            .O(n8191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_13 (.CI(n50596), .I0(n2099), .I1(n2272), .CO(n50597));
    SB_LUT4 add_2793_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n50595), 
            .O(n8191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_12 (.CI(n50595), .I0(n2100), .I1(n2144), .CO(n50596));
    SB_LUT4 add_2793_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n50594), 
            .O(n8191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_11 (.CI(n50594), .I0(n2101), .I1(n2013), .CO(n50595));
    SB_LUT4 add_2793_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n50593), 
            .O(n8191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_10 (.CI(n50593), .I0(n2102), .I1(n1879), .CO(n50594));
    SB_LUT4 add_2793_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n50592), 
            .O(n8191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_9 (.CI(n50592), .I0(n2103), .I1(n1742), .CO(n50593));
    SB_LUT4 add_2793_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n50591), 
            .O(n8191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_8 (.CI(n50591), .I0(n2104), .I1(n1602), .CO(n50592));
    SB_LUT4 add_2793_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n50590), 
            .O(n8191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_7 (.CI(n50590), .I0(n2105), .I1(n1459), .CO(n50591));
    SB_LUT4 add_2793_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n50589), 
            .O(n8191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_6 (.CI(n50589), .I0(n2106), .I1(n1460), .CO(n50590));
    SB_LUT4 add_2793_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n50588), 
            .O(n8191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_5 (.CI(n50588), .I0(n2107), .I1(n1011), .CO(n50589));
    SB_LUT4 add_2793_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n50587), 
            .O(n8191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_4 (.CI(n50587), .I0(n2108), .I1(n856), .CO(n50588));
    SB_LUT4 add_2793_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n50586), 
            .O(n8191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_3 (.CI(n50586), .I0(n2109), .I1(n698), .CO(n50587));
    SB_LUT4 add_2793_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n50586));
    SB_LUT4 add_2792_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n50585), 
            .O(n8165[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n50584), 
            .O(n8165[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_13 (.CI(n50584), .I0(n1967), .I1(n2144), .CO(n50585));
    SB_LUT4 add_2792_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n50583), 
            .O(n8165[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_12 (.CI(n50583), .I0(n1968), .I1(n2013), .CO(n50584));
    SB_LUT4 add_2792_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n50582), 
            .O(n8165[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_11 (.CI(n50582), .I0(n1969), .I1(n1879), .CO(n50583));
    SB_LUT4 add_2792_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n50581), 
            .O(n8165[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_10 (.CI(n50581), .I0(n1970), .I1(n1742), .CO(n50582));
    SB_LUT4 add_2792_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n50580), 
            .O(n8165[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_9 (.CI(n50580), .I0(n1971), .I1(n1602), .CO(n50581));
    SB_LUT4 add_2792_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n50579), 
            .O(n8165[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_8 (.CI(n50579), .I0(n1972), .I1(n1459), .CO(n50580));
    SB_LUT4 add_2792_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n50578), 
            .O(n8165[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_7 (.CI(n50578), .I0(n1973), .I1(n1460), .CO(n50579));
    SB_LUT4 add_2792_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n50577), 
            .O(n8165[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_6 (.CI(n50577), .I0(n1974), .I1(n1011), .CO(n50578));
    SB_LUT4 add_2792_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n50576), 
            .O(n8165[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_5 (.CI(n50576), .I0(n1975), .I1(n856), .CO(n50577));
    SB_LUT4 add_2792_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n50575), 
            .O(n8165[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_4 (.CI(n50575), .I0(n1976), .I1(n698), .CO(n50576));
    SB_LUT4 add_2792_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n50574), 
            .O(n8165[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_3 (.CI(n50574), .I0(n1977), .I1(n858), .CO(n50575));
    SB_LUT4 add_2792_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8165[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50574));
    SB_LUT4 add_2791_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n50573), 
            .O(n8139[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n50572), 
            .O(n8139[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_12 (.CI(n50572), .I0(n1832), .I1(n2013), .CO(n50573));
    SB_LUT4 add_2791_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n50571), 
            .O(n8139[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_11 (.CI(n50571), .I0(n1833), .I1(n1879), .CO(n50572));
    SB_LUT4 add_2791_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n50570), 
            .O(n8139[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_10 (.CI(n50570), .I0(n1834), .I1(n1742), .CO(n50571));
    SB_LUT4 add_2791_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n50569), 
            .O(n8139[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_9 (.CI(n50569), .I0(n1835), .I1(n1602), .CO(n50570));
    SB_LUT4 add_2791_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n50568), 
            .O(n8139[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_8 (.CI(n50568), .I0(n1836), .I1(n1459), .CO(n50569));
    SB_LUT4 add_2791_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n50567), 
            .O(n8139[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_7 (.CI(n50567), .I0(n1837), .I1(n1460), .CO(n50568));
    SB_LUT4 add_2791_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n50566), 
            .O(n8139[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_6 (.CI(n50566), .I0(n1838), .I1(n1011), .CO(n50567));
    SB_LUT4 add_2791_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n50565), 
            .O(n8139[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_5 (.CI(n50565), .I0(n1839), .I1(n856), .CO(n50566));
    SB_LUT4 add_2791_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n50564), 
            .O(n8139[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_4 (.CI(n50564), .I0(n1840), .I1(n698), .CO(n50565));
    SB_LUT4 add_2791_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n50563), 
            .O(n8139[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_3 (.CI(n50563), .I0(n1841), .I1(n858), .CO(n50564));
    SB_LUT4 add_2791_2_lut (.I0(n58478), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2791_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50563));
    SB_LUT4 add_2790_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n50562), 
            .O(n8113[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n50561), 
            .O(n8113[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_10 (.CI(n50561), .I0(n1694), .I1(n1879), .CO(n50562));
    SB_LUT4 add_2790_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n50560), 
            .O(n8113[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_9 (.CI(n50560), .I0(n1695), .I1(n1742), .CO(n50561));
    SB_LUT4 add_2790_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n50559), 
            .O(n8113[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_8 (.CI(n50559), .I0(n1696), .I1(n1602), .CO(n50560));
    SB_LUT4 add_2790_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n50558), 
            .O(n8113[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_7 (.CI(n50558), .I0(n1697), .I1(n1459), .CO(n50559));
    SB_LUT4 add_2790_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n50557), 
            .O(n8113[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_6 (.CI(n50557), .I0(n1698), .I1(n1460), .CO(n50558));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n49659), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n50556), 
            .O(n8113[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_5 (.CI(n50556), .I0(n1699), .I1(n1011), .CO(n50557));
    SB_LUT4 add_2790_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n50555), 
            .O(n8113[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_4 (.CI(n50555), .I0(n1700), .I1(n856), .CO(n50556));
    SB_LUT4 add_2790_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n50554), 
            .O(n8113[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_3 (.CI(n50554), .I0(n1701), .I1(n698), .CO(n50555));
    SB_LUT4 add_2790_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8113[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n50554));
    SB_LUT4 add_2789_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n50553), 
            .O(n8087[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2789_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n50552), 
            .O(n8087[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_10 (.CI(n50552), .I0(n1553), .I1(n1742), .CO(n50553));
    SB_LUT4 add_2789_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n50551), 
            .O(n8087[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_9 (.CI(n50551), .I0(n1554), .I1(n1602), .CO(n50552));
    SB_LUT4 add_2789_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n50550), 
            .O(n8087[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_8 (.CI(n50550), .I0(n1555), .I1(n1459), .CO(n50551));
    SB_LUT4 add_2789_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n50549), 
            .O(n8087[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_7 (.CI(n50549), .I0(n1556), .I1(n1460), .CO(n50550));
    SB_LUT4 add_2789_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n50548), 
            .O(n8087[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_6 (.CI(n50548), .I0(n1557), .I1(n1011), .CO(n50549));
    SB_LUT4 add_2789_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n50547), 
            .O(n8087[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_5 (.CI(n50547), .I0(n1558), .I1(n856), .CO(n50548));
    SB_LUT4 add_2789_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n50546), 
            .O(n8087[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_4 (.CI(n50546), .I0(n1559), .I1(n698), .CO(n50547));
    SB_LUT4 add_2789_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n50545), 
            .O(n8087[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53714_2_lut_4_lut (.I0(n68587), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25663), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i53714_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY add_2789_3 (.CI(n50545), .I0(n1560), .I1(n858), .CO(n50546));
    SB_LUT4 i53695_2_lut_4_lut (.I0(n68479), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25657), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i53695_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 add_2789_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8087[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50545));
    SB_LUT4 add_2788_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n50544), 
            .O(n8061[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2788_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n50543), 
            .O(n8061[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_9 (.CI(n50543), .I0(n1409), .I1(n1602), .CO(n50544));
    SB_LUT4 add_2788_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n50542), 
            .O(n8061[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_8 (.CI(n50542), .I0(n1410), .I1(n1459), .CO(n50543));
    SB_LUT4 add_2788_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n50541), 
            .O(n8061[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_7 (.CI(n50541), .I0(n1411), .I1(n1460), .CO(n50542));
    SB_LUT4 add_2788_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n50540), 
            .O(n8061[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_6 (.CI(n50540), .I0(n1412), .I1(n1011), .CO(n50541));
    SB_LUT4 add_2788_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n50539), 
            .O(n8061[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_5 (.CI(n50539), .I0(n1413), .I1(n856), .CO(n50540));
    SB_LUT4 add_2788_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n50538), 
            .O(n8061[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_4 (.CI(n50538), .I0(n1414), .I1(n698), .CO(n50539));
    SB_LUT4 add_2788_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n50537), 
            .O(n8061[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_3 (.CI(n50537), .I0(n1415), .I1(n858), .CO(n50538));
    SB_LUT4 add_2788_2_lut (.I0(n58487), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2788_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50537));
    SB_LUT4 add_2787_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n50536), 
            .O(n8035[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2787_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n50535), 
            .O(n8035[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1004 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4940), 
            .I3(\r_SM_Main[0] ), .O(n60748));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'hfeff;
    SB_CARRY add_2787_8 (.CI(n50535), .I0(n1262), .I1(n1459), .CO(n50536));
    SB_LUT4 i1_4_lut_adj_1005 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n60748), .O(n58925));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1005.LUT_INIT = 16'hfffe;
    SB_CARRY sub_38_add_2_11 (.CI(n49659), .I0(n294[9]), .I1(VCC_net), 
            .CO(n49660));
    SB_LUT4 i1_2_lut_4_lut_adj_1006 (.I0(n68479), .I1(baudrate[17]), .I2(n2596), 
            .I3(n60692), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1006.LUT_INIT = 16'h7100;
    SB_LUT4 add_2787_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n50534), 
            .O(n8035[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_7 (.CI(n50534), .I0(n1263), .I1(n1460), .CO(n50535));
    SB_LUT4 add_2787_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n50533), 
            .O(n8035[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_6 (.CI(n50533), .I0(n1264), .I1(n1011), .CO(n50534));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n49658), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2787_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n50532), 
            .O(n8035[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_5 (.CI(n50532), .I0(n1265), .I1(n856), .CO(n50533));
    SB_LUT4 add_2787_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n50531), 
            .O(n8035[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_4 (.CI(n50531), .I0(n1266), .I1(n698), .CO(n50532));
    SB_LUT4 add_2787_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n50530), 
            .O(n8035[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_3 (.CI(n50530), .I0(n1267), .I1(n858), .CO(n50531));
    SB_LUT4 add_2787_2_lut (.I0(n58491), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2787_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50530));
    SB_LUT4 add_2786_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n50529), 
            .O(n8009[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2786_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n50528), 
            .O(n8009[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_7 (.CI(n50528), .I0(n1112), .I1(n1460), .CO(n50529));
    SB_LUT4 add_2786_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n50527), 
            .O(n8009[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_6 (.CI(n50527), .I0(n1113), .I1(n1011), .CO(n50528));
    SB_LUT4 add_2786_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n50526), 
            .O(n8009[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_5 (.CI(n50526), .I0(n1114), .I1(n856), .CO(n50527));
    SB_CARRY sub_38_add_2_10 (.CI(n49658), .I0(n294[8]), .I1(VCC_net), 
            .CO(n49659));
    SB_LUT4 add_2786_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n50525), 
            .O(n8009[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_4 (.CI(n50525), .I0(n1115), .I1(n698), .CO(n50526));
    SB_LUT4 add_2786_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n50524), 
            .O(n8009[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_3 (.CI(n50524), .I0(n1116), .I1(n858), .CO(n50525));
    SB_LUT4 add_2786_2_lut (.I0(n58495), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2786_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50524));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n49657), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n49657), .I0(n294[7]), .I1(VCC_net), 
            .CO(n49658));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n49656), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n49656), .I0(n294[6]), .I1(VCC_net), 
            .CO(n49657));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n49655), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n49655), .I0(n294[5]), .I1(VCC_net), 
            .CO(n49656));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n49654), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n49654), .I0(n294[4]), .I1(VCC_net), 
            .CO(n49655));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n49653), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n49653), .I0(n294[3]), .I1(VCC_net), 
            .CO(n49654));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n49652), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n49652), .I0(n294[2]), .I1(VCC_net), 
            .CO(n49653));
    SB_LUT4 i47151_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), .I2(n62864), 
            .I3(GND_net), .O(n62870));
    defparam i47151_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n49651), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n49651), .I0(n294[1]), .I1(VCC_net), 
            .CO(n49652));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n59626), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n59626), .I1(GND_net), 
            .CO(n49651));
    SB_LUT4 i46930_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), .I2(n25657), 
            .I3(GND_net), .O(n62648));
    defparam i46930_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i53541_4_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(n6), .I3(n60115), .O(n58373));
    defparam i53541_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i50259_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5168), .I2(n25692), 
            .I3(GND_net), .O(n65987));   // verilog/uart_rx.v(119[33:55])
    defparam i50259_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_1007 (.I0(n25682), .I1(n48_adj_5159), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5169));
    defparam i1_3_lut_4_lut_adj_1007.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_4_lut_adj_1008 (.I0(n68008), .I1(baudrate[16]), .I2(n2476), 
            .I3(n60690), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1008.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n62278));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i53692_2_lut_4_lut (.I0(n68008), .I1(baudrate[16]), .I2(n2476), 
            .I3(n62602), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i53692_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i47122_1_lut (.I0(n62840), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58478));
    defparam i47122_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5578_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam i5578_2_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i7242_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n20994));   // verilog/uart_rx.v(119[33:55])
    defparam i7242_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8061[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8061[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8061[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8061[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8061[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8061[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8061[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8061[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50896_3_lut_4_lut (.I0(n962), .I1(baudrate[1]), .I2(n48_adj_5175), 
            .I3(n25605), .O(n1115));
    defparam i50896_3_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i5749_2_lut_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), 
            .I3(baudrate[1]), .O(n42_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam i5749_2_lut_4_lut.LUT_INIT = 16'hb2bb;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52192_3_lut (.I0(n32_adj_5177), .I1(baudrate[5]), .I2(n39_adj_5174), 
            .I3(GND_net), .O(n67920));   // verilog/uart_rx.v(119[33:55])
    defparam i52192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52193_3_lut (.I0(n67920), .I1(baudrate[6]), .I2(n41_adj_5173), 
            .I3(GND_net), .O(n67921));   // verilog/uart_rx.v(119[33:55])
    defparam i52193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51602_4_lut (.I0(n41_adj_5173), .I1(n39_adj_5174), .I2(n37_adj_5172), 
            .I3(n66435), .O(n67330));
    defparam i51602_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52266_3_lut (.I0(n34_adj_5178), .I1(baudrate[4]), .I2(n37_adj_5172), 
            .I3(GND_net), .O(n67994));   // verilog/uart_rx.v(119[33:55])
    defparam i52266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51335_3_lut (.I0(n67921), .I1(baudrate[7]), .I2(n43_adj_5171), 
            .I3(GND_net), .O(n67063));   // verilog/uart_rx.v(119[33:55])
    defparam i51335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5747_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11428));   // verilog/uart_rx.v(119[33:55])
    defparam i5747_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i52493_4_lut (.I0(n67063), .I1(n67994), .I2(n43_adj_5171), 
            .I3(n67330), .O(n68221));   // verilog/uart_rx.v(119[33:55])
    defparam i52493_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52494_3_lut (.I0(n68221), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n68222));   // verilog/uart_rx.v(119[33:55])
    defparam i52494_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n68222), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8035[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8035[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8035[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8035[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8035[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8035[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8035[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52196_3_lut (.I0(n34_adj_5183), .I1(baudrate[5]), .I2(n41_adj_5181), 
            .I3(GND_net), .O(n67924));   // verilog/uart_rx.v(119[33:55])
    defparam i52196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52197_3_lut (.I0(n67924), .I1(baudrate[6]), .I2(n43_adj_5179), 
            .I3(GND_net), .O(n67925));   // verilog/uart_rx.v(119[33:55])
    defparam i52197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51610_4_lut (.I0(n43_adj_5179), .I1(n41_adj_5181), .I2(n39_adj_5182), 
            .I3(n66445), .O(n67338));
    defparam i51610_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5184), .I1(baudrate[4]), 
            .I2(n39_adj_5182), .I3(GND_net), .O(n38_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51331_3_lut (.I0(n67925), .I1(baudrate[7]), .I2(n45_adj_5180), 
            .I3(GND_net), .O(n67059));   // verilog/uart_rx.v(119[33:55])
    defparam i51331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52260_4_lut (.I0(n67059), .I1(n38_adj_5185), .I2(n45_adj_5180), 
            .I3(n67338), .O(n67988));   // verilog/uart_rx.v(119[33:55])
    defparam i52260_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i42771_1_lut (.I0(n25657), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58457));
    defparam i42771_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1009 (.I0(n68447), .I1(baudrate[15]), .I2(n2353), 
            .I3(n60688), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1009.LUT_INIT = 16'h7100;
    SB_LUT4 i53688_2_lut_4_lut (.I0(n68447), .I1(baudrate[15]), .I2(n2353), 
            .I3(n62648), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i53688_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50747_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4937), .I3(\o_Rx_DV_N_3488[8] ), .O(n65682));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50747_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8009[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50863_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n57075), 
            .I3(r_SM_Main[0]), .O(n65688));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50863_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i50744_4_lut (.I0(n65682), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65679));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50744_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8009[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8009[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50750_4_lut (.I0(n65688), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65685));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50750_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n65685), .I1(n65679), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_5166));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8009[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8009[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8009[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5188), .I1(baudrate[4]), 
            .I2(n41_adj_5186), .I3(GND_net), .O(n40_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52633_4_lut (.I0(n40_adj_5189), .I1(n36_adj_5187), .I2(n41_adj_5186), 
            .I3(n66452), .O(n68361));   // verilog/uart_rx.v(119[33:55])
    defparam i52633_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52634_3_lut (.I0(n68361), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n68362));   // verilog/uart_rx.v(119[33:55])
    defparam i52634_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52496_3_lut (.I0(n68362), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n68224));   // verilog/uart_rx.v(119[33:55])
    defparam i52496_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46931_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25657), .I3(GND_net), .O(n58465));
    defparam i46931_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_4_lut_adj_1010 (.I0(n68346), .I1(baudrate[14]), .I2(n2227), 
            .I3(n60686), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1010.LUT_INIT = 16'h7100;
    SB_LUT4 i46885_1_lut_2_lut (.I0(baudrate[17]), .I1(n25657), .I2(GND_net), 
            .I3(GND_net), .O(n58461));
    defparam i46885_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_4_lut_adj_1011 (.I0(n68428), .I1(baudrate[18]), .I2(n2713), 
            .I3(n60694), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1011.LUT_INIT = 16'h7100;
    SB_LUT4 i53700_2_lut_4_lut (.I0(n68428), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25660), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i53700_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i42767_1_lut (.I0(n25660), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58453));
    defparam i42767_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5190));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4937), 
            .O(n15_adj_5191));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5191), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5190), 
            .I3(n57317), .O(n69846));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61158), .O(n61164));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61164), .O(n61170));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'hfffe;
    SB_LUT4 i52925_2_lut_3_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n27996));
    defparam i52925_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61142), .O(n61148));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61148), .O(n61154));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61078), .O(n61084));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61084), .O(n61090));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1018 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4940), 
            .I3(GND_net), .O(n60714));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_adj_1018.LUT_INIT = 16'hfefe;
    SB_LUT4 i5763_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n58926), .I3(n44_adj_5192), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i5763_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i742_4_lut (.I0(n58193), .I1(n294[18]), .I2(n46), .I3(baudrate[5]), 
            .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5193), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_3_lut_adj_1019 (.I0(n25605), .I1(n48_adj_5175), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1019.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1020 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n60714), .O(\r_SM_Main_2__N_3536[1] ));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 i7250_4_lut (.I0(n960), .I1(n11428), .I2(n21004), .I3(baudrate[3]), 
            .O(n21006));   // verilog/uart_rx.v(119[33:55])
    defparam i7250_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5192), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i5741_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam i5741_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i7249_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21004));   // verilog/uart_rx.v(119[33:55])
    defparam i7249_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5176), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5196), .I1(baudrate[4]), 
            .I2(n43_adj_5194), .I3(GND_net), .O(n42_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52621_4_lut (.I0(n42_adj_5197), .I1(n38_adj_5195), .I2(n43_adj_5194), 
            .I3(n66458), .O(n68349));   // verilog/uart_rx.v(119[33:55])
    defparam i52621_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52622_3_lut (.I0(n68349), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n68350));   // verilog/uart_rx.v(119[33:55])
    defparam i52622_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5592_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n58972), .I3(n44_adj_5198), 
            .O(n46_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam i5592_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i639_4_lut (.I0(n58191), .I1(n294[19]), .I2(n46_adj_5199), 
            .I3(baudrate[4]), .O(n58193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n62274));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5170), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i7243_4_lut (.I0(n804), .I1(n42960), .I2(n20994), .I3(baudrate[2]), 
            .O(n20996));   // verilog/uart_rx.v(119[33:55])
    defparam i7243_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5198), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i42763_1_lut (.I0(n25663), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58449));
    defparam i42763_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n62276));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1023 (.I0(n62166), .I1(n62162), .I2(n62164), 
            .I3(n62160), .O(n62146));
    defparam i1_4_lut_adj_1023.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1024 (.I0(n62274), .I1(n62030), .I2(n62158), 
            .I3(n62020), .O(n25666));
    defparam i1_4_lut_adj_1024.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n62012), .I1(n25666), .I2(n62146), 
            .I3(n62010), .O(n25605));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 i28999_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n58498));   // verilog/uart_rx.v(119[33:55])
    defparam i28999_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n58498), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52200_3_lut (.I0(n42_adj_5200), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n67928));   // verilog/uart_rx.v(119[33:55])
    defparam i52200_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52201_3_lut (.I0(n67928), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n67929));   // verilog/uart_rx.v(119[33:55])
    defparam i52201_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47150_1_lut (.I0(n62868), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58445));
    defparam i47150_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50695_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n66423));   // verilog/uart_rx.v(119[33:55])
    defparam i50695_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n67929), .I1(baudrate[5]), 
            .I2(n58193), .I3(GND_net), .O(n48_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53124_2_lut (.I0(n48_adj_5175), .I1(n25605), .I2(GND_net), 
            .I3(GND_net), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i53124_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i42755_1_lut (.I0(n25666), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58441));
    defparam i42755_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(n62276), .I1(n62278), .I2(n62114), 
            .I3(n62274), .O(n25670));
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1027 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4937), 
            .I3(\o_Rx_DV_N_3488[8] ), .O(n60672));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1028 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n60672), .O(r_SM_Main_2__N_3446[1]));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n61774));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_267_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5201));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(r_Clock_Count[3]), .I1(n3_adj_5201), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n61774), .O(n61778));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'hffde;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61062), .O(n61068));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_267_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61068), .O(n61074));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1033 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n61110), .O(n61116));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1033.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n61116), .O(n61122));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i534_3_lut (.I0(n58189), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n58191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n61778), .O(n61782));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'hffde;
    SB_LUT4 equal_267_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5202));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i535_4_lut (.I0(n68641), .I1(n44_adj_5169), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 i50904_4_lut (.I0(n25682), .I1(n65987), .I2(n48_adj_5159), 
            .I3(baudrate[0]), .O(n804));
    defparam i50904_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(r_Clock_Count[6]), .I1(n8_adj_5202), 
            .I2(n61782), .I3(\o_Rx_DV_N_3488[7] ), .O(n57075));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'hfdfe;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8399[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n60115));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i47147_2_lut (.I0(baudrate[8]), .I1(n62864), .I2(GND_net), 
            .I3(GND_net), .O(n62866));
    defparam i47147_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1037 (.I0(n25692), .I1(n48_adj_5168), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1037.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52202_3_lut (.I0(n42_adj_5203), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n67930));   // verilog/uart_rx.v(119[33:55])
    defparam i52202_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52203_3_lut (.I0(n67930), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n67931));   // verilog/uart_rx.v(119[33:55])
    defparam i52203_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n67931), .I1(baudrate[4]), 
            .I2(n58191), .I3(GND_net), .O(n48_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60115), .O(n60806));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60806), .O(n60812));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i47063_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n57075), .I2(GND_net), 
            .I3(GND_net), .O(n62782));
    defparam i47063_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8399[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47169_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n62782), .O(n62888));
    defparam i47169_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n60812), .I1(r_SM_Main_2__N_3446[1]), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n62888), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n11645));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n11645), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8399[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8399[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53159_2_lut_4_lut (.I0(n68220), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25636), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i53159_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8399[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8399[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8399[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46884_2_lut (.I0(baudrate[17]), .I1(n25657), .I2(GND_net), 
            .I3(GND_net), .O(n62602));
    defparam i46884_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1040 (.I0(n62010), .I1(n62166), .I2(baudrate[16]), 
            .I3(n42960), .O(n61274));
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'h0100;
    SB_LUT4 i50985_3_lut (.I0(n58984), .I1(n59856), .I2(baudrate[2]), 
            .I3(GND_net), .O(n65628));   // verilog/uart_rx.v(119[33:55])
    defparam i50985_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i50847_4_lut (.I0(n58258), .I1(n61274), .I2(n62012), .I3(n61328), 
            .O(n65629));   // verilog/uart_rx.v(119[33:55])
    defparam i50847_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n65629), .I1(n65628), .I2(n294[21]), 
            .I3(n62602), .O(n58189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n62272));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n61008));
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'h0100;
    SB_LUT4 i47107_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n62826));
    defparam i47107_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(n58258), .I1(n61008), .I2(n62272), 
            .I3(baudrate[16]), .O(n61036));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h0004;
    SB_LUT4 i47177_4_lut (.I0(n62826), .I1(n62748), .I2(n62752), .I3(n62586), 
            .O(n62896));
    defparam i47177_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52913_4_lut (.I0(n62884), .I1(n65985), .I2(n62896), .I3(n61036), 
            .O(n68641));
    defparam i52913_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n62164));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n61356));
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1046 (.I0(n61356), .I1(n62172), .I2(n62134), 
            .I3(GND_net), .O(n25663));
    defparam i1_3_lut_adj_1046.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n62004));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n62002));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n61328));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1050 (.I0(n61328), .I1(n62002), .I2(n62004), 
            .I3(n62000), .O(n61340));
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1051 (.I0(n61340), .I1(n25663), .I2(n61332), 
            .I3(n62174), .O(n25692));
    defparam i1_4_lut_adj_1051.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n65705), .I1(baudrate[2]), 
            .I2(n68641), .I3(n48_adj_5159), .O(n46_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5204), .I1(baudrate[3]), 
            .I2(n58189), .I3(GND_net), .O(n48_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53121_2_lut (.I0(n48_adj_5168), .I1(n25692), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i53121_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n62162));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n62166));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n61998));
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n62000));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'heeee;
    SB_LUT4 i47043_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n62762));
    defparam i47043_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47165_4_lut (.I0(n62762), .I1(n61332), .I2(n62000), .I3(baudrate[9]), 
            .O(n62884));
    defparam i47165_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28992_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42962));
    defparam i28992_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28990_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42960));
    defparam i28990_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n62172), .I1(n60660), .I2(n60658), 
            .I3(n62162), .O(n25657));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1057 (.I0(baudrate[17]), .I1(n62788), .I2(baudrate[2]), 
            .I3(n42960), .O(n60618));
    defparam i1_4_lut_adj_1057.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(n62838), .I1(n60618), .I2(n25657), 
            .I3(n62748), .O(n59856));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8399[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1059 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n42962), .O(n60952));
    defparam i1_4_lut_adj_1059.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1060 (.I0(n60952), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n60970));
    defparam i1_4_lut_adj_1060.LUT_INIT = 16'h0002;
    SB_LUT4 i47179_4_lut (.I0(n62832), .I1(n62748), .I2(n62752), .I3(n62586), 
            .O(n62898));
    defparam i47179_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8399[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n62884), .I1(n62898), .I2(n58258), 
            .I3(n60970), .O(n58984));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n58984), .I1(baudrate[2]), 
            .I2(n59856), .I3(GND_net), .O(n48_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53707_2_lut (.I0(n48_adj_5159), .I1(n25682), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i53707_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_3_lut_4_lut_adj_1062 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61094));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1062.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut_4_lut_adj_1063 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61046));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1063.LUT_INIT = 16'hffbf;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8399[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n62112));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'heeee;
    SB_LUT4 i42574_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n58258));
    defparam i42574_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47089_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n62808));
    defparam i47089_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i47149_4_lut (.I0(n62808), .I1(n62158), .I2(n62806), .I3(n62112), 
            .O(n62868));
    defparam i47149_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46867_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62584));
    defparam i46867_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47119_4_lut (.I0(n61192), .I1(n61188), .I2(n61190), .I3(n61186), 
            .O(n62838));
    defparam i47119_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47183_4_lut (.I0(n62868), .I1(n62748), .I2(n58258), .I3(baudrate[4]), 
            .O(n62902));
    defparam i47183_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52942_4_lut (.I0(n62838), .I1(n62586), .I2(n62902), .I3(n62584), 
            .O(n62906));
    defparam i52942_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_1065 (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[2] ), .I3(GND_net), .O(n4));
    defparam i1_2_lut_3_lut_adj_1065.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8399[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8399[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8399[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8399[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1066 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n60658));
    defparam i1_3_lut_4_lut_adj_1066.LUT_INIT = 16'hfffe;
    SB_LUT4 i47113_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n62832));
    defparam i47113_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47148_1_lut_2_lut (.I0(baudrate[8]), .I1(n62864), .I2(GND_net), 
            .I3(GND_net), .O(n58491));
    defparam i47148_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8399[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8399[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8425[20]), .I3(n294[1]), .O(n41_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8399[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8425[19]), .I3(n294[1]), .O(n39_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8425[17]), .I3(n294[1]), .O(n35_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8425[18]), .I3(n294[1]), .O(n37_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8425[14]), .I3(n294[1]), .O(n29_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8425[15]), .I3(n294[1]), .O(n31_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8399[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50304_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n66032));
    defparam i50304_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8425[11]), .I3(n294[1]), .O(n23_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8425[12]), .I3(n294[1]), .O(n25_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i50337_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n66065));
    defparam i50337_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8425[16]), .I3(n294[1]), .O(n33_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8425[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8399[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8399[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8373[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8425[21]), .I3(n294[1]), .O(n43_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8425[22]), .I3(n294[1]), .O(n45_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8373[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8373[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8373[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8373[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8373[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8425[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i50410_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n66138));
    defparam i50410_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8373[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8373[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8425[8]), .I3(n294[1]), .O(n17_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8373[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8425[9]), .I3(n294[1]), .O(n19_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8373[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8373[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50377_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n66105));
    defparam i50377_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8373[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50450_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n66178));
    defparam i50450_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8425[10]), .I3(n294[1]), .O(n21_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50429_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n66157));
    defparam i50429_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8373[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8373[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50541_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n66269));
    defparam i50541_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8425[5]), .I3(n294[1]), .O(n11_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8373[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50547_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n66275));
    defparam i50547_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1067 (.I0(n61196), .I1(n62870), .I2(baudrate[0]), 
            .I3(n48_adj_5152), .O(n962));
    defparam i1_3_lut_4_lut_adj_1067.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8425[6]), .I3(n294[1]), .O(n13_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8425[7]), .I3(n294[1]), .O(n15_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8373[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8373[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50575_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n66303));
    defparam i50575_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8347[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8347[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1068 (.I0(n62000), .I1(n62840), .I2(n8087[14]), 
            .I3(n48_adj_5151), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1068.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8425[13]), .I3(n294[1]), .O(n27_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8347[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8347[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(baudrate[24]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n62118));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n62160));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n62116));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n61214));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n62020));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62158));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'heeee;
    SB_LUT4 i50195_4_lut (.I0(n27_adj_5222), .I1(n15_adj_5221), .I2(n13_adj_5220), 
            .I3(n11_adj_5219), .O(n65923));
    defparam i50195_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n62158), .I1(n62020), .I2(n61214), 
            .I3(baudrate[19]), .O(n61234));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8347[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1076 (.I0(n61234), .I1(n62116), .I2(n62160), 
            .I3(n62118), .O(n25660));
    defparam i1_4_lut_adj_1076.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n62586));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut_adj_1078 (.I0(n61188), .I1(n62650), .I2(n8165[11]), 
            .I3(n48_adj_5024), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1078.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8347[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n61188));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n61186));
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n61190));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n61192));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n61196));
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'heeee;
    SB_LUT4 i50203_4_lut (.I0(n21_adj_5218), .I1(n19_adj_5217), .I2(n17_adj_5216), 
            .I3(n9), .O(n65931));
    defparam i50203_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8347[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5214), .I3(GND_net), .O(n16_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8347[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n61194));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8347[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47069_2_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n62788));
    defparam i47069_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1085 (.I0(n61190), .I1(n61186), .I2(n61188), 
            .I3(n62586), .O(n61208));
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(n62788), .I1(n61194), .I2(n61196), 
            .I3(n61192), .O(n61210));
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8347[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1087 (.I0(n61210), .I1(n25660), .I2(n61208), 
            .I3(GND_net), .O(n25682));
    defparam i1_3_lut_adj_1087.LUT_INIT = 16'hfefe;
    SB_LUT4 i50164_2_lut (.I0(n43_adj_5214), .I1(n19_adj_5217), .I2(GND_net), 
            .I3(GND_net), .O(n65892));
    defparam i50164_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53051_3_lut (.I0(n25682), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25593));   // verilog/uart_rx.v(119[33:55])
    defparam i53051_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8347[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8347[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5216), .I3(GND_net), .O(n8_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8347[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5223), .I1(baudrate[22]), 
            .I2(n45_adj_5215), .I3(GND_net), .O(n24_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8347[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8425[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8347[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50217_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n65945));
    defparam i50217_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8347[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8347[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8321[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50579_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n66307));
    defparam i50579_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8321[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8321[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51091_4_lut (.I0(n13_adj_5220), .I1(n11_adj_5219), .I2(n9), 
            .I3(n65945), .O(n66819));
    defparam i51091_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51087_4_lut (.I0(n19_adj_5217), .I1(n17_adj_5216), .I2(n15_adj_5221), 
            .I3(n66819), .O(n66815));
    defparam i51087_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8321[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50595_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n66323));
    defparam i50595_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8321[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52451_4_lut (.I0(n25_adj_5212), .I1(n23_adj_5211), .I2(n21_adj_5218), 
            .I3(n66815), .O(n68179));
    defparam i52451_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51830_4_lut (.I0(n31_adj_5210), .I1(n29_adj_5209), .I2(n27_adj_5222), 
            .I3(n68179), .O(n67558));
    defparam i51830_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8321[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8321[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52670_4_lut (.I0(n37_adj_5208), .I1(n35_adj_5207), .I2(n33_adj_5213), 
            .I3(n67558), .O(n68398));
    defparam i52670_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8321[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8321[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5213), .I3(GND_net), .O(n12_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8321[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8321[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50601_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n66329));
    defparam i50601_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n60702), .I3(n48_adj_4993), .O(n4_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52385_3_lut (.I0(n4_adj_5227), .I1(baudrate[13]), .I2(n27_adj_5222), 
            .I3(GND_net), .O(n68113));   // verilog/uart_rx.v(119[33:55])
    defparam i52385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52386_3_lut (.I0(n68113), .I1(baudrate[14]), .I2(n29_adj_5209), 
            .I3(GND_net), .O(n68114));   // verilog/uart_rx.v(119[33:55])
    defparam i52386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1088 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61062));
    defparam i1_3_lut_4_lut_adj_1088.LUT_INIT = 16'hfff7;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_1089 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61110));
    defparam i1_3_lut_4_lut_adj_1089.LUT_INIT = 16'hff7f;
    SB_LUT4 i50618_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n66346));
    defparam i50618_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50185_2_lut (.I0(n33_adj_5213), .I1(n15_adj_5221), .I2(GND_net), 
            .I3(GND_net), .O(n65913));
    defparam i50185_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8321[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8321[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_5220), .I3(GND_net), .O(n10_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8321[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8321[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50622_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n66350));
    defparam i50622_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_5226), .I1(baudrate[17]), 
            .I2(n35_adj_5207), .I3(GND_net), .O(n30_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1090 (.I0(baudrate[2]), .I1(n42_adj_5170), 
            .I2(baudrate[3]), .I3(n20996), .O(n58972));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1090.LUT_INIT = 16'hff4f;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8321[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8295[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8269[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8295[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53193_2_lut_4_lut (.I0(n68483), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25645), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i53193_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i5585_2_lut_3_lut (.I0(baudrate[2]), .I1(n42_adj_5170), .I2(n20996), 
            .I3(GND_net), .O(n44_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam i5585_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 i1_2_lut_4_lut_adj_1091 (.I0(n68350), .I1(baudrate[6]), .I2(n1111), 
            .I3(n60678), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1091.LUT_INIT = 16'h7100;
    SB_LUT4 i53664_2_lut_4_lut (.I0(n68350), .I1(baudrate[6]), .I2(n1111), 
            .I3(n62870), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i53664_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i50730_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n66458));   // verilog/uart_rx.v(119[33:55])
    defparam i50730_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i53685_2_lut_4_lut (.I0(n68346), .I1(baudrate[14]), .I2(n2227), 
            .I3(n62650), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i53685_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut_adj_1092 (.I0(baudrate[3]), .I1(n42_adj_5176), 
            .I2(baudrate[4]), .I3(n21006), .O(n58926));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1092.LUT_INIT = 16'hff4f;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8295[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50187_4_lut (.I0(n33_adj_5213), .I1(n31_adj_5210), .I2(n29_adj_5209), 
            .I3(n65923), .O(n65915));
    defparam i50187_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i5756_2_lut_3_lut (.I0(baudrate[3]), .I1(n42_adj_5176), .I2(n21006), 
            .I3(GND_net), .O(n44_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam i5756_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8295[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8295[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52736_4_lut (.I0(n30_adj_5229), .I1(n10_adj_5228), .I2(n35_adj_5207), 
            .I3(n65913), .O(n68464));   // verilog/uart_rx.v(119[33:55])
    defparam i52736_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_3_lut_4_lut_adj_1093 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61142));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1093.LUT_INIT = 16'hfffd;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8295[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1094 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61078));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1094.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1095 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61158));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1095.LUT_INIT = 16'hffef;
    SB_LUT4 i50653_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n66381));
    defparam i50653_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52316_3_lut (.I0(n68114), .I1(baudrate[15]), .I2(n31_adj_5210), 
            .I3(GND_net), .O(n68044));   // verilog/uart_rx.v(119[33:55])
    defparam i52316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1096 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n61126));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1096.LUT_INIT = 16'hfffe;
    SB_LUT4 i52854_4_lut (.I0(n68044), .I1(n68464), .I2(n35_adj_5207), 
            .I3(n65915), .O(n68582));   // verilog/uart_rx.v(119[33:55])
    defparam i52854_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8295[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52855_3_lut (.I0(n68582), .I1(baudrate[18]), .I2(n37_adj_5208), 
            .I3(GND_net), .O(n68583));   // verilog/uart_rx.v(119[33:55])
    defparam i52855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8295[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8295[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8295[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1097 (.I0(n68534), .I1(baudrate[11]), .I2(n1831), 
            .I3(n60684), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1097.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8295[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52389_3_lut (.I0(n6_adj_5236), .I1(baudrate[10]), .I2(n21_adj_5218), 
            .I3(GND_net), .O(n68117));   // verilog/uart_rx.v(119[33:55])
    defparam i52389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8295[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8295[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52390_3_lut (.I0(n68117), .I1(baudrate[11]), .I2(n23_adj_5211), 
            .I3(GND_net), .O(n68118));   // verilog/uart_rx.v(119[33:55])
    defparam i52390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8295[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5020));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8295[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5015));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50169_4_lut (.I0(n43_adj_5214), .I1(n25_adj_5212), .I2(n23_adj_5211), 
            .I3(n65931), .O(n65897));
    defparam i50169_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8295[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50670_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n66398));
    defparam i50670_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51952_4_lut (.I0(n24_adj_5225), .I1(n8_adj_5224), .I2(n45_adj_5215), 
            .I3(n65892), .O(n67680));   // verilog/uart_rx.v(119[33:55])
    defparam i51952_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8295[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52314_3_lut (.I0(n68118), .I1(baudrate[12]), .I2(n25_adj_5212), 
            .I3(GND_net), .O(n68042));   // verilog/uart_rx.v(119[33:55])
    defparam i52314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50476_4_lut (.I0(n37_adj_5245), .I1(n25_adj_5244), .I2(n23_adj_5243), 
            .I3(n21_adj_5242), .O(n66204));
    defparam i50476_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51436_4_lut (.I0(n19_adj_5241), .I1(n17_adj_5240), .I2(n2729), 
            .I3(baudrate[2]), .O(n67164));
    defparam i51436_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52796_3_lut (.I0(n68583), .I1(baudrate[19]), .I2(n39_adj_5206), 
            .I3(GND_net), .O(n68524));   // verilog/uart_rx.v(119[33:55])
    defparam i52796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50171_4_lut (.I0(n43_adj_5214), .I1(n41_adj_5205), .I2(n39_adj_5206), 
            .I3(n68398), .O(n65899));
    defparam i50171_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51974_4_lut (.I0(n25_adj_5244), .I1(n23_adj_5243), .I2(n21_adj_5242), 
            .I3(n67164), .O(n67702));
    defparam i51974_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51970_4_lut (.I0(n31_adj_5239), .I1(n29_adj_5238), .I2(n27_adj_5237), 
            .I3(n67702), .O(n67698));
    defparam i51970_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50478_4_lut (.I0(n37_adj_5245), .I1(n35_adj_5235), .I2(n33_adj_5234), 
            .I3(n67698), .O(n66206));
    defparam i50478_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50635_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n66363));
    defparam i50635_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52555_4_lut (.I0(n68042), .I1(n67680), .I2(n45_adj_5215), 
            .I3(n65897), .O(n68283));   // verilog/uart_rx.v(119[33:55])
    defparam i52555_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52140_3_lut (.I0(n14_adj_5246), .I1(baudrate[13]), .I2(n37_adj_5245), 
            .I3(GND_net), .O(n67868));   // verilog/uart_rx.v(119[33:55])
    defparam i52140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52788_3_lut (.I0(n68524), .I1(baudrate[20]), .I2(n41_adj_5205), 
            .I3(GND_net), .O(n40_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam i52788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52141_3_lut (.I0(n67868), .I1(baudrate[14]), .I2(n39_adj_5232), 
            .I3(GND_net), .O(n67869));   // verilog/uart_rx.v(119[33:55])
    defparam i52141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_5150), .I1(baudrate[17]), 
            .I2(n45_adj_5231), .I3(GND_net), .O(n40_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50472_4_lut (.I0(n43_adj_5233), .I1(n41_adj_5230), .I2(n39_adj_5232), 
            .I3(n66204), .O(n66200));
    defparam i50472_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52283_4_lut (.I0(n40_adj_5248), .I1(n20_adj_5149), .I2(n45_adj_5231), 
            .I3(n66196), .O(n68011));   // verilog/uart_rx.v(119[33:55])
    defparam i52283_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n60630));
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'heeee;
    SB_LUT4 i51395_3_lut (.I0(n67869), .I1(baudrate[15]), .I2(n41_adj_5230), 
            .I3(GND_net), .O(n67123));   // verilog/uart_rx.v(119[33:55])
    defparam i51395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8425[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5148), .I1(baudrate[9]), 
            .I2(n29_adj_5238), .I3(GND_net), .O(n26_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52557_4_lut (.I0(n40_adj_5247), .I1(n68283), .I2(n45_adj_5215), 
            .I3(n65899), .O(n68285));   // verilog/uart_rx.v(119[33:55])
    defparam i52557_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52653_4_lut (.I0(n26_adj_5249), .I1(n16_adj_5147), .I2(n29_adj_5238), 
            .I3(n66219), .O(n68381));   // verilog/uart_rx.v(119[33:55])
    defparam i52653_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52654_3_lut (.I0(n68381), .I1(baudrate[10]), .I2(n31_adj_5239), 
            .I3(GND_net), .O(n68382));   // verilog/uart_rx.v(119[33:55])
    defparam i52654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52448_3_lut (.I0(n68382), .I1(baudrate[11]), .I2(n33_adj_5234), 
            .I3(GND_net), .O(n68176));   // verilog/uart_rx.v(119[33:55])
    defparam i52448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1099 (.I0(n62272), .I1(n62118), .I2(n60630), 
            .I3(n62114), .O(n60638));
    defparam i1_4_lut_adj_1099.LUT_INIT = 16'hfffe;
    SB_LUT4 i53252_4_lut (.I0(n60638), .I1(n68285), .I2(baudrate[23]), 
            .I3(n3253), .O(n59626));   // verilog/uart_rx.v(119[33:55])
    defparam i53252_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 i52325_4_lut (.I0(n43_adj_5233), .I1(n41_adj_5230), .I2(n39_adj_5232), 
            .I3(n66206), .O(n68053));
    defparam i52325_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52698_4_lut (.I0(n67123), .I1(n68011), .I2(n45_adj_5231), 
            .I3(n66200), .O(n68426));   // verilog/uart_rx.v(119[33:55])
    defparam i52698_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51393_3_lut (.I0(n68176), .I1(baudrate[12]), .I2(n35_adj_5235), 
            .I3(GND_net), .O(n67121));   // verilog/uart_rx.v(119[33:55])
    defparam i51393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52700_4_lut (.I0(n67121), .I1(n68426), .I2(n45_adj_5231), 
            .I3(n68053), .O(n68428));   // verilog/uart_rx.v(119[33:55])
    defparam i52700_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8269[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8269[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8269[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8269[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8269[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53725_2_lut_4_lut (.I0(n68395), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25670), .O(n294[1]));
    defparam i53725_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8269[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8269[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8269[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1100 (.I0(n68224), .I1(baudrate[7]), .I2(n1261), 
            .I3(n60680), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1100.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5070));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8269[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8269[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8269[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8269[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8269[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53670_2_lut_4_lut (.I0(n68224), .I1(baudrate[7]), .I2(n1261), 
            .I3(n62866), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i53670_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8269[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50724_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n66452));   // verilog/uart_rx.v(119[33:55])
    defparam i50724_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1101 (.I0(n67988), .I1(baudrate[8]), .I2(n1408), 
            .I3(n60682), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1101.LUT_INIT = 16'h7100;
    SB_LUT4 i53673_2_lut_4_lut (.I0(n67988), .I1(baudrate[8]), .I2(n1408), 
            .I3(n62864), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i53673_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50717_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n66445));   // verilog/uart_rx.v(119[33:55])
    defparam i50717_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8243[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8243[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8243[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8243[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53679_2_lut_4_lut (.I0(n68534), .I1(baudrate[11]), .I2(n1831), 
            .I3(n62840), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i53679_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8243[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50707_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n66435));   // verilog/uart_rx.v(119[33:55])
    defparam i50707_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8243[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8243[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8243[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8243[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8243[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50245_4_lut (.I0(n29_adj_5256), .I1(n17_adj_5255), .I2(n15_adj_5254), 
            .I3(n13_adj_5253), .O(n65973));
    defparam i50245_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8243[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8243[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47121_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n62650), .I3(baudrate[12]), .O(n62840));
    defparam i47121_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53682_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n62650), .I3(n48_adj_5024), .O(n294[11]));
    defparam i53682_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8217[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8217[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46932_2_lut_4_lut (.I0(baudrate[15]), .I1(baudrate[16]), .I2(baudrate[17]), 
            .I3(n25657), .O(n62650));
    defparam i46932_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8217[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8217[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51182_4_lut (.I0(n11_adj_5251), .I1(n9_adj_5250), .I2(n3171), 
            .I3(baudrate[2]), .O(n66910));
    defparam i51182_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8217[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51866_4_lut (.I0(n17_adj_5255), .I1(n15_adj_5254), .I2(n13_adj_5253), 
            .I3(n66910), .O(n67594));
    defparam i51866_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8217[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51864_4_lut (.I0(n23_c), .I1(n21), .I2(n19_adj_5252), .I3(n67594), 
            .O(n67592));
    defparam i51864_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50252_4_lut (.I0(n29_adj_5256), .I1(n27_c), .I2(n25), .I3(n67592), 
            .O(n65980));
    defparam i50252_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8217[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8217[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8217[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52395_3_lut (.I0(n6_adj_5257), .I1(baudrate[13]), .I2(n29_adj_5256), 
            .I3(GND_net), .O(n68123));   // verilog/uart_rx.v(119[33:55])
    defparam i52395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50230_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n65958));
    defparam i50230_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[10] , \PID_CONTROLLER.integral_23__N_3715[0] , 
            GND_net, \Ki[11] , \Ki[12] , \Ki[13] , \Kp[0] , \Kp[1] , 
            \Ki[14] , n365, control_update, duty, clk16MHz, reset, 
            IntegralLimit, n155, \Kp[5] , PWMLimit, \Kp[6] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[7] , \Kp[12] , \Kp[8] , \Kp[13] , 
            \Ki[1] , \PID_CONTROLLER.integral_23__N_3715[16] , \Ki[15] , 
            \Ki[2] , \Ki[3] , \Kp[14] , \Ki[4] , \Kp[15] , \Ki[5] , 
            \Ki[6] , \Ki[7] , \Kp[3] , deadband, n380, n379, setpoint, 
            \motor_state[10] , \motor_state[9] , \motor_state[8] , \motor_state[7] , 
            n41756, \PID_CONTROLLER.integral_23__N_3715[23] , \motor_state[5] , 
            \Kp[2] , \Kp[4] , \motor_state[4] , n42305, \motor_state[2] , 
            \PID_CONTROLLER.integral_23__N_3715[22] , \PID_CONTROLLER.integral_23__N_3715[21] , 
            \PID_CONTROLLER.integral_23__N_3715[20] , n212, n213, n214, 
            \motor_state[1] , n4, n37308, n11610, \PID_CONTROLLER.integral_23__N_3715[15] , 
            \PID_CONTROLLER.integral_23__N_3715[14] , \Ki[0] , \motor_state[0] , 
            VCC_net, \Ki[8] , \PID_CONTROLLER.integral , \Ki[9] , n38, 
            n29669, n110, n30497, n30496, n30495, n30494, n30493, 
            n30491, n30489, n30488, n30487, n30486, n30485, n30484, 
            n30483, n30482, n30481, n30480, n30479, n30478, n30477, 
            n30476, n30475, n30474, n30473, \PID_CONTROLLER.integral_23__N_3715[13] , 
            \PID_CONTROLLER.integral_23__N_3715[12] , n27722, n53, n459, 
            n460, \motor_state[23] , \motor_state[22] , \motor_state[21] , 
            n219, \motor_state[20] , \PID_CONTROLLER.integral_23__N_3715[11] , 
            \motor_state[19] , n490, n417, \motor_state[18] , n20203, 
            n344, \motor_state[17] , n20204, n271, n20205, n198, 
            n56, n125, n20, \motor_state[15] , \motor_state[14] , 
            n405, \motor_state[13] , \motor_state[12] , n43, \motor_state[11] , 
            \PID_CONTROLLER.integral_23__N_3715[10] , n4_adj_7, n30, \PID_CONTROLLER.integral_23__N_3715[9] , 
            \PID_CONTROLLER.integral_23__N_3715[8] , \PID_CONTROLLER.integral_23__N_3715[7] , 
            \PID_CONTROLLER.integral_23__N_3715[6] , n6, n36852, n4_adj_8, 
            n36823, \PID_CONTROLLER.integral_23__N_3715[5] , \PID_CONTROLLER.integral_23__N_3715[4] , 
            \PID_CONTROLLER.integral_23__N_3715[3] , \PID_CONTROLLER.integral_23__N_3715[2] , 
            \PID_CONTROLLER.integral_23__N_3715[1] , n43450, n20253, n49420, 
            n20283, n35, n4_adj_9, n32) /* synthesis syn_module_defined=1 */ ;
    input \Ki[10] ;
    output \PID_CONTROLLER.integral_23__N_3715[0] ;
    input GND_net;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Kp[0] ;
    input \Kp[1] ;
    input \Ki[14] ;
    output n365;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input [23:0]IntegralLimit;
    output n155;
    input \Kp[5] ;
    input [23:0]PWMLimit;
    input \Kp[6] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[7] ;
    input \Kp[12] ;
    input \Kp[8] ;
    input \Kp[13] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.integral_23__N_3715[16] ;
    input \Ki[15] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Kp[14] ;
    input \Ki[4] ;
    input \Kp[15] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Kp[3] ;
    input [23:0]deadband;
    output n380;
    output n379;
    input [23:0]setpoint;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input n41756;
    output \PID_CONTROLLER.integral_23__N_3715[23] ;
    input \motor_state[5] ;
    input \Kp[2] ;
    input \Kp[4] ;
    input \motor_state[4] ;
    input n42305;
    input \motor_state[2] ;
    output \PID_CONTROLLER.integral_23__N_3715[22] ;
    output \PID_CONTROLLER.integral_23__N_3715[21] ;
    output \PID_CONTROLLER.integral_23__N_3715[20] ;
    output n212;
    output n213;
    output n214;
    input \motor_state[1] ;
    input n4;
    input n37308;
    output n11610;
    output \PID_CONTROLLER.integral_23__N_3715[15] ;
    output \PID_CONTROLLER.integral_23__N_3715[14] ;
    input \Ki[0] ;
    input \motor_state[0] ;
    input VCC_net;
    input \Ki[8] ;
    output [23:0]\PID_CONTROLLER.integral ;
    input \Ki[9] ;
    input n38;
    input n29669;
    input n110;
    input n30497;
    input n30496;
    input n30495;
    input n30494;
    input n30493;
    input n30491;
    input n30489;
    input n30488;
    input n30487;
    input n30486;
    input n30485;
    input n30484;
    input n30483;
    input n30482;
    input n30481;
    input n30480;
    input n30479;
    input n30478;
    input n30477;
    input n30476;
    input n30475;
    input n30474;
    input n30473;
    output \PID_CONTROLLER.integral_23__N_3715[13] ;
    input \PID_CONTROLLER.integral_23__N_3715[12] ;
    input n27722;
    input n53;
    output n459;
    output n460;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    output n219;
    input \motor_state[20] ;
    output \PID_CONTROLLER.integral_23__N_3715[11] ;
    input \motor_state[19] ;
    input n490;
    input n417;
    input \motor_state[18] ;
    input n20203;
    input n344;
    input \motor_state[17] ;
    input n20204;
    input n271;
    input n20205;
    input n198;
    input n56;
    input n125;
    input n20;
    input \motor_state[15] ;
    input \motor_state[14] ;
    output n405;
    input \motor_state[13] ;
    input \motor_state[12] ;
    output n43;
    input \motor_state[11] ;
    output \PID_CONTROLLER.integral_23__N_3715[10] ;
    input n4_adj_7;
    output n30;
    output \PID_CONTROLLER.integral_23__N_3715[9] ;
    output \PID_CONTROLLER.integral_23__N_3715[8] ;
    output \PID_CONTROLLER.integral_23__N_3715[7] ;
    output \PID_CONTROLLER.integral_23__N_3715[6] ;
    input n6;
    input n36852;
    input n4_adj_8;
    input n36823;
    output \PID_CONTROLLER.integral_23__N_3715[5] ;
    output \PID_CONTROLLER.integral_23__N_3715[4] ;
    output \PID_CONTROLLER.integral_23__N_3715[3] ;
    output \PID_CONTROLLER.integral_23__N_3715[2] ;
    output \PID_CONTROLLER.integral_23__N_3715[1] ;
    output n43450;
    output n20253;
    output n49420;
    output n20283;
    output n35;
    input n4_adj_9;
    input n32;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n731, n804, n877, n49623;
    wire [47:0]n257;
    wire [47:0]n306;
    
    wire n49624;
    wire [10:0]n19161;
    wire [9:0]n19425;
    
    wire n767, n49810, n950;
    wire [23:0]n356;
    wire [23:0]n382;
    
    wire n69902;
    wire [23:0]n1;
    wire [4:0]n20165;
    
    wire n1023, n49338, n66659, n67830, n69928, n68339;
    wire [23:0]n49;
    
    wire n49622, n49695;
    wire [23:0]n1_adj_4984;
    
    wire n49696;
    wire [17:0]n15745;
    wire [16:0]n16429;
    
    wire n527, n50005;
    wire [23:0]n130;
    wire [23:0]n182;
    
    wire n181;
    wire [23:0]n207;
    
    wire n375;
    wire [23:0]n1_adj_4985;
    
    wire n448, n688, n761, n834, n521, n907, n594, n980, n122, 
        n1096, n667, n195, n268, n740, n813, n886, n959, n1032, 
        n341, n1105, n95, n414, n26, n487, n560, n69893, n68551, 
        n69890, n19, n10;
    wire [2:0]n20265;
    
    wire n4_adj_4449;
    wire [3:0]n20225;
    
    wire n11, n9, n66734, n17_adj_4450, n15_adj_4451, n13_adj_4452, 
        n67520, n23, n21, n67518, n6_c, n62, n131, n204, n50006, 
        n49811, n49694, n29, n27, n25, n66714, n65620, n454, 
        n50004, n6_adj_4453, n694, n49809, n381, n50003, n308, 
        n50002, n49693, n621, n49808, n67986, n35_c, n14_adj_4455, 
        counter_31__N_3714, n235, n50001, n49568, n49569, n12_adj_4456, 
        n49692, n548, n49807, n37, n32_c, n162, n50000, n49567, 
        n66710, n49621, n66569, n34, n475, n49806, n49691, n31, 
        n67987, n20_c, n89, n49566, n33, n66701, n49690, n402, 
        n49805, n49565, n329, n49804, n49620, n49689, n256, n49803, 
        n66696, n68351, n49564, n66862, n6_adj_4460, n183, n49802, 
        n49688, n67976, n41, n110_adj_4462, n734, n49619, n49687, 
        n831, n49686, n904, n49563, n49618, n49685, n49684, n168, 
        n241, n314, n387_adj_4470, n460_c, n533, n606, n679, n752, 
        n825, n49617, n49562;
    wire [8:0]n19744;
    wire [7:0]n19905;
    
    wire n700, n49986, n49683, n627, n49985, n49682, n898, n49616, 
        n971, n554, n49984, n1044, n1117, n481, n49983, n408, 
        n49982, n49615, n49561, n335_adj_4476, n49981, n49681, n262, 
        n49980, n67977, n49560, n189_adj_4478, n49979, n47, n116, 
        n49680;
    wire [15:0]n17041;
    
    wire n49978, n49977, n49614, n1114, n49976, n49559, n49679, 
        n1041, n49975, n67974, n92, n23_adj_4485, n165, n968, 
        n49974, n60589, n11608, n238, n311, n895, n49973, n384, 
        n457, n822, n49972, n530, n67975, n69898, n67476, n66649, 
        n749, n49971, n676, n49970, n69924, n603, n49969, n49968, 
        n49967, n30_c, n10_adj_4486, n66637, n68416;
    wire [23:0]n436;
    
    wire n27922, n49966, n49965, n49964, n66872, n49963, n49678, 
        n27917, n27912, n68537, n68538, n68499, n69912, n67482, 
        n66613, n24_adj_4488, n8_adj_4489, n69888, n66611, n67584, 
        n49613, n66870, n66615, n68211, n27907, n66878, n27902, 
        n49677, n49612, n27897, n49611, n49676, n27892, n27887;
    wire [14:0]n17585;
    
    wire n49950, n49610, n49949, n49948, n49947, n49675, n49946, 
        n41_adj_4494, n39, n49945, n49944, n49943, n45, n37_adj_4495, 
        n49942, n23_adj_4496, n8_adj_4497, n67990, n67991, n65796, 
        n66720, n67582, n66860, n68115, n68535, n68153, n68596, 
        n68597, n68451, n68365, n68366, n68406, n62222, n47_adj_4498, 
        n49941, n49940, n49609, n49939, n67963, n49938, n25_adj_4499, 
        n43_c, n29_adj_4500, n31_adj_4501, n35_adj_4502, n33_adj_4503, 
        n11_adj_4504, n49937, n49936, n27882;
    wire [0:0]n12229;
    wire [21:0]n12736;
    
    wire n51238, n51237, n51236, n51235, n51234, n51233, n51232, 
        n51231, n51230, n27877, n51229, n51228, n51227, n49608, 
        n51226, n51225, n658, n51224, n585, n51223, n512, n51222, 
        n439, n51221, n366_adj_4505, n51220, n293_adj_4506, n51219, 
        n220, n51218, n27872, n147, n51217, n5_adj_4508, n74;
    wire [20:0]n13704;
    
    wire n51216, n51215, n51214, n51213, n51212, n51211, n51210, 
        n13_adj_4509, n1099, n51209, n15_adj_4511, n1026, n51208, 
        n953, n51207, n880, n51206, n807, n51205, n734_adj_4512, 
        n51204, n661, n51203, n588, n51202, n515, n51201, n442, 
        n51200, n27_adj_4513, n369_adj_4514, n51199, n296_adj_4515, 
        n51198, n223, n51197, n150, n51196, n9_adj_4517, n8_adj_4518, 
        n77;
    wire [19:0]n14585;
    
    wire n51195, n51194, n17_adj_4519, n51193, n51192, n51191, n51190, 
        n1102, n51189, n1029, n51188, n19_adj_4520, n956, n51187, 
        n883, n51186, n810, n51185, n737, n51184, n664, n51183, 
        n27867, n21_adj_4521, n66088, n591, n51182, n518, n51181, 
        n445, n51180, n372_adj_4522, n51179, n299_adj_4523, n51178, 
        n226, n51177, n153, n51176, n11_adj_4524, n80;
    wire [8:0]n19645;
    
    wire n770, n51175, n697, n51174, n66069, n624, n51173, n12_adj_4525, 
        n10_adj_4526, n551, n51172, n478, n51171, n405_c, n51170, 
        n332_adj_4527, n51169, n259, n51168, n27862, n49607, n186_adj_4528, 
        n51167, n30_adj_4529, n44_adj_4530, n113, n27857;
    wire [18:0]n15384;
    
    wire n51166, n51165, n51164, n51163, n66121, n67006, n51162, 
        n1105_adj_4532, n51161, n66988, n1032_adj_4533, n51160, n959_adj_4534, 
        n51159, n886_adj_4535, n51158, n813_adj_4536, n51157, n68235, 
        n740_adj_4537, n51156, n67620, n667_adj_4538, n51155, n594_adj_4539, 
        n51154, n521_adj_4540, n51153, n68412, n16_adj_4541, n6_adj_4542, 
        n67668, n67669, n8_adj_4543, n24_adj_4544, n66030, n66024, 
        n67578, n66850, n4_adj_4546, n67664, n67665, n66059, n66057, 
        n68149, n66852, n68502, n68503, n68421, n66035, n68203, 
        n66858, n68404, n41_adj_4547, n39_adj_4548, n45_adj_4549, 
        n43_adj_4550, n29_adj_4551, n31_adj_4552, n25_adj_4553, n66485, 
        n11_adj_4555, n13_adj_4556, n15_adj_4557, n27_adj_4558, n9_adj_4559, 
        n17_adj_4560, n19_adj_4561, n21_adj_4562, n23_adj_4563, n33_adj_4564, 
        n35_adj_4565, n37_adj_4566, n66006, n65918, n12_adj_4567, 
        n448_adj_4568, n51152, n375_adj_4569, n51151, n302_adj_4570, 
        n51150, n49606, n229, n51149, n156, n51148, n14_adj_4571, 
        n83;
    wire [17:0]n16105;
    
    wire n51147, n51146, n66502, n27852, n10_adj_4572, n30_adj_4573, 
        n51145, n51144, n1108, n51143, n1035, n51142, n962, n51141, 
        n889, n51140, n816, n51139, n743, n51138, n670, n51137, 
        n597, n51136, n524, n51135, n451_adj_4574, n51134;
    wire [6:0]n20032;
    
    wire n630, n49924, n378_adj_4575, n51133, n49605, n305, n51132, 
        n232, n51131, n27847, n159, n51130, n17_adj_4576, n86;
    wire [7:0]n19825;
    
    wire n700_adj_4578, n51129, n27842, n27837, n27832, n557, n49923, 
        n627_adj_4582, n51128, n554_adj_4583, n51127, n481_adj_4584, 
        n51126, n408_adj_4585, n51125, n335_adj_4586, n51124, n262_adj_4587, 
        n51123, n484, n49922, n411, n49921, n66022, n66920, n27827, 
        n66914, n27822, n189_adj_4589, n51122, n68199, n47_adj_4590, 
        n116_adj_4591;
    wire [0:0]n11650;
    wire [21:0]n12157;
    
    wire n50187;
    wire [16:0]n16752;
    
    wire n51121, n51120, n51119, n1111, n51118, n50186, n1038, 
        n51117, n338_adj_4592, n49920, n67554, n965, n51116, n68396, 
        n892, n51115, n819, n51114, n50185, n50184, n746, n51113, 
        n265, n49919, n192_adj_4593, n49918, n50_adj_4594, n119_adj_4595, 
        n673, n51112, n16_adj_4596, n807_adj_4597, n600, n51111, 
        n50183, n527_adj_4598, n51110, n6_adj_4599, n68197, n50182;
    wire [13:0]n18065;
    
    wire n1120, n49917, n454_adj_4600, n51109, n1047, n49916, n381_adj_4601, 
        n51108, n50181, n974, n49915, n308_adj_4602, n51107, n50180, 
        n235_adj_4603, n51106, n901, n49914, n1096_adj_4604, n50179, 
        n828, n49913, n162_adj_4605, n51105, n20_adj_4606, n89_adj_4607, 
        n755, n49912;
    wire [15:0]n17329;
    
    wire n51104, n51103, n682, n49911, n1023_adj_4608, n50178, n1114_adj_4609, 
        n51102, n950_adj_4610, n50177, n68198, n877_adj_4611, n50176, 
        n804_adj_4612, n50175, n1041_adj_4613, n51101, n968_adj_4614, 
        n51100, n731_adj_4615, n50174, n49604, n658_adj_4616, n50173, 
        n585_adj_4617, n50172, n895_adj_4618, n51099, n512_adj_4619, 
        n50171, n609, n49910, n822_adj_4620, n51098, n749_adj_4621, 
        n51097, n439_adj_4622, n50170, n676_adj_4623, n51096, n603_adj_4624, 
        n51095, n530_adj_4625, n51094, n457_adj_4626, n51093, n384_adj_4627, 
        n51092, n366_adj_4628, n50169, n536, n49909, n293_adj_4629, 
        n50168, n463, n49908, n49603, n8_adj_4630, n220_adj_4631, 
        n50167, n147_adj_4632, n50166, n5_adj_4633, n74_adj_4634, 
        n311_adj_4635, n51091, n238_adj_4636, n51090, n165_adj_4637, 
        n51089, n23_adj_4638, n92_adj_4639;
    wire [6:0]n19969;
    
    wire n630_adj_4640, n51088, n557_adj_4641, n51087, n24_adj_4642, 
        n65870, n484_adj_4643, n51086, n65855, n67580, n411_adj_4644, 
        n51085, n338_adj_4645, n51084, n265_adj_4646, n51083, n192_adj_4647, 
        n51082, n50_adj_4648, n119_adj_4649;
    wire [14:0]n17840;
    
    wire n51081, n1117_adj_4650, n51080, n1044_adj_4651, n51079, n67897, 
        n971_adj_4652, n51078, n390_adj_4653, n49907, n4_adj_4654, 
        n898_adj_4655, n51077, n825_adj_4656, n51076, n752_adj_4657, 
        n51075, n679_adj_4658, n51074, n68157, n606_adj_4659, n51073, 
        n977, n68158, n1050, n533_adj_4660, n51072, n460_adj_4661, 
        n51071, n387_adj_4662, n51070, n317, n49906, n314_adj_4663, 
        n51069, n241_adj_4664, n51068, n168_adj_4665, n51067, n27817, 
        n26_adj_4667, n95_adj_4668;
    wire [13:0]n18289;
    
    wire n1120_adj_4669, n51066, n1047_adj_4670, n51065, n974_adj_4671, 
        n51064, n901_adj_4672, n51063, n828_adj_4673, n51062, n755_adj_4674, 
        n51061, n682_adj_4675, n51060, n609_adj_4676, n51059, n536_adj_4677, 
        n51058, n463_adj_4678, n51057, n390_adj_4679, n51056, n244, 
        n49905, n317_adj_4680, n51055, n244_adj_4681, n51054, n171, 
        n51053, n29_adj_4682, n98;
    wire [5:0]n20081;
    
    wire n560_adj_4683, n51052, n487_adj_4684, n51051, n65905, n414_adj_4685, 
        n51050, n65901, n68449, n67899, n68574, n68575, n68542, 
        n341_adj_4686, n51049, n268_adj_4687, n51048, n65872, n195_adj_4688, 
        n51047, n171_adj_4689, n49904, n53_c, n122_adj_4690;
    wire [12:0]n18680;
    
    wire n1050_adj_4691, n51046, n977_adj_4692, n51045, n904_adj_4693, 
        n51044, n831_adj_4694, n51043, n67902, n40_adj_4695, n68207, 
        n758, n51042, n29_adj_4696, n98_adj_4697, n685, n51041, 
        n612, n51040, n539, n51039, n466, n51038, n393_adj_4698, 
        n51037, n320, n51036, n49602, n247, n51035, n174, n51034, 
        n32_adj_4699, n101;
    wire [11:0]n19017;
    
    wire n980_adj_4700, n51033, n907_adj_4701, n51032, n834_adj_4702, 
        n51031;
    wire [20:0]n13220;
    
    wire n50148, n761_adj_4703, n51030, n688_adj_4704, n51029, n615, 
        n51028, n50147, n542, n51027, n469, n51026, n50146, n396_adj_4705, 
        n51025, n50145, n50144, n323, n51024, n250, n51023, n177, 
        n51022, n50143, n35_adj_4706, n104, n59281, n490_c, n51021, 
        n50142, n417_c, n51020, n344_adj_4707, n51019, n271_c, n51018, 
        n198_adj_4708, n51017, n56_adj_4709, n125_adj_4710;
    wire [10:0]n19304;
    
    wire n910, n51016, n837, n51015, n764, n51014, n691, n51013, 
        n618, n51012, n545, n51011, n1099_adj_4711, n50141, n472, 
        n51010, n1026_adj_4712, n50140, n399, n51009, n326, n51008, 
        n253, n51007, n953_adj_4713, n50139, n180, n51006, n107_adj_4715;
    wire [9:0]n19545;
    
    wire n840, n51005, n767_adj_4716, n51004, n694_adj_4717, n51003, 
        n621_adj_4718, n51002, n548_adj_4719, n51001, n475_adj_4720, 
        n51000, n402_adj_4721, n50999, n329_adj_4722, n50998, n256_adj_4723, 
        n50997, n183_adj_4724, n50996, n41_adj_4725, n880_adj_4727, 
        n50138, n49601;
    wire [31:0]n51;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    wire [12:0]n18485;
    
    wire n49893, n49892, n49600, n50137, n50869, n50868, n50867, 
        n50866, n50865, n50864, n50863, n50862, n50861, n50860, 
        n50859, n50858, n50857, n50856, n50855, n50854, n50853, 
        n50852, n50851, n50850, n50849, n50848, n50847, n50846, 
        n50845, n50844, n50843, n50842, n50841, n50840, n50839, 
        n49891, n49890, n50136, n758_adj_4753, n49889, n661_adj_4754, 
        n50135, n588_adj_4755, n50134, n515_adj_4756, n50133, n49743, 
        n442_adj_4757, n50132, n685_adj_4758, n49888, n369_adj_4759, 
        n50131, n49742, n612_adj_4760, n49887, n296_adj_4761, n50130, 
        n223_adj_4762, n50129, n49599, n150_adj_4763, n50128, n8_adj_4764, 
        n77_adj_4765, n49741, n539_adj_4767, n49886;
    wire [19:0]n14145;
    
    wire n50127, n466_adj_4768, n49885, n50126, n50125, n393_adj_4769, 
        n49884, n50124, n49740, n49739, n50123, n50122, n1102_adj_4772, 
        n50121, n1029_adj_4773, n50120, n956_adj_4774, n50119, n883_adj_4775, 
        n50118, n810_adj_4776, n50117, n320_adj_4777, n49883, n49738, 
        n737_adj_4779, n50116, n49598, n664_adj_4780, n50115, n591_adj_4781, 
        n50114, n49737, n518_adj_4783, n50113, n445_adj_4784, n50112, 
        n247_adj_4785, n49882, n174_adj_4786, n49881, n372_adj_4787, 
        n50111, n32_adj_4788, n101_adj_4789, n299_adj_4790, n50110, 
        n226_adj_4791, n50109, n49597, n153_adj_4792, n50108, n49736, 
        n11_adj_4794, n80_adj_4795, n49735, n49596, n49734, n49595, 
        n49733;
    wire [18:0]n14985;
    
    wire n50091, n49594;
    wire [5:0]n20129;
    
    wire n49871, n49593, n50090, n49870, n49732, n50089, n50088, 
        n49592, n50087, n49869, n50086, n49868, n49591, n50085, 
        n50084, n50083, n49590, n49731, n50082, n50081, n49867, 
        n49866, n49730, n49589, n50080, n49588;
    wire [11:0]n18849;
    
    wire n49865, n50079, n49864, n49729, n50078, n49863, n49862, 
        n49861, n49728, n50077, n49727, n50076, n49726, n615_adj_4799, 
        n49860, n542_adj_4800, n49859, n302_adj_4801, n50075, n49587, 
        n469_adj_4802, n49858, n229_adj_4803, n50074, n396_adj_4804, 
        n49857, n156_adj_4805, n50073, n49725, n323_adj_4807, n49856, 
        n250_adj_4808, n49855, n177_adj_4809, n49854, n49724, n14_adj_4811, 
        n83_adj_4812, n35_adj_4813, n104_adj_4814, n49586, n49723, 
        n49722, n49585, n49584, n49721, n49583, n910_adj_4820, n49845, 
        n837_adj_4823, n49844, n764_adj_4824, n49843, n691_adj_4825, 
        n49842;
    wire [23:0]n1_adj_4986;
    
    wire n49720, n770_adj_4827, n50057, n697_adj_4828, n50056, n49719, 
        n49582, n618_adj_4830, n49841, n624_adj_4831, n50055, n49718, 
        n545_adj_4833, n49840, n551_adj_4834, n50054, n478_adj_4835, 
        n50053, n405_adj_4836, n50052, n332_adj_4837, n50051, n259_adj_4838, 
        n50050, n472_adj_4839, n49839, n186_adj_4840, n50049, n399_adj_4841, 
        n49838, n44_adj_4842, n113_adj_4843, n326_adj_4844, n49837, 
        n50048, n49717, n50047, n253_adj_4846, n49836, n50046, n49716, 
        n50045, n49581, n1108_adj_4848, n50044, n1035_adj_4849, n50043, 
        n49715, n962_adj_4851, n50042, n180_adj_4852, n49835, n889_adj_4853, 
        n50041, n816_adj_4854, n50040, n49580, n38_adj_4855, n107_adj_4856, 
        n743_adj_4857, n50039, n670_adj_4858, n50038, n597_adj_4859, 
        n50037, n49714, n49713, n524_adj_4862, n50036, n451_adj_4863, 
        n50035, n49579, n378_adj_4864, n50034, n305_adj_4865, n50033, 
        n49712, n232_adj_4867, n50032, n49711, n159_adj_4869, n50031, 
        n17_adj_4870, n86_adj_4871, n49578, n49577, n60309, n49827;
    wire [4:0]n20200;
    
    wire n49826, n49710, n49709, n49576, n49825, n49575, n49824, 
        n49823, n49708, n49707, n49706, n49705, n49574, n49573, 
        n49704, n49703, n49702, n49627, n49701, n49572, n49700, 
        n49626, n50016, n50015, n49699, n50014, n49698, n49625, 
        n49571, n49570, n1111_adj_4896, n50013, n1038_adj_4897, n50012, 
        n37293, n25_adj_4900, n23_adj_4901, n21_adj_4902, n19_adj_4903, 
        n13_adj_4904, n15_adj_4905, n17_adj_4906, n6_adj_4907, n7_adj_4908, 
        n9_adj_4909;
    wire [1:0]n20289;
    
    wire n11_adj_4910, n5_adj_4911, n965_adj_4912, n50011, n66605, 
        n66601, n892_adj_4913, n50010, n10_adj_4914, n62242, n62244, 
        n210_adj_4915, n62248, n49454, n49697, n62252, n8_adj_4917, 
        n4_adj_4918, n12_adj_4920, n8_adj_4921, n819_adj_4923, n50009, 
        n746_adj_4924, n50008, n673_adj_4925, n50007, n6_adj_4926, 
        n16_adj_4927, n66599, n68353, n68354, n68248, n68101, n66603, 
        n68151, n66882, n68363, n600_adj_4929, n68364, n840_adj_4931, 
        n6_adj_4932, n66542;
    wire [3:0]n20249;
    wire [1:0]n20297;
    wire [2:0]n20280;
    
    wire n62200, n62202, n8_adj_4936, n6_adj_4937, n62208, n49260, 
        n60055, n60322, n4_adj_4938, n20_adj_4939, n26_adj_4940, n12_adj_4941, 
        n59546, n10_adj_4942, n9_adj_4943, n24_adj_4944, n28_adj_4945, 
        n23_adj_4946, n49388, n41_adj_4949, n39_adj_4950, n45_adj_4951, 
        n43_adj_4952, n37_adj_4953, n29_adj_4954, n31_adj_4955, n23_adj_4956, 
        n25_adj_4958, n35_adj_4959, n33_adj_4960, n9_adj_4961, n17_adj_4962, 
        n19_adj_4963, n21_adj_4964, n11_adj_4965, n13_adj_4966, n15_adj_4967, 
        n27_adj_4968, n66526, n66514, n12_adj_4969, n10_adj_4970, 
        n30_adj_4971, n67420, n67410, n68321, n67796, n68438, n67960, 
        n16_adj_4972, n8_adj_4973, n24_adj_4974, n67961, n66487, n67588, 
        n66887, n67958, n67959, n66506, n68355, n66889, n68539, 
        n68540, n68495, n66489, n68215, n66895, n68408, n68409, 
        n409, n43_adj_4976, n37_adj_4977, n39_adj_4978, n41_adj_4979, 
        n67964, n67965, n67430, n67908, n66884, n67962, n66680, 
        n67488, n69904, n49235, n12_adj_4981, n66665, n67484, n69917, 
        n16_adj_4982, n66684, n4_adj_4983, n69943, n66682, n69936, 
        n67836, n69939, n67486, n68107;
    
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_21 (.CI(n49623), .I0(n257[19]), .I1(n306[19]), .CO(n49624));
    SB_LUT4 add_6442_11_lut (.I0(GND_net), .I1(n19425[8]), .I2(n767), 
            .I3(n49810), .O(n19161[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i29_rep_79_2_lut (.I0(n356[14]), .I1(n382[14]), 
            .I2(GND_net), .I3(GND_net), .O(n69902));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i29_rep_79_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35401_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n20165[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35401_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35403_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n49338));   // verilog/motorControl.v(50[18:24])
    defparam i35403_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i52102_4_lut (.I0(n365), .I1(n69902), .I2(n382[15]), .I3(n66659), 
            .O(n67830));
    defparam i52102_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i33_rep_105_2_lut (.I0(n356[16]), .I1(n382[16]), 
            .I2(GND_net), .I3(GND_net), .O(n69928));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i33_rep_105_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52611_4_lut (.I0(n356[17]), .I1(n69928), .I2(n382[17]), .I3(n67830), 
            .O(n68339));
    defparam i52611_4_lut.LUT_INIT = 16'hffde;
    SB_DFFER result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n49[0]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n306[18]), 
            .I3(n49622), .O(n356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_23 (.CI(n49695), .I0(GND_net), .I1(n1_adj_4984[21]), 
            .CO(n49696));
    SB_LUT4 add_6239_8_lut (.I0(GND_net), .I1(n16429[5]), .I2(n527), .I3(n50005), 
            .O(n15745[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[0] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[7]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[8]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[9]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[10]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[11]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[12]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i37_rep_70_2_lut (.I0(n356[18]), .I1(n382[18]), 
            .I2(GND_net), .I3(GND_net), .O(n69893));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i37_rep_70_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52823_4_lut (.I0(n356[19]), .I1(n69893), .I2(n382[19]), .I3(n68339), 
            .O(n68551));
    defparam i52823_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i41_rep_67_2_lut (.I0(n356[20]), .I1(n382[20]), 
            .I2(GND_net), .I3(GND_net), .O(n69890));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i41_rep_67_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n356[5]), .I1(n356[9]), .I2(n19), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[19]), .I2(n20265[1]), 
            .I3(n4_adj_4449), .O(n20225[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i51006_4_lut (.I0(n11), .I1(n9), .I2(deadband[3]), .I3(n356[3]), 
            .O(n66734));
    defparam i51006_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51792_4_lut (.I0(n17_adj_4450), .I1(n15_adj_4451), .I2(n13_adj_4452), 
            .I3(n66734), .O(n67520));
    defparam i51792_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51790_4_lut (.I0(n23), .I1(n21), .I2(n19), .I3(n67520), 
            .O(n67518));
    defparam i51790_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35363_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[19]), .I2(n4_adj_4449), 
            .I3(n20265[1]), .O(n6_c));   // verilog/motorControl.v(50[18:24])
    defparam i35363_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i35355_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n20265[0]), 
            .O(n4_adj_4449));   // verilog/motorControl.v(50[18:24])
    defparam i35355_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_964 (.I0(n62), .I1(n131), .I2(n204), .I3(n20265[0]), 
            .O(n20225[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_964.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[13]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6239_8 (.CI(n50005), .I0(n16429[5]), .I1(n527), .CO(n50006));
    SB_CARRY add_6442_11 (.CI(n49810), .I0(n19425[8]), .I1(n767), .CO(n49811));
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[20]), 
            .I3(n49694), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50986_4_lut (.I0(n29), .I1(n27), .I2(n25), .I3(n67518), 
            .O(n66714));
    defparam i50986_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50248_4_lut (.I0(deadband[1]), .I1(n380), .I2(n379), .I3(deadband[0]), 
            .O(n65620));   // verilog/motorControl.v(51[12:29])
    defparam i50248_4_lut.LUT_INIT = 16'h50d4;
    SB_LUT4 add_6239_7_lut (.I0(GND_net), .I1(n16429[4]), .I2(n454), .I3(n50004), 
            .O(n15745[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i6_3_lut (.I0(n65620), .I1(n356[2]), .I2(deadband[2]), 
            .I3(GND_net), .O(n6_adj_4453));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6442_10_lut (.I0(GND_net), .I1(n19425[7]), .I2(n694), 
            .I3(n49809), .O(n19161[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_7 (.CI(n50004), .I0(n16429[4]), .I1(n454), .CO(n50005));
    SB_CARRY add_6442_10 (.CI(n49809), .I0(n19425[7]), .I1(n694), .CO(n49810));
    SB_CARRY add_18_20 (.CI(n49622), .I0(n257[18]), .I1(n306[18]), .CO(n49623));
    SB_CARRY unary_minus_13_add_3_22 (.CI(n49694), .I0(GND_net), .I1(n1_adj_4984[20]), 
            .CO(n49695));
    SB_LUT4 add_6239_6_lut (.I0(GND_net), .I1(n16429[3]), .I2(n381), .I3(n50003), 
            .O(n15745[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_6 (.CI(n50003), .I0(n16429[3]), .I1(n381), .CO(n50004));
    SB_LUT4 add_6239_5_lut (.I0(GND_net), .I1(n16429[2]), .I2(n308), .I3(n50002), 
            .O(n15745[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[19]), 
            .I3(n49693), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_9_lut (.I0(GND_net), .I1(n19425[6]), .I2(n621), .I3(n49808), 
            .O(n19161[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_5 (.CI(n50002), .I0(n16429[2]), .I1(n308), .CO(n50003));
    SB_CARRY unary_minus_13_add_3_21 (.CI(n49693), .I0(GND_net), .I1(n1_adj_4984[19]), 
            .CO(n49694));
    SB_LUT4 i52258_3_lut (.I0(n6_adj_4453), .I1(n356[14]), .I2(n29), .I3(GND_net), 
            .O(n67986));   // verilog/motorControl.v(51[12:29])
    defparam i52258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i14_3_lut (.I0(n356[8]), .I1(n356[17]), .I2(n35_c), 
            .I3(GND_net), .O(n14_adj_4455));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(23[10] 30[6])
    SB_LUT4 add_6239_4_lut (.I0(GND_net), .I1(n16429[1]), .I2(n235), .I3(n50001), 
            .O(n15745[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_9 (.CI(n49808), .I0(n19425[6]), .I1(n621), .CO(n49809));
    SB_CARRY sub_8_add_2_12 (.CI(n49568), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n49569));
    SB_CARRY add_6239_4 (.CI(n50001), .I0(n16429[1]), .I1(n235), .CO(n50002));
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n356[6]), .I1(n356[7]), .I2(n15_adj_4451), 
            .I3(GND_net), .O(n12_adj_4456));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[18]), 
            .I3(n49692), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_8_lut (.I0(GND_net), .I1(n19425[5]), .I2(n548), .I3(n49807), 
            .O(n19161[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n49692), .I0(GND_net), .I1(n1_adj_4984[18]), 
            .CO(n49693));
    SB_LUT4 LessThan_19_i32_3_lut (.I0(n14_adj_4455), .I1(n356[18]), .I2(n37), 
            .I3(GND_net), .O(n32_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6239_3_lut (.I0(GND_net), .I1(n16429[0]), .I2(n162), .I3(n50000), 
            .O(n15745[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_3 (.CI(n50000), .I0(n16429[0]), .I1(n162), .CO(n50001));
    SB_CARRY add_6442_8 (.CI(n49807), .I0(n19425[5]), .I1(n548), .CO(n49808));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n49567), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50982_4_lut (.I0(n29), .I1(n17_adj_4450), .I2(n15_adj_4451), 
            .I3(n13_adj_4452), .O(n66710));
    defparam i50982_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n306[17]), 
            .I3(n49621), .O(n356[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50841_3_lut_4_lut (.I0(PWMLimit[17]), .I1(n356[17]), .I2(n356[16]), 
            .I3(PWMLimit[16]), .O(n66569));   // verilog/motorControl.v(52[14:29])
    defparam i50841_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i34_3_lut_3_lut (.I0(PWMLimit[17]), .I1(n356[17]), 
            .I2(n356[16]), .I3(GND_net), .O(n34));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY sub_8_add_2_11 (.CI(n49567), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n49568));
    SB_LUT4 add_6442_7_lut (.I0(GND_net), .I1(n19425[4]), .I2(n475), .I3(n49806), 
            .O(n19161[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[17]), 
            .I3(n49691), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52259_3_lut (.I0(n67986), .I1(n365), .I2(n31), .I3(GND_net), 
            .O(n67987));   // verilog/motorControl.v(51[12:29])
    defparam i52259_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n49691), .I0(GND_net), .I1(n1_adj_4984[17]), 
            .CO(n49692));
    SB_LUT4 add_6239_2_lut (.I0(GND_net), .I1(n20_c), .I2(n89), .I3(GND_net), 
            .O(n15745[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n49566), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50973_4_lut (.I0(n35_c), .I1(n33), .I2(n31), .I3(n66710), 
            .O(n66701));
    defparam i50973_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[16]), 
            .I3(n49690), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_7 (.CI(n49806), .I0(n19425[4]), .I1(n475), .CO(n49807));
    SB_CARRY sub_8_add_2_10 (.CI(n49566), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n49567));
    SB_LUT4 add_6442_6_lut (.I0(GND_net), .I1(n19425[3]), .I2(n402), .I3(n49805), 
            .O(n19161[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n49621), .I0(n257[17]), .I1(n306[17]), .CO(n49622));
    SB_CARRY add_6239_2 (.CI(GND_net), .I0(n20_c), .I1(n89), .CO(n50000));
    SB_CARRY unary_minus_13_add_3_18 (.CI(n49690), .I0(GND_net), .I1(n1_adj_4984[16]), 
            .CO(n49691));
    SB_CARRY add_6442_6 (.CI(n49805), .I0(n19425[3]), .I1(n402), .CO(n49806));
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n49565), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_5_lut (.I0(GND_net), .I1(n19425[2]), .I2(n329), .I3(n49804), 
            .O(n19161[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n306[16]), 
            .I3(n49620), .O(n356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[15]), 
            .I3(n49689), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_5 (.CI(n49804), .I0(n19425[2]), .I1(n329), .CO(n49805));
    SB_LUT4 add_6442_4_lut (.I0(GND_net), .I1(n19425[1]), .I2(n256), .I3(n49803), 
            .O(n19161[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_9 (.CI(n49565), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n49566));
    SB_LUT4 i52623_4_lut (.I0(n32_c), .I1(n12_adj_4456), .I2(n37), .I3(n66696), 
            .O(n68351));   // verilog/motorControl.v(51[12:29])
    defparam i52623_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6442_4 (.CI(n49803), .I0(n19425[1]), .I1(n256), .CO(n49804));
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(n41756), 
            .I3(n49564), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51134_3_lut (.I0(n67987), .I1(n356[16]), .I2(n33), .I3(GND_net), 
            .O(n66862));   // verilog/motorControl.v(51[12:29])
    defparam i51134_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n49689), .I0(GND_net), .I1(n1_adj_4984[15]), 
            .CO(n49690));
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n382[2]), .I1(n382[3]), .I2(n356[3]), 
            .I3(GND_net), .O(n6_adj_4460));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_18_18 (.CI(n49620), .I0(n257[16]), .I1(n306[16]), .CO(n49621));
    SB_LUT4 add_6442_3_lut (.I0(GND_net), .I1(n19425[0]), .I2(n183), .I3(n49802), 
            .O(n19161[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_3 (.CI(n49802), .I0(n19425[0]), .I1(n183), .CO(n49803));
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[14]), 
            .I3(n49688), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52248_3_lut (.I0(n6_adj_4460), .I1(n382[10]), .I2(n356[10]), 
            .I3(GND_net), .O(n67976));   // verilog/motorControl.v(51[33:53])
    defparam i52248_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6442_2_lut (.I0(GND_net), .I1(n41), .I2(n110_adj_4462), 
            .I3(GND_net), .O(n19161[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_8 (.CI(n49564), .I0(setpoint[6]), .I1(n41756), 
            .CO(n49565));
    SB_CARRY add_6442_2 (.CI(GND_net), .I0(n41), .I1(n110_adj_4462), .CO(n49802));
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n306[15]), 
            .I3(n49619), .O(n365)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_16 (.CI(n49688), .I0(GND_net), .I1(n1_adj_4984[14]), 
            .CO(n49689));
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[13]), 
            .I3(n49687), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[23] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n49687), .I0(GND_net), .I1(n1_adj_4984[13]), 
            .CO(n49688));
    SB_CARRY add_18_17 (.CI(n49619), .I0(n257[15]), .I1(n306[15]), .CO(n49620));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[12]), 
            .I3(n49686), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n49686), .I0(GND_net), .I1(n1_adj_4984[12]), 
            .CO(n49687));
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n49563), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n306[14]), 
            .I3(n49618), .O(n356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n49563), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n49564));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[11]), 
            .I3(n49685), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_16 (.CI(n49618), .I0(n257[14]), .I1(n306[14]), .CO(n49619));
    SB_CARRY unary_minus_13_add_3_13 (.CI(n49685), .I0(GND_net), .I1(n1_adj_4984[11]), 
            .CO(n49686));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[10]), 
            .I3(n49684), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4470));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n49684), .I0(GND_net), .I1(n1_adj_4984[10]), 
            .CO(n49685));
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n306[13]), 
            .I3(n49617), .O(n356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_15 (.CI(n49617), .I0(n257[13]), .I1(n306[13]), .CO(n49618));
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n49562), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6491_10_lut (.I0(GND_net), .I1(n19905[7]), .I2(n700), 
            .I3(n49986), .O(n19744[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[9]), 
            .I3(n49683), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[0]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n49683), .I0(GND_net), .I1(n1_adj_4984[9]), 
            .CO(n49684));
    SB_LUT4 add_6491_9_lut (.I0(GND_net), .I1(n19905[6]), .I2(n627), .I3(n49985), 
            .O(n19744[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_6 (.CI(n49562), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n49563));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[8]), 
            .I3(n49682), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_9 (.CI(n49985), .I0(n19905[6]), .I1(n627), .CO(n49986));
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[1]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n306[12]), 
            .I3(n49616), .O(n356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6491_8_lut (.I0(GND_net), .I1(n19905[5]), .I2(n554), .I3(n49984), 
            .O(n19744[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6491_8 (.CI(n49984), .I0(n19905[5]), .I1(n554), .CO(n49985));
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6491_7_lut (.I0(GND_net), .I1(n19905[4]), .I2(n481), .I3(n49983), 
            .O(n19744[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[2]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_18_14 (.CI(n49616), .I0(n257[12]), .I1(n306[12]), .CO(n49617));
    SB_CARRY add_6491_7 (.CI(n49983), .I0(n19905[4]), .I1(n481), .CO(n49984));
    SB_CARRY unary_minus_13_add_3_10 (.CI(n49682), .I0(GND_net), .I1(n1_adj_4984[8]), 
            .CO(n49683));
    SB_LUT4 add_6491_6_lut (.I0(GND_net), .I1(n19905[3]), .I2(n408), .I3(n49982), 
            .O(n19744[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n306[11]), 
            .I3(n49615), .O(n356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(n42305), 
            .I3(n49561), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_6 (.CI(n49982), .I0(n19905[3]), .I1(n408), .CO(n49983));
    SB_LUT4 add_6491_5_lut (.I0(GND_net), .I1(n19905[2]), .I2(n335_adj_4476), 
            .I3(n49981), .O(n19744[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[7]), 
            .I3(n49681), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_5 (.CI(n49981), .I0(n19905[2]), .I1(n335_adj_4476), 
            .CO(n49982));
    SB_LUT4 add_6491_4_lut (.I0(GND_net), .I1(n19905[1]), .I2(n262), .I3(n49980), 
            .O(n19744[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_4 (.CI(n49980), .I0(n19905[1]), .I1(n262), .CO(n49981));
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[3]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52249_3_lut (.I0(n67976), .I1(n382[11]), .I2(n356[11]), .I3(GND_net), 
            .O(n67977));   // verilog/motorControl.v(51[33:53])
    defparam i52249_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_8_add_2_5 (.CI(n49561), .I0(setpoint[3]), .I1(n42305), 
            .CO(n49562));
    SB_LUT4 sub_8_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(\motor_state[2] ), 
            .I3(n49560), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_13 (.CI(n49615), .I0(n257[11]), .I1(n306[11]), .CO(n49616));
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[22] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[21] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6491_3_lut (.I0(GND_net), .I1(n19905[0]), .I2(n189_adj_4478), 
            .I3(n49979), .O(n19744[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[14]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[20] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n212));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6491_3 (.CI(n49979), .I0(n19905[0]), .I1(n189_adj_4478), 
            .CO(n49980));
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n213));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6491_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n19744[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n214));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n49681), .I0(GND_net), .I1(n1_adj_4984[7]), 
            .CO(n49682));
    SB_CARRY add_6491_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n49979));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[6]), 
            .I3(n49680), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[15]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6274_18_lut (.I0(GND_net), .I1(n17041[15]), .I2(GND_net), 
            .I3(n49978), .O(n16429[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_8 (.CI(n49680), .I0(GND_net), .I1(n1_adj_4984[6]), 
            .CO(n49681));
    SB_LUT4 add_6274_17_lut (.I0(GND_net), .I1(n17041[14]), .I2(GND_net), 
            .I3(n49977), .O(n16429[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_17 (.CI(n49977), .I0(n17041[14]), .I1(GND_net), 
            .CO(n49978));
    SB_CARRY sub_8_add_2_4 (.CI(n49560), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n49561));
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n306[10]), 
            .I3(n49614), .O(n356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6274_16_lut (.I0(GND_net), .I1(n17041[13]), .I2(n1114), 
            .I3(n49976), .O(n16429[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(\motor_state[1] ), 
            .I3(n49559), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[5]), 
            .I3(n49679), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_16 (.CI(n49976), .I0(n17041[13]), .I1(n1114), .CO(n49977));
    SB_LUT4 add_6274_15_lut (.I0(GND_net), .I1(n17041[12]), .I2(n1041), 
            .I3(n49975), .O(n16429[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52246_3_lut (.I0(n4), .I1(n382[13]), .I2(n356[13]), .I3(GND_net), 
            .O(n67974));   // verilog/motorControl.v(51[33:53])
    defparam i52246_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[4]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4485));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6274_15 (.CI(n49975), .I0(n17041[12]), .I1(n1041), .CO(n49976));
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6274_14_lut (.I0(GND_net), .I1(n17041[11]), .I2(n968), 
            .I3(n49974), .O(n16429[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29349_4_lut (.I0(PWMLimit[1]), .I1(n60589), .I2(n37308), 
            .I3(n11608), .O(n49[1]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29349_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6274_14 (.CI(n49974), .I0(n17041[11]), .I1(n968), .CO(n49975));
    SB_LUT4 add_6274_13_lut (.I0(GND_net), .I1(n17041[10]), .I2(n895), 
            .I3(n49973), .O(n16429[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_12 (.CI(n49614), .I0(n257[10]), .I1(n306[10]), .CO(n49615));
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6274_13 (.CI(n49973), .I0(n17041[10]), .I1(n895), .CO(n49974));
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6274_12_lut (.I0(GND_net), .I1(n17041[9]), .I2(n822), 
            .I3(n49972), .O(n16429[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_12 (.CI(n49972), .I0(n17041[9]), .I1(n822), .CO(n49973));
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52247_3_lut (.I0(n67974), .I1(n382[14]), .I2(n356[14]), .I3(GND_net), 
            .O(n67975));   // verilog/motorControl.v(51[33:53])
    defparam i52247_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50921_4_lut (.I0(n356[16]), .I1(n69898), .I2(n382[16]), .I3(n67476), 
            .O(n66649));
    defparam i50921_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_6274_11_lut (.I0(GND_net), .I1(n17041[8]), .I2(n749), 
            .I3(n49971), .O(n16429[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_7 (.CI(n49679), .I0(GND_net), .I1(n1_adj_4984[5]), 
            .CO(n49680));
    SB_CARRY add_6274_11 (.CI(n49971), .I0(n17041[8]), .I1(n749), .CO(n49972));
    SB_LUT4 add_6274_10_lut (.I0(GND_net), .I1(n17041[7]), .I2(n676), 
            .I3(n49970), .O(n16429[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_10 (.CI(n49970), .I0(n17041[7]), .I1(n676), .CO(n49971));
    SB_LUT4 LessThan_21_i35_rep_101_2_lut (.I0(n356[17]), .I1(n382[17]), 
            .I2(GND_net), .I3(GND_net), .O(n69924));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i35_rep_101_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6274_9_lut (.I0(GND_net), .I1(n17041[6]), .I2(n603), .I3(n49969), 
            .O(n16429[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_9 (.CI(n49969), .I0(n17041[6]), .I1(n603), .CO(n49970));
    SB_LUT4 add_6274_8_lut (.I0(GND_net), .I1(n17041[5]), .I2(n530), .I3(n49968), 
            .O(n16429[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6274_8 (.CI(n49968), .I0(n17041[5]), .I1(n530), .CO(n49969));
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6274_7_lut (.I0(GND_net), .I1(n17041[4]), .I2(n457), .I3(n49967), 
            .O(n16429[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6274_7 (.CI(n49967), .I0(n17041[4]), .I1(n457), .CO(n49968));
    SB_LUT4 i52688_4_lut (.I0(n30_c), .I1(n10_adj_4486), .I2(n69924), 
            .I3(n66637), .O(n68416));   // verilog/motorControl.v(51[33:53])
    defparam i52688_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13856_3_lut (.I0(n356[2]), .I1(n436[2]), .I2(n11610), .I3(GND_net), 
            .O(n27922));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29348_4_lut (.I0(PWMLimit[2]), .I1(n60589), .I2(n27922), 
            .I3(n11608), .O(n49[2]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29348_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6274_6_lut (.I0(GND_net), .I1(n17041[3]), .I2(n384), .I3(n49966), 
            .O(n16429[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_6 (.CI(n49966), .I0(n17041[3]), .I1(n384), .CO(n49967));
    SB_LUT4 add_6274_5_lut (.I0(GND_net), .I1(n17041[2]), .I2(n311), .I3(n49965), 
            .O(n16429[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_5 (.CI(n49965), .I0(n17041[2]), .I1(n311), .CO(n49966));
    SB_LUT4 add_6274_4_lut (.I0(GND_net), .I1(n17041[1]), .I2(n238), .I3(n49964), 
            .O(n16429[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_4 (.CI(n49964), .I0(n17041[1]), .I1(n238), .CO(n49965));
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51144_3_lut (.I0(n67975), .I1(n382[15]), .I2(n365), .I3(GND_net), 
            .O(n66872));   // verilog/motorControl.v(51[33:53])
    defparam i51144_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6274_3_lut (.I0(GND_net), .I1(n17041[0]), .I2(n165), .I3(n49963), 
            .O(n16429[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6274_3 (.CI(n49963), .I0(n17041[0]), .I1(n165), .CO(n49964));
    SB_LUT4 add_6274_2_lut (.I0(GND_net), .I1(n23_adj_4485), .I2(n92), 
            .I3(GND_net), .O(n16429[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6274_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[4]), 
            .I3(n49678), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13851_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n11610), .I3(GND_net), 
            .O(n27917));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13851_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6274_2 (.CI(GND_net), .I0(n23_adj_4485), .I1(n92), .CO(n49963));
    SB_LUT4 i29347_4_lut (.I0(PWMLimit[3]), .I1(n60589), .I2(n27917), 
            .I3(n11608), .O(n49[3]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29347_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13846_3_lut (.I0(n356[4]), .I1(n436[4]), .I2(n11610), .I3(GND_net), 
            .O(n27912));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52809_4_lut (.I0(n66872), .I1(n68416), .I2(n69924), .I3(n66649), 
            .O(n68537));   // verilog/motorControl.v(51[33:53])
    defparam i52809_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29346_4_lut (.I0(PWMLimit[4]), .I1(n60589), .I2(n27912), 
            .I3(n11608), .O(n49[4]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29346_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[5]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[6]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52810_3_lut (.I0(n68537), .I1(n382[18]), .I2(n356[18]), .I3(GND_net), 
            .O(n68538));   // verilog/motorControl.v(51[33:53])
    defparam i52810_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52771_3_lut (.I0(n68538), .I1(n382[19]), .I2(n356[19]), .I3(GND_net), 
            .O(n68499));   // verilog/motorControl.v(51[33:53])
    defparam i52771_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50885_4_lut (.I0(n356[21]), .I1(n69912), .I2(n382[21]), .I3(n67482), 
            .O(n66613));
    defparam i50885_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[15] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4478));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51856_4_lut (.I0(n24_adj_4488), .I1(n8_adj_4489), .I2(n69888), 
            .I3(n66611), .O(n67584));   // verilog/motorControl.v(51[33:53])
    defparam i51856_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n306[9]), .I3(n49613), 
            .O(n356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[7]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4476));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51142_3_lut (.I0(n67977), .I1(n382[12]), .I2(n356[12]), .I3(GND_net), 
            .O(n66870));   // verilog/motorControl.v(51[33:53])
    defparam i51142_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_13_add_3_6 (.CI(n49678), .I0(GND_net), .I1(n1_adj_4984[4]), 
            .CO(n49679));
    SB_LUT4 i50887_4_lut (.I0(n356[21]), .I1(n69890), .I2(n382[21]), .I3(n68551), 
            .O(n66615));
    defparam i50887_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_18_11 (.CI(n49613), .I0(n257[9]), .I1(n306[9]), .CO(n49614));
    SB_LUT4 LessThan_21_i45_rep_65_2_lut (.I0(n356[22]), .I1(n382[22]), 
            .I2(GND_net), .I3(GND_net), .O(n69888));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i45_rep_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52483_4_lut (.I0(n66870), .I1(n67584), .I2(n69888), .I3(n66613), 
            .O(n68211));   // verilog/motorControl.v(51[33:53])
    defparam i52483_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13841_3_lut (.I0(n356[5]), .I1(n436[5]), .I2(n11610), .I3(GND_net), 
            .O(n27907));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29345_4_lut (.I0(PWMLimit[5]), .I1(n60589), .I2(n27907), 
            .I3(n11608), .O(n49[5]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29345_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i51150_3_lut (.I0(n68499), .I1(n382[20]), .I2(n356[20]), .I3(GND_net), 
            .O(n66878));   // verilog/motorControl.v(51[33:53])
    defparam i51150_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13836_3_lut (.I0(n356[6]), .I1(n436[6]), .I2(n11610), .I3(GND_net), 
            .O(n27902));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29344_4_lut (.I0(PWMLimit[6]), .I1(n60589), .I2(n27902), 
            .I3(n11608), .O(n49[6]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29344_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[3]), 
            .I3(n49677), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n306[8]), .I3(n49612), 
            .O(n356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_10 (.CI(n49612), .I0(n257[8]), .I1(n306[8]), .CO(n49613));
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[8]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_13_add_3_5 (.CI(n49677), .I0(GND_net), .I1(n1_adj_4984[3]), 
            .CO(n49678));
    SB_CARRY sub_8_add_2_3 (.CI(n49559), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n49560));
    SB_LUT4 sub_8_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(\motor_state[0] ), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13831_3_lut (.I0(n356[7]), .I1(n436[7]), .I2(n11610), .I3(GND_net), 
            .O(n27897));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n306[7]), .I3(n49611), 
            .O(n356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29343_4_lut (.I0(PWMLimit[7]), .I1(n60589), .I2(n27897), 
            .I3(n11608), .O(n49[7]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29343_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[2]), 
            .I3(n49676), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n49559));
    SB_LUT4 i13826_3_lut (.I0(n356[8]), .I1(n436[8]), .I2(n11610), .I3(GND_net), 
            .O(n27892));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29342_4_lut (.I0(PWMLimit[8]), .I1(n60589), .I2(n27892), 
            .I3(n11608), .O(n49[8]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29342_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13821_3_lut (.I0(n356[9]), .I1(n436[9]), .I2(n11610), .I3(GND_net), 
            .O(n27887));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_9 (.CI(n49611), .I0(n257[7]), .I1(n306[7]), .CO(n49612));
    SB_LUT4 i29341_4_lut (.I0(PWMLimit[9]), .I1(n60589), .I2(n27887), 
            .I3(n11608), .O(n49[9]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29341_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6307_17_lut (.I0(GND_net), .I1(n17585[14]), .I2(GND_net), 
            .I3(n49950), .O(n17041[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n306[6]), .I3(n49610), 
            .O(n356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_16_lut (.I0(GND_net), .I1(n17585[13]), .I2(n1117), 
            .I3(n49949), .O(n17041[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_16 (.CI(n49949), .I0(n17585[13]), .I1(n1117), .CO(n49950));
    SB_CARRY unary_minus_13_add_3_4 (.CI(n49676), .I0(GND_net), .I1(n1_adj_4984[2]), 
            .CO(n49677));
    SB_LUT4 add_6307_15_lut (.I0(GND_net), .I1(n17585[12]), .I2(n1044), 
            .I3(n49948), .O(n17041[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_15 (.CI(n49948), .I0(n17585[12]), .I1(n1044), .CO(n49949));
    SB_LUT4 add_6307_14_lut (.I0(GND_net), .I1(n17585[11]), .I2(n971), 
            .I3(n49947), .O(n17041[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[1]), 
            .I3(n49675), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_14 (.CI(n49947), .I0(n17585[11]), .I1(n971), .CO(n49948));
    SB_LUT4 add_6307_13_lut (.I0(GND_net), .I1(n17585[10]), .I2(n898), 
            .I3(n49946), .O(n17041[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_3 (.CI(n49675), .I0(GND_net), .I1(n1_adj_4984[1]), 
            .CO(n49676));
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_13 (.CI(n49946), .I0(n17585[10]), .I1(n898), .CO(n49947));
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[9]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4494));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6307_12_lut (.I0(GND_net), .I1(n17585[9]), .I2(n825), 
            .I3(n49945), .O(n17041[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4984[0]), 
            .CO(n49675));
    SB_CARRY add_6307_12 (.CI(n49945), .I0(n17585[9]), .I1(n825), .CO(n49946));
    SB_LUT4 add_6307_11_lut (.I0(GND_net), .I1(n17585[8]), .I2(n752), 
            .I3(n49944), .O(n17041[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_11 (.CI(n49944), .I0(n17585[8]), .I1(n752), .CO(n49945));
    SB_CARRY add_18_8 (.CI(n49610), .I0(n257[6]), .I1(n306[6]), .CO(n49611));
    SB_LUT4 add_6307_10_lut (.I0(GND_net), .I1(n17585[7]), .I2(n679), 
            .I3(n49943), .O(n17041[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6307_10 (.CI(n49943), .I0(n17585[7]), .I1(n679), .CO(n49944));
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4495));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6307_9_lut (.I0(GND_net), .I1(n17585[6]), .I2(n606), .I3(n49942), 
            .O(n17041[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4496));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6307_9 (.CI(n49942), .I0(n17585[6]), .I1(n606), .CO(n49943));
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n356[3]), .I1(n356[4]), .I2(n9), 
            .I3(GND_net), .O(n8_adj_4497));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52262_3_lut (.I0(n8_adj_4497), .I1(n356[11]), .I2(n23), .I3(GND_net), 
            .O(n67990));   // verilog/motorControl.v(51[12:29])
    defparam i52262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52263_3_lut (.I0(n67990), .I1(n356[12]), .I2(n25), .I3(GND_net), 
            .O(n67991));   // verilog/motorControl.v(51[12:29])
    defparam i52263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50992_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n65796), 
            .O(n66720));
    defparam i50992_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51854_3_lut (.I0(n10), .I1(n356[10]), .I2(n21), .I3(GND_net), 
            .O(n67582));   // verilog/motorControl.v(51[12:29])
    defparam i51854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51132_3_lut (.I0(n67991), .I1(n356[13]), .I2(n27), .I3(GND_net), 
            .O(n66860));   // verilog/motorControl.v(51[12:29])
    defparam i51132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52387_4_lut (.I0(n35_c), .I1(n33), .I2(n31), .I3(n66714), 
            .O(n68115));
    defparam i52387_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52807_4_lut (.I0(n66862), .I1(n68351), .I2(n37), .I3(n66701), 
            .O(n68535));   // verilog/motorControl.v(51[12:29])
    defparam i52807_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52425_4_lut (.I0(n66860), .I1(n67582), .I2(n27), .I3(n66720), 
            .O(n68153));   // verilog/motorControl.v(51[12:29])
    defparam i52425_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52868_4_lut (.I0(n68153), .I1(n68535), .I2(n37), .I3(n68115), 
            .O(n68596));   // verilog/motorControl.v(51[12:29])
    defparam i52868_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52869_3_lut (.I0(n68596), .I1(n356[19]), .I2(deadband[19]), 
            .I3(GND_net), .O(n68597));   // verilog/motorControl.v(51[12:29])
    defparam i52869_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52723_3_lut (.I0(n68597), .I1(n356[20]), .I2(deadband[20]), 
            .I3(GND_net), .O(n68451));   // verilog/motorControl.v(51[12:29])
    defparam i52723_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52637_3_lut (.I0(n68451), .I1(n356[21]), .I2(deadband[21]), 
            .I3(GND_net), .O(n68365));   // verilog/motorControl.v(51[12:29])
    defparam i52637_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52638_3_lut (.I0(n68365), .I1(n356[22]), .I2(deadband[22]), 
            .I3(GND_net), .O(n68366));   // verilog/motorControl.v(51[12:29])
    defparam i52638_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52678_4_lut (.I0(n66878), .I1(n68211), .I2(n69888), .I3(n66615), 
            .O(n68406));   // verilog/motorControl.v(51[33:53])
    defparam i52678_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut (.I0(n68366), .I1(control_update), .I2(deadband[23]), 
            .I3(n356[23]), .O(n62222));
    defparam i1_4_lut.LUT_INIT = 16'h4c04;
    SB_LUT4 i1_4_lut_adj_965 (.I0(n62222), .I1(n68406), .I2(n356[23]), 
            .I3(n47_adj_4498), .O(n60589));
    defparam i1_4_lut_adj_965.LUT_INIT = 16'h0a22;
    SB_LUT4 add_6307_8_lut (.I0(GND_net), .I1(n17585[5]), .I2(n533), .I3(n49941), 
            .O(n17041[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_8 (.CI(n49941), .I0(n17585[5]), .I1(n533), .CO(n49942));
    SB_LUT4 add_6307_7_lut (.I0(GND_net), .I1(n17585[4]), .I2(n460_c), 
            .I3(n49940), .O(n17041[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n306[5]), .I3(n49609), 
            .O(n356[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_7 (.CI(n49940), .I0(n17585[4]), .I1(n460_c), .CO(n49941));
    SB_LUT4 add_6307_6_lut (.I0(GND_net), .I1(n17585[3]), .I2(n387_adj_4470), 
            .I3(n49939), .O(n17041[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_6 (.CI(n49939), .I0(n17585[3]), .I1(n387_adj_4470), 
            .CO(n49940));
    SB_LUT4 i5967_2_lut_4_lut (.I0(control_update), .I1(n67963), .I2(PWMLimit[23]), 
            .I3(n356[23]), .O(n11608));
    defparam i5967_2_lut_4_lut.LUT_INIT = 16'h2a02;
    SB_LUT4 add_6307_5_lut (.I0(GND_net), .I1(n17585[2]), .I2(n314), .I3(n49938), 
            .O(n17041[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_5 (.CI(n49938), .I0(n17585[2]), .I1(n314), .CO(n49939));
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4499));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_c));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4500));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4501));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4502));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4503));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4504));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6307_4_lut (.I0(GND_net), .I1(n17585[1]), .I2(n241), .I3(n49937), 
            .O(n17041[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_4 (.CI(n49937), .I0(n17585[1]), .I1(n241), .CO(n49938));
    SB_LUT4 add_6307_3_lut (.I0(GND_net), .I1(n17585[0]), .I2(n168), .I3(n49936), 
            .O(n17041[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13816_3_lut (.I0(n356[10]), .I1(n436[10]), .I2(n11610), .I3(GND_net), 
            .O(n27882));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13816_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6307_3 (.CI(n49936), .I0(n17585[0]), .I1(n168), .CO(n49937));
    SB_LUT4 i29340_4_lut (.I0(PWMLimit[10]), .I1(n60589), .I2(n27882), 
            .I3(n11608), .O(n49[10]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29340_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3715[23] ), 
            .I1(n12736[21]), .I2(GND_net), .I3(n51238), .O(n12229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n12736[20]), .I2(GND_net), 
            .I3(n51237), .O(n306[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_23 (.CI(n51237), .I0(n12736[20]), .I1(GND_net), 
            .CO(n51238));
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n12736[19]), .I2(GND_net), 
            .I3(n51236), .O(n306[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_22 (.CI(n51236), .I0(n12736[19]), .I1(GND_net), 
            .CO(n51237));
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n12736[18]), .I2(GND_net), 
            .I3(n51235), .O(n306[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n17041[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_21 (.CI(n51235), .I0(n12736[18]), .I1(GND_net), 
            .CO(n51236));
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n12736[17]), .I2(GND_net), 
            .I3(n51234), .O(n306[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n49936));
    SB_CARRY mult_17_add_1225_20 (.CI(n51234), .I0(n12736[17]), .I1(GND_net), 
            .CO(n51235));
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n12736[16]), .I2(GND_net), 
            .I3(n51233), .O(n306[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n51233), .I0(n12736[16]), .I1(GND_net), 
            .CO(n51234));
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n12736[15]), .I2(GND_net), 
            .I3(n51232), .O(n306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n51232), .I0(n12736[15]), .I1(GND_net), 
            .CO(n51233));
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n12736[14]), .I2(GND_net), 
            .I3(n51231), .O(n306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_17 (.CI(n51231), .I0(n12736[14]), .I1(GND_net), 
            .CO(n51232));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n12736[13]), .I2(n1096), 
            .I3(n51230), .O(n306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13811_3_lut (.I0(n356[11]), .I1(n436[11]), .I2(n11610), .I3(GND_net), 
            .O(n27877));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13811_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_17_add_1225_16 (.CI(n51230), .I0(n12736[13]), .I1(n1096), 
            .CO(n51231));
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n12736[12]), .I2(n1023), 
            .I3(n51229), .O(n306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29339_4_lut (.I0(PWMLimit[11]), .I1(n60589), .I2(n27877), 
            .I3(n11608), .O(n49[11]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29339_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY mult_17_add_1225_15 (.CI(n51229), .I0(n12736[12]), .I1(n1023), 
            .CO(n51230));
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n12736[11]), .I2(n950), 
            .I3(n51228), .O(n306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_14 (.CI(n51228), .I0(n12736[11]), .I1(n950), 
            .CO(n51229));
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n12736[10]), .I2(n877), 
            .I3(n51227), .O(n306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_13 (.CI(n51227), .I0(n12736[10]), .I1(n877), 
            .CO(n51228));
    SB_CARRY add_18_7 (.CI(n49609), .I0(n257[5]), .I1(n306[5]), .CO(n49610));
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n306[4]), .I3(n49608), 
            .O(n356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n12736[9]), .I2(n804), 
            .I3(n51226), .O(n306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_12 (.CI(n51226), .I0(n12736[9]), .I1(n804), 
            .CO(n51227));
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n12736[8]), .I2(n731), 
            .I3(n51225), .O(n306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_11 (.CI(n51225), .I0(n12736[8]), .I1(n731), 
            .CO(n51226));
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n12736[7]), .I2(n658), 
            .I3(n51224), .O(n306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_10 (.CI(n51224), .I0(n12736[7]), .I1(n658), 
            .CO(n51225));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n12736[6]), .I2(n585), 
            .I3(n51223), .O(n306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_9 (.CI(n51223), .I0(n12736[6]), .I1(n585), 
            .CO(n51224));
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n12736[5]), .I2(n512), 
            .I3(n51222), .O(n306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_8 (.CI(n51222), .I0(n12736[5]), .I1(n512), 
            .CO(n51223));
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n12736[4]), .I2(n439), 
            .I3(n51221), .O(n306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_7 (.CI(n51221), .I0(n12736[4]), .I1(n439), 
            .CO(n51222));
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n12736[3]), .I2(n366_adj_4505), 
            .I3(n51220), .O(n306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_6 (.CI(n51220), .I0(n12736[3]), .I1(n366_adj_4505), 
            .CO(n51221));
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n12736[2]), .I2(n293_adj_4506), 
            .I3(n51219), .O(n306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_5 (.CI(n51219), .I0(n12736[2]), .I1(n293_adj_4506), 
            .CO(n51220));
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n12736[1]), .I2(n220), 
            .I3(n51218), .O(n306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13806_3_lut (.I0(n356[12]), .I1(n436[12]), .I2(n11610), .I3(GND_net), 
            .O(n27872));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13806_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_17_add_1225_4 (.CI(n51218), .I0(n12736[1]), .I1(n220), 
            .CO(n51219));
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n12736[0]), .I2(n147), 
            .I3(n51217), .O(n306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_3 (.CI(n51217), .I0(n12736[0]), .I1(n147), 
            .CO(n51218));
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4508), .I2(n74), 
            .I3(GND_net), .O(n306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5_adj_4508), .I1(n74), 
            .CO(n51217));
    SB_LUT4 add_6100_23_lut (.I0(GND_net), .I1(n13704[20]), .I2(GND_net), 
            .I3(n51216), .O(n12736[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6100_22_lut (.I0(GND_net), .I1(n13704[19]), .I2(GND_net), 
            .I3(n51215), .O(n12736[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_22 (.CI(n51215), .I0(n13704[19]), .I1(GND_net), 
            .CO(n51216));
    SB_LUT4 add_6100_21_lut (.I0(GND_net), .I1(n13704[18]), .I2(GND_net), 
            .I3(n51214), .O(n12736[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_21 (.CI(n51214), .I0(n13704[18]), .I1(GND_net), 
            .CO(n51215));
    SB_LUT4 add_6100_20_lut (.I0(GND_net), .I1(n13704[17]), .I2(GND_net), 
            .I3(n51213), .O(n12736[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_20 (.CI(n51213), .I0(n13704[17]), .I1(GND_net), 
            .CO(n51214));
    SB_LUT4 add_6100_19_lut (.I0(GND_net), .I1(n13704[16]), .I2(GND_net), 
            .I3(n51212), .O(n12736[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29338_4_lut (.I0(PWMLimit[12]), .I1(n60589), .I2(n27872), 
            .I3(n11608), .O(n49[12]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29338_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6100_19 (.CI(n51212), .I0(n13704[16]), .I1(GND_net), 
            .CO(n51213));
    SB_LUT4 add_6100_18_lut (.I0(GND_net), .I1(n13704[15]), .I2(GND_net), 
            .I3(n51211), .O(n12736[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_18 (.CI(n51211), .I0(n13704[15]), .I1(GND_net), 
            .CO(n51212));
    SB_LUT4 add_6100_17_lut (.I0(GND_net), .I1(n13704[14]), .I2(GND_net), 
            .I3(n51210), .O(n12736[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4509));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6100_17 (.CI(n51210), .I0(n13704[14]), .I1(GND_net), 
            .CO(n51211));
    SB_LUT4 add_6100_16_lut (.I0(GND_net), .I1(n13704[13]), .I2(n1099), 
            .I3(n51209), .O(n12736[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4511));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6100_16 (.CI(n51209), .I0(n13704[13]), .I1(n1099), .CO(n51210));
    SB_LUT4 add_6100_15_lut (.I0(GND_net), .I1(n13704[12]), .I2(n1026), 
            .I3(n51208), .O(n12736[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_15 (.CI(n51208), .I0(n13704[12]), .I1(n1026), .CO(n51209));
    SB_LUT4 add_6100_14_lut (.I0(GND_net), .I1(n13704[11]), .I2(n953), 
            .I3(n51207), .O(n12736[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_14 (.CI(n51207), .I0(n13704[11]), .I1(n953), .CO(n51208));
    SB_LUT4 add_6100_13_lut (.I0(GND_net), .I1(n13704[10]), .I2(n880), 
            .I3(n51206), .O(n12736[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_13 (.CI(n51206), .I0(n13704[10]), .I1(n880), .CO(n51207));
    SB_LUT4 add_6100_12_lut (.I0(GND_net), .I1(n13704[9]), .I2(n807), 
            .I3(n51205), .O(n12736[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_12 (.CI(n51205), .I0(n13704[9]), .I1(n807), .CO(n51206));
    SB_LUT4 add_6100_11_lut (.I0(GND_net), .I1(n13704[8]), .I2(n734_adj_4512), 
            .I3(n51204), .O(n12736[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_11 (.CI(n51204), .I0(n13704[8]), .I1(n734_adj_4512), 
            .CO(n51205));
    SB_LUT4 add_6100_10_lut (.I0(GND_net), .I1(n13704[7]), .I2(n661), 
            .I3(n51203), .O(n12736[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_10 (.CI(n51203), .I0(n13704[7]), .I1(n661), .CO(n51204));
    SB_LUT4 add_6100_9_lut (.I0(GND_net), .I1(n13704[6]), .I2(n588), .I3(n51202), 
            .O(n12736[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_9 (.CI(n51202), .I0(n13704[6]), .I1(n588), .CO(n51203));
    SB_LUT4 add_6100_8_lut (.I0(GND_net), .I1(n13704[5]), .I2(n515), .I3(n51201), 
            .O(n12736[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_8 (.CI(n51201), .I0(n13704[5]), .I1(n515), .CO(n51202));
    SB_LUT4 add_6100_7_lut (.I0(GND_net), .I1(n13704[4]), .I2(n442), .I3(n51200), 
            .O(n12736[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4513));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6100_7 (.CI(n51200), .I0(n13704[4]), .I1(n442), .CO(n51201));
    SB_LUT4 add_6100_6_lut (.I0(GND_net), .I1(n13704[3]), .I2(n369_adj_4514), 
            .I3(n51199), .O(n12736[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_6 (.CI(n51199), .I0(n13704[3]), .I1(n369_adj_4514), 
            .CO(n51200));
    SB_LUT4 add_6100_5_lut (.I0(GND_net), .I1(n13704[2]), .I2(n296_adj_4515), 
            .I3(n51198), .O(n12736[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_5 (.CI(n51198), .I0(n13704[2]), .I1(n296_adj_4515), 
            .CO(n51199));
    SB_LUT4 add_6100_4_lut (.I0(GND_net), .I1(n13704[1]), .I2(n223), .I3(n51197), 
            .O(n12736[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_4 (.CI(n51197), .I0(n13704[1]), .I1(n223), .CO(n51198));
    SB_LUT4 add_6100_3_lut (.I0(GND_net), .I1(n13704[0]), .I2(n150), .I3(n51196), 
            .O(n12736[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_3 (.CI(n51196), .I0(n13704[0]), .I1(n150), .CO(n51197));
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4517));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6100_2_lut (.I0(GND_net), .I1(n8_adj_4518), .I2(n77), 
            .I3(GND_net), .O(n12736[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_2 (.CI(GND_net), .I0(n8_adj_4518), .I1(n77), .CO(n51196));
    SB_LUT4 add_6143_22_lut (.I0(GND_net), .I1(n14585[19]), .I2(GND_net), 
            .I3(n51195), .O(n13704[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6143_21_lut (.I0(GND_net), .I1(n14585[18]), .I2(GND_net), 
            .I3(n51194), .O(n13704[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_21 (.CI(n51194), .I0(n14585[18]), .I1(GND_net), 
            .CO(n51195));
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4519));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6143_20_lut (.I0(GND_net), .I1(n14585[17]), .I2(GND_net), 
            .I3(n51193), .O(n13704[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_20 (.CI(n51193), .I0(n14585[17]), .I1(GND_net), 
            .CO(n51194));
    SB_LUT4 add_6143_19_lut (.I0(GND_net), .I1(n14585[16]), .I2(GND_net), 
            .I3(n51192), .O(n13704[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_19 (.CI(n51192), .I0(n14585[16]), .I1(GND_net), 
            .CO(n51193));
    SB_LUT4 add_6143_18_lut (.I0(GND_net), .I1(n14585[15]), .I2(GND_net), 
            .I3(n51191), .O(n13704[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_18 (.CI(n51191), .I0(n14585[15]), .I1(GND_net), 
            .CO(n51192));
    SB_LUT4 add_6143_17_lut (.I0(GND_net), .I1(n14585[14]), .I2(GND_net), 
            .I3(n51190), .O(n13704[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_17 (.CI(n51190), .I0(n14585[14]), .I1(GND_net), 
            .CO(n51191));
    SB_LUT4 add_6143_16_lut (.I0(GND_net), .I1(n14585[13]), .I2(n1102), 
            .I3(n51189), .O(n13704[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_16 (.CI(n51189), .I0(n14585[13]), .I1(n1102), .CO(n51190));
    SB_LUT4 add_6143_15_lut (.I0(GND_net), .I1(n14585[12]), .I2(n1029), 
            .I3(n51188), .O(n13704[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4520));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6143_15 (.CI(n51188), .I0(n14585[12]), .I1(n1029), .CO(n51189));
    SB_LUT4 add_6143_14_lut (.I0(GND_net), .I1(n14585[11]), .I2(n956), 
            .I3(n51187), .O(n13704[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_14 (.CI(n51187), .I0(n14585[11]), .I1(n956), .CO(n51188));
    SB_LUT4 add_6143_13_lut (.I0(GND_net), .I1(n14585[10]), .I2(n883), 
            .I3(n51186), .O(n13704[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_13 (.CI(n51186), .I0(n14585[10]), .I1(n883), .CO(n51187));
    SB_LUT4 add_6143_12_lut (.I0(GND_net), .I1(n14585[9]), .I2(n810), 
            .I3(n51185), .O(n13704[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_12 (.CI(n51185), .I0(n14585[9]), .I1(n810), .CO(n51186));
    SB_LUT4 add_6143_11_lut (.I0(GND_net), .I1(n14585[8]), .I2(n737), 
            .I3(n51184), .O(n13704[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_11 (.CI(n51184), .I0(n14585[8]), .I1(n737), .CO(n51185));
    SB_LUT4 add_6143_10_lut (.I0(GND_net), .I1(n14585[7]), .I2(n664), 
            .I3(n51183), .O(n13704[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13801_3_lut (.I0(n356[13]), .I1(n436[13]), .I2(n11610), .I3(GND_net), 
            .O(n27867));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4521));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50360_4_lut (.I0(n21_adj_4521), .I1(n19_adj_4520), .I2(n17_adj_4519), 
            .I3(n9_adj_4517), .O(n66088));
    defparam i50360_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6143_10 (.CI(n51183), .I0(n14585[7]), .I1(n664), .CO(n51184));
    SB_CARRY add_18_6 (.CI(n49608), .I0(n257[4]), .I1(n306[4]), .CO(n49609));
    SB_LUT4 add_6143_9_lut (.I0(GND_net), .I1(n14585[6]), .I2(n591), .I3(n51182), 
            .O(n13704[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_9 (.CI(n51182), .I0(n14585[6]), .I1(n591), .CO(n51183));
    SB_LUT4 add_6143_8_lut (.I0(GND_net), .I1(n14585[5]), .I2(n518), .I3(n51181), 
            .O(n13704[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_8 (.CI(n51181), .I0(n14585[5]), .I1(n518), .CO(n51182));
    SB_LUT4 add_6143_7_lut (.I0(GND_net), .I1(n14585[4]), .I2(n445), .I3(n51180), 
            .O(n13704[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_7 (.CI(n51180), .I0(n14585[4]), .I1(n445), .CO(n51181));
    SB_LUT4 add_6143_6_lut (.I0(GND_net), .I1(n14585[3]), .I2(n372_adj_4522), 
            .I3(n51179), .O(n13704[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_6 (.CI(n51179), .I0(n14585[3]), .I1(n372_adj_4522), 
            .CO(n51180));
    SB_LUT4 i29337_4_lut (.I0(PWMLimit[13]), .I1(n60589), .I2(n27867), 
            .I3(n11608), .O(n49[13]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29337_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6143_5_lut (.I0(GND_net), .I1(n14585[2]), .I2(n299_adj_4523), 
            .I3(n51178), .O(n13704[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_5 (.CI(n51178), .I0(n14585[2]), .I1(n299_adj_4523), 
            .CO(n51179));
    SB_LUT4 add_6143_4_lut (.I0(GND_net), .I1(n14585[1]), .I2(n226), .I3(n51177), 
            .O(n13704[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_4 (.CI(n51177), .I0(n14585[1]), .I1(n226), .CO(n51178));
    SB_LUT4 add_6143_3_lut (.I0(GND_net), .I1(n14585[0]), .I2(n153), .I3(n51176), 
            .O(n13704[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_3 (.CI(n51176), .I0(n14585[0]), .I1(n153), .CO(n51177));
    SB_LUT4 add_6143_2_lut (.I0(GND_net), .I1(n11_adj_4524), .I2(n80), 
            .I3(GND_net), .O(n13704[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_2 (.CI(GND_net), .I0(n11_adj_4524), .I1(n80), .CO(n51176));
    SB_LUT4 add_6463_11_lut (.I0(GND_net), .I1(n19645[8]), .I2(n770), 
            .I3(n51175), .O(n19425[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6463_10_lut (.I0(GND_net), .I1(n19645[7]), .I2(n697), 
            .I3(n51174), .O(n19425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_10 (.CI(n51174), .I0(n19645[7]), .I1(n697), .CO(n51175));
    SB_LUT4 i50341_4_lut (.I0(n27_adj_4513), .I1(n15_adj_4511), .I2(n13_adj_4509), 
            .I3(n11_adj_4504), .O(n66069));
    defparam i50341_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6463_9_lut (.I0(GND_net), .I1(n19645[6]), .I2(n624), .I3(n51173), 
            .O(n19425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_4503), 
            .I3(GND_net), .O(n12_adj_4525));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6463_9 (.CI(n51173), .I0(n19645[6]), .I1(n624), .CO(n51174));
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_4509), 
            .I3(GND_net), .O(n10_adj_4526));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6463_8_lut (.I0(GND_net), .I1(n19645[5]), .I2(n551), .I3(n51172), 
            .O(n19425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_8 (.CI(n51172), .I0(n19645[5]), .I1(n551), .CO(n51173));
    SB_LUT4 add_6463_7_lut (.I0(GND_net), .I1(n19645[4]), .I2(n478), .I3(n51171), 
            .O(n19425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_7 (.CI(n51171), .I0(n19645[4]), .I1(n478), .CO(n51172));
    SB_LUT4 add_6463_6_lut (.I0(GND_net), .I1(n19645[3]), .I2(n405_c), 
            .I3(n51170), .O(n19425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_6 (.CI(n51170), .I0(n19645[3]), .I1(n405_c), .CO(n51171));
    SB_LUT4 add_6463_5_lut (.I0(GND_net), .I1(n19645[2]), .I2(n332_adj_4527), 
            .I3(n51169), .O(n19425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_5 (.CI(n51169), .I0(n19645[2]), .I1(n332_adj_4527), 
            .CO(n51170));
    SB_LUT4 add_6463_4_lut (.I0(GND_net), .I1(n19645[1]), .I2(n259), .I3(n51168), 
            .O(n19425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13796_3_lut (.I0(n356[14]), .I1(n436[14]), .I2(n11610), .I3(GND_net), 
            .O(n27862));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13796_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6463_4 (.CI(n51168), .I0(n19645[1]), .I1(n259), .CO(n51169));
    SB_LUT4 i29336_4_lut (.I0(PWMLimit[14]), .I1(n60589), .I2(n27862), 
            .I3(n11608), .O(n49[14]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29336_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n306[3]), .I3(n49607), 
            .O(n356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6463_3_lut (.I0(GND_net), .I1(n19645[0]), .I2(n186_adj_4528), 
            .I3(n51167), .O(n19425[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_3 (.CI(n51167), .I0(n19645[0]), .I1(n186_adj_4528), 
            .CO(n51168));
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_4525), .I1(n130[17]), .I2(n35_adj_4502), 
            .I3(GND_net), .O(n30_adj_4529));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6463_2_lut (.I0(GND_net), .I1(n44_adj_4530), .I2(n113), 
            .I3(GND_net), .O(n19425[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6463_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6463_2 (.CI(GND_net), .I0(n44_adj_4530), .I1(n113), .CO(n51167));
    SB_LUT4 i13791_3_lut (.I0(n365), .I1(n436[15]), .I2(n11610), .I3(GND_net), 
            .O(n27857));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6183_21_lut (.I0(GND_net), .I1(n15384[18]), .I2(GND_net), 
            .I3(n51166), .O(n14585[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6183_20_lut (.I0(GND_net), .I1(n15384[17]), .I2(GND_net), 
            .I3(n51165), .O(n14585[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29335_4_lut (.I0(PWMLimit[15]), .I1(n60589), .I2(n27857), 
            .I3(n11608), .O(n49[15]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29335_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6183_20 (.CI(n51165), .I0(n15384[17]), .I1(GND_net), 
            .CO(n51166));
    SB_LUT4 add_6183_19_lut (.I0(GND_net), .I1(n15384[16]), .I2(GND_net), 
            .I3(n51164), .O(n14585[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_19 (.CI(n51164), .I0(n15384[16]), .I1(GND_net), 
            .CO(n51165));
    SB_LUT4 add_6183_18_lut (.I0(GND_net), .I1(n15384[15]), .I2(GND_net), 
            .I3(n51163), .O(n14585[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51278_4_lut (.I0(n13_adj_4509), .I1(n11_adj_4504), .I2(n9_adj_4517), 
            .I3(n66121), .O(n67006));
    defparam i51278_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_6183_18 (.CI(n51163), .I0(n15384[15]), .I1(GND_net), 
            .CO(n51164));
    SB_LUT4 add_6183_17_lut (.I0(GND_net), .I1(n15384[14]), .I2(GND_net), 
            .I3(n51162), .O(n14585[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_17 (.CI(n51162), .I0(n15384[14]), .I1(GND_net), 
            .CO(n51163));
    SB_LUT4 add_6183_16_lut (.I0(GND_net), .I1(n15384[13]), .I2(n1105_adj_4532), 
            .I3(n51161), .O(n14585[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51260_4_lut (.I0(n19_adj_4520), .I1(n17_adj_4519), .I2(n15_adj_4511), 
            .I3(n67006), .O(n66988));
    defparam i51260_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_6183_16 (.CI(n51161), .I0(n15384[13]), .I1(n1105_adj_4532), 
            .CO(n51162));
    SB_LUT4 add_6183_15_lut (.I0(GND_net), .I1(n15384[12]), .I2(n1032_adj_4533), 
            .I3(n51160), .O(n14585[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_15 (.CI(n51160), .I0(n15384[12]), .I1(n1032_adj_4533), 
            .CO(n51161));
    SB_LUT4 add_6183_14_lut (.I0(GND_net), .I1(n15384[11]), .I2(n959_adj_4534), 
            .I3(n51159), .O(n14585[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_14 (.CI(n51159), .I0(n15384[11]), .I1(n959_adj_4534), 
            .CO(n51160));
    SB_LUT4 add_6183_13_lut (.I0(GND_net), .I1(n15384[10]), .I2(n886_adj_4535), 
            .I3(n51158), .O(n14585[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_13 (.CI(n51158), .I0(n15384[10]), .I1(n886_adj_4535), 
            .CO(n51159));
    SB_LUT4 add_6183_12_lut (.I0(GND_net), .I1(n15384[9]), .I2(n813_adj_4536), 
            .I3(n51157), .O(n14585[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_12 (.CI(n51157), .I0(n15384[9]), .I1(n813_adj_4536), 
            .CO(n51158));
    SB_LUT4 i52507_4_lut (.I0(n25_adj_4499), .I1(n23_adj_4496), .I2(n21_adj_4521), 
            .I3(n66988), .O(n68235));
    defparam i52507_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6183_11_lut (.I0(GND_net), .I1(n15384[8]), .I2(n740_adj_4537), 
            .I3(n51156), .O(n14585[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51892_4_lut (.I0(n31_adj_4501), .I1(n29_adj_4500), .I2(n27_adj_4513), 
            .I3(n68235), .O(n67620));
    defparam i51892_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_6183_11 (.CI(n51156), .I0(n15384[8]), .I1(n740_adj_4537), 
            .CO(n51157));
    SB_LUT4 add_6183_10_lut (.I0(GND_net), .I1(n15384[7]), .I2(n667_adj_4538), 
            .I3(n51155), .O(n14585[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_10 (.CI(n51155), .I0(n15384[7]), .I1(n667_adj_4538), 
            .CO(n51156));
    SB_LUT4 add_6183_9_lut (.I0(GND_net), .I1(n15384[6]), .I2(n594_adj_4539), 
            .I3(n51154), .O(n14585[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_9 (.CI(n51154), .I0(n15384[6]), .I1(n594_adj_4539), 
            .CO(n51155));
    SB_LUT4 add_6183_8_lut (.I0(GND_net), .I1(n15384[5]), .I2(n521_adj_4540), 
            .I3(n51153), .O(n14585[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52684_4_lut (.I0(n37_adj_4495), .I1(n35_adj_4502), .I2(n33_adj_4503), 
            .I3(n67620), .O(n68412));
    defparam i52684_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43_c), 
            .I3(GND_net), .O(n16_adj_4541));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51940_3_lut (.I0(n6_adj_4542), .I1(n130[10]), .I2(n21_adj_4521), 
            .I3(GND_net), .O(n67668));   // verilog/motorControl.v(45[12:34])
    defparam i51940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51941_3_lut (.I0(n67668), .I1(n130[11]), .I2(n23_adj_4496), 
            .I3(GND_net), .O(n67669));   // verilog/motorControl.v(45[12:34])
    defparam i51941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_4519), 
            .I3(GND_net), .O(n8_adj_4543));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_4541), .I1(n130[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4544));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50302_4_lut (.I0(n43_c), .I1(n25_adj_4499), .I2(n23_adj_4496), 
            .I3(n66088), .O(n66030));
    defparam i50302_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51850_4_lut (.I0(n24_adj_4544), .I1(n8_adj_4543), .I2(n45), 
            .I3(n66024), .O(n67578));   // verilog/motorControl.v(45[12:34])
    defparam i51850_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51122_3_lut (.I0(n67669), .I1(n130[12]), .I2(n25_adj_4499), 
            .I3(GND_net), .O(n66850));   // verilog/motorControl.v(45[12:34])
    defparam i51122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4546));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i51936_3_lut (.I0(n4_adj_4546), .I1(n130[13]), .I2(n27_adj_4513), 
            .I3(GND_net), .O(n67664));   // verilog/motorControl.v(45[12:34])
    defparam i51936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51937_3_lut (.I0(n67664), .I1(n130[14]), .I2(n29_adj_4500), 
            .I3(GND_net), .O(n67665));   // verilog/motorControl.v(45[12:34])
    defparam i51937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50331_4_lut (.I0(n33_adj_4503), .I1(n31_adj_4501), .I2(n29_adj_4500), 
            .I3(n66069), .O(n66059));
    defparam i50331_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52421_4_lut (.I0(n30_adj_4529), .I1(n10_adj_4526), .I2(n35_adj_4502), 
            .I3(n66057), .O(n68149));   // verilog/motorControl.v(45[12:34])
    defparam i52421_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51124_3_lut (.I0(n67665), .I1(n130[15]), .I2(n31_adj_4501), 
            .I3(GND_net), .O(n66852));   // verilog/motorControl.v(45[12:34])
    defparam i51124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52774_4_lut (.I0(n66852), .I1(n68149), .I2(n35_adj_4502), 
            .I3(n66059), .O(n68502));   // verilog/motorControl.v(45[12:34])
    defparam i52774_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52775_3_lut (.I0(n68502), .I1(n130[18]), .I2(n37_adj_4495), 
            .I3(GND_net), .O(n68503));   // verilog/motorControl.v(45[12:34])
    defparam i52775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52693_3_lut (.I0(n68503), .I1(n130[19]), .I2(n39), .I3(GND_net), 
            .O(n68421));   // verilog/motorControl.v(45[12:34])
    defparam i52693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50307_4_lut (.I0(n43_c), .I1(n41_adj_4494), .I2(n39), .I3(n68412), 
            .O(n66035));
    defparam i50307_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52475_4_lut (.I0(n66850), .I1(n67578), .I2(n45), .I3(n66030), 
            .O(n68203));   // verilog/motorControl.v(45[12:34])
    defparam i52475_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51130_3_lut (.I0(n68421), .I1(n130[20]), .I2(n41_adj_4494), 
            .I3(GND_net), .O(n66858));   // verilog/motorControl.v(45[12:34])
    defparam i51130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52676_4_lut (.I0(n66858), .I1(n68203), .I2(n45), .I3(n66035), 
            .O(n68404));   // verilog/motorControl.v(45[12:34])
    defparam i52676_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52677_3_lut (.I0(n68404), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(45[12:34])
    defparam i52677_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4547));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4548));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4549));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4550));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4551));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4552));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4553));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50757_2_lut_4_lut (.I0(n356[21]), .I1(n436[21]), .I2(n356[9]), 
            .I3(n436[9]), .O(n66485));
    defparam i50757_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4555));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4556));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4557));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4558));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4559));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4560));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4561));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4562));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4563));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4564));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4565));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4566));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50278_4_lut (.I0(n21_adj_4562), .I1(n19_adj_4561), .I2(n17_adj_4560), 
            .I3(n9_adj_4559), .O(n66006));
    defparam i50278_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50190_4_lut (.I0(n27_adj_4558), .I1(n15_adj_4557), .I2(n13_adj_4556), 
            .I3(n11_adj_4555), .O(n65918));
    defparam i50190_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_4564), 
            .I3(GND_net), .O(n12_adj_4567));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6183_8 (.CI(n51153), .I0(n15384[5]), .I1(n521_adj_4540), 
            .CO(n51154));
    SB_LUT4 add_6183_7_lut (.I0(GND_net), .I1(n15384[4]), .I2(n448_adj_4568), 
            .I3(n51152), .O(n14585[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_7 (.CI(n51152), .I0(n15384[4]), .I1(n448_adj_4568), 
            .CO(n51153));
    SB_LUT4 add_6183_6_lut (.I0(GND_net), .I1(n15384[3]), .I2(n375_adj_4569), 
            .I3(n51151), .O(n14585[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_6 (.CI(n51151), .I0(n15384[3]), .I1(n375_adj_4569), 
            .CO(n51152));
    SB_CARRY add_18_5 (.CI(n49607), .I0(n257[3]), .I1(n306[3]), .CO(n49608));
    SB_LUT4 add_6183_5_lut (.I0(GND_net), .I1(n15384[2]), .I2(n302_adj_4570), 
            .I3(n51150), .O(n14585[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_5 (.CI(n51150), .I0(n15384[2]), .I1(n302_adj_4570), 
            .CO(n51151));
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n306[2]), .I3(n49606), 
            .O(n356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6183_4_lut (.I0(GND_net), .I1(n15384[1]), .I2(n229), .I3(n51149), 
            .O(n14585[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_4 (.CI(n51149), .I0(n15384[1]), .I1(n229), .CO(n51150));
    SB_LUT4 add_6183_3_lut (.I0(GND_net), .I1(n15384[0]), .I2(n156), .I3(n51148), 
            .O(n14585[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_3 (.CI(n51148), .I0(n15384[0]), .I1(n156), .CO(n51149));
    SB_LUT4 add_6183_2_lut (.I0(GND_net), .I1(n14_adj_4571), .I2(n83), 
            .I3(GND_net), .O(n14585[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_2 (.CI(GND_net), .I0(n14_adj_4571), .I1(n83), .CO(n51148));
    SB_LUT4 add_6221_20_lut (.I0(GND_net), .I1(n16105[17]), .I2(GND_net), 
            .I3(n51147), .O(n15384[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6221_19_lut (.I0(GND_net), .I1(n16105[16]), .I2(GND_net), 
            .I3(n51146), .O(n15384[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50774_2_lut_4_lut (.I0(n356[16]), .I1(n436[16]), .I2(n356[7]), 
            .I3(n436[7]), .O(n66502));
    defparam i50774_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i13786_3_lut (.I0(n356[16]), .I1(n436[16]), .I2(n11610), .I3(GND_net), 
            .O(n27852));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29334_4_lut (.I0(PWMLimit[16]), .I1(n60589), .I2(n27852), 
            .I3(n11608), .O(n49[16]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29334_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_4556), 
            .I3(GND_net), .O(n10_adj_4572));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_4567), .I1(n182[17]), .I2(n35_adj_4565), 
            .I3(GND_net), .O(n30_adj_4573));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6221_19 (.CI(n51146), .I0(n16105[16]), .I1(GND_net), 
            .CO(n51147));
    SB_LUT4 add_6221_18_lut (.I0(GND_net), .I1(n16105[15]), .I2(GND_net), 
            .I3(n51145), .O(n15384[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_18 (.CI(n51145), .I0(n16105[15]), .I1(GND_net), 
            .CO(n51146));
    SB_LUT4 add_6221_17_lut (.I0(GND_net), .I1(n16105[14]), .I2(GND_net), 
            .I3(n51144), .O(n15384[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_17 (.CI(n51144), .I0(n16105[14]), .I1(GND_net), 
            .CO(n51145));
    SB_LUT4 add_6221_16_lut (.I0(GND_net), .I1(n16105[13]), .I2(n1108), 
            .I3(n51143), .O(n15384[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_16 (.CI(n51143), .I0(n16105[13]), .I1(n1108), .CO(n51144));
    SB_LUT4 add_6221_15_lut (.I0(GND_net), .I1(n16105[12]), .I2(n1035), 
            .I3(n51142), .O(n15384[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_15 (.CI(n51142), .I0(n16105[12]), .I1(n1035), .CO(n51143));
    SB_LUT4 add_6221_14_lut (.I0(GND_net), .I1(n16105[11]), .I2(n962), 
            .I3(n51141), .O(n15384[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_14 (.CI(n51141), .I0(n16105[11]), .I1(n962), .CO(n51142));
    SB_LUT4 add_6221_13_lut (.I0(GND_net), .I1(n16105[10]), .I2(n889), 
            .I3(n51140), .O(n15384[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_13 (.CI(n51140), .I0(n16105[10]), .I1(n889), .CO(n51141));
    SB_LUT4 add_6221_12_lut (.I0(GND_net), .I1(n16105[9]), .I2(n816), 
            .I3(n51139), .O(n15384[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_12 (.CI(n51139), .I0(n16105[9]), .I1(n816), .CO(n51140));
    SB_LUT4 add_6221_11_lut (.I0(GND_net), .I1(n16105[8]), .I2(n743), 
            .I3(n51138), .O(n15384[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_11 (.CI(n51138), .I0(n16105[8]), .I1(n743), .CO(n51139));
    SB_LUT4 add_6221_10_lut (.I0(GND_net), .I1(n16105[7]), .I2(n670), 
            .I3(n51137), .O(n15384[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_10 (.CI(n51137), .I0(n16105[7]), .I1(n670), .CO(n51138));
    SB_LUT4 add_6221_9_lut (.I0(GND_net), .I1(n16105[6]), .I2(n597), .I3(n51136), 
            .O(n15384[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_9 (.CI(n51136), .I0(n16105[6]), .I1(n597), .CO(n51137));
    SB_LUT4 add_6221_8_lut (.I0(GND_net), .I1(n16105[5]), .I2(n524), .I3(n51135), 
            .O(n15384[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_8 (.CI(n51135), .I0(n16105[5]), .I1(n524), .CO(n51136));
    SB_LUT4 add_6221_7_lut (.I0(GND_net), .I1(n16105[4]), .I2(n451_adj_4574), 
            .I3(n51134), .O(n15384[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_7 (.CI(n51134), .I0(n16105[4]), .I1(n451_adj_4574), 
            .CO(n51135));
    SB_CARRY add_18_4 (.CI(n49606), .I0(n257[2]), .I1(n306[2]), .CO(n49607));
    SB_LUT4 add_6507_9_lut (.I0(GND_net), .I1(n20032[6]), .I2(n630), .I3(n49924), 
            .O(n19905[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6221_6_lut (.I0(GND_net), .I1(n16105[3]), .I2(n378_adj_4575), 
            .I3(n51133), .O(n15384[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_6 (.CI(n51133), .I0(n16105[3]), .I1(n378_adj_4575), 
            .CO(n51134));
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n306[1]), .I3(n49605), 
            .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6221_5_lut (.I0(GND_net), .I1(n16105[2]), .I2(n305), .I3(n51132), 
            .O(n15384[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_5 (.CI(n51132), .I0(n16105[2]), .I1(n305), .CO(n51133));
    SB_CARRY add_18_3 (.CI(n49605), .I0(n257[1]), .I1(n306[1]), .CO(n49606));
    SB_LUT4 add_6221_4_lut (.I0(GND_net), .I1(n16105[1]), .I2(n232), .I3(n51131), 
            .O(n15384[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13781_3_lut (.I0(n356[17]), .I1(n436[17]), .I2(n11610), .I3(GND_net), 
            .O(n27847));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13781_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6221_4 (.CI(n51131), .I0(n16105[1]), .I1(n232), .CO(n51132));
    SB_LUT4 add_6221_3_lut (.I0(GND_net), .I1(n16105[0]), .I2(n159), .I3(n51130), 
            .O(n15384[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_3 (.CI(n51130), .I0(n16105[0]), .I1(n159), .CO(n51131));
    SB_LUT4 add_6221_2_lut (.I0(GND_net), .I1(n17_adj_4576), .I2(n86), 
            .I3(GND_net), .O(n15384[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29333_4_lut (.I0(PWMLimit[17]), .I1(n60589), .I2(n27847), 
            .I3(n11608), .O(n49[17]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29333_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n306[0]), .I3(GND_net), 
            .O(n380)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_2 (.CI(GND_net), .I0(n17_adj_4576), .I1(n86), .CO(n51130));
    SB_LUT4 add_6482_10_lut (.I0(GND_net), .I1(n19825[7]), .I2(n700_adj_4578), 
            .I3(n51129), .O(n19645[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13776_3_lut (.I0(n356[18]), .I1(n436[18]), .I2(n11610), .I3(GND_net), 
            .O(n27842));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29332_4_lut (.I0(PWMLimit[18]), .I1(n60589), .I2(n27842), 
            .I3(n11608), .O(n49[18]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29332_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13771_3_lut (.I0(n356[19]), .I1(n436[19]), .I2(n11610), .I3(GND_net), 
            .O(n27837));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29331_4_lut (.I0(PWMLimit[19]), .I1(n60589), .I2(n27837), 
            .I3(n11608), .O(n49[19]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29331_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13766_3_lut (.I0(n356[20]), .I1(n436[20]), .I2(n11610), .I3(GND_net), 
            .O(n27832));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29330_4_lut (.I0(PWMLimit[20]), .I1(n60589), .I2(n27832), 
            .I3(n11608), .O(n49[20]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29330_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6507_8_lut (.I0(GND_net), .I1(n20032[5]), .I2(n557), .I3(n49923), 
            .O(n19905[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6482_9_lut (.I0(GND_net), .I1(n19825[6]), .I2(n627_adj_4582), 
            .I3(n51128), .O(n19645[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_9 (.CI(n51128), .I0(n19825[6]), .I1(n627_adj_4582), 
            .CO(n51129));
    SB_LUT4 add_6482_8_lut (.I0(GND_net), .I1(n19825[5]), .I2(n554_adj_4583), 
            .I3(n51127), .O(n19645[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_8 (.CI(n51127), .I0(n19825[5]), .I1(n554_adj_4583), 
            .CO(n51128));
    SB_LUT4 add_6482_7_lut (.I0(GND_net), .I1(n19825[4]), .I2(n481_adj_4584), 
            .I3(n51126), .O(n19645[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_7 (.CI(n51126), .I0(n19825[4]), .I1(n481_adj_4584), 
            .CO(n51127));
    SB_LUT4 add_6482_6_lut (.I0(GND_net), .I1(n19825[3]), .I2(n408_adj_4585), 
            .I3(n51125), .O(n19645[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_6 (.CI(n51125), .I0(n19825[3]), .I1(n408_adj_4585), 
            .CO(n51126));
    SB_LUT4 add_6482_5_lut (.I0(GND_net), .I1(n19825[2]), .I2(n335_adj_4586), 
            .I3(n51124), .O(n19645[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_8 (.CI(n49923), .I0(n20032[5]), .I1(n557), .CO(n49924));
    SB_CARRY add_6482_5 (.CI(n51124), .I0(n19825[2]), .I1(n335_adj_4586), 
            .CO(n51125));
    SB_LUT4 add_6482_4_lut (.I0(GND_net), .I1(n19825[1]), .I2(n262_adj_4587), 
            .I3(n51123), .O(n19645[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6507_7_lut (.I0(GND_net), .I1(n20032[4]), .I2(n484), .I3(n49922), 
            .O(n19905[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_7 (.CI(n49922), .I0(n20032[4]), .I1(n484), .CO(n49923));
    SB_LUT4 add_6507_6_lut (.I0(GND_net), .I1(n20032[3]), .I2(n411), .I3(n49921), 
            .O(n19905[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_6 (.CI(n49921), .I0(n20032[3]), .I1(n411), .CO(n49922));
    SB_LUT4 i51192_4_lut (.I0(n13_adj_4556), .I1(n11_adj_4555), .I2(n9_adj_4559), 
            .I3(n66022), .O(n66920));
    defparam i51192_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i13761_3_lut (.I0(n356[21]), .I1(n436[21]), .I2(n11610), .I3(GND_net), 
            .O(n27827));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51186_4_lut (.I0(n19_adj_4561), .I1(n17_adj_4560), .I2(n15_adj_4557), 
            .I3(n66920), .O(n66914));
    defparam i51186_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29329_4_lut (.I0(PWMLimit[21]), .I1(n60589), .I2(n27827), 
            .I3(n11608), .O(n49[21]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29329_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6482_4 (.CI(n51123), .I0(n19825[1]), .I1(n262_adj_4587), 
            .CO(n51124));
    SB_LUT4 i13756_3_lut (.I0(n356[22]), .I1(n436[22]), .I2(n11610), .I3(GND_net), 
            .O(n27822));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6482_3_lut (.I0(GND_net), .I1(n19825[0]), .I2(n189_adj_4589), 
            .I3(n51122), .O(n19645[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29328_4_lut (.I0(PWMLimit[22]), .I1(n60589), .I2(n27822), 
            .I3(n11608), .O(n49[22]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29328_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6482_3 (.CI(n51122), .I0(n19825[0]), .I1(n189_adj_4589), 
            .CO(n51123));
    SB_LUT4 i52471_4_lut (.I0(n25_adj_4553), .I1(n23_adj_4563), .I2(n21_adj_4562), 
            .I3(n66914), .O(n68199));
    defparam i52471_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6482_2_lut (.I0(GND_net), .I1(n47_adj_4590), .I2(n116_adj_4591), 
            .I3(GND_net), .O(n19645[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_2 (.CI(GND_net), .I0(n47_adj_4590), .I1(n116_adj_4591), 
            .CO(n51122));
    SB_LUT4 mult_16_add_1225_24_lut (.I0(n1[23]), .I1(n12157[21]), .I2(GND_net), 
            .I3(n50187), .O(n11650[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6257_19_lut (.I0(GND_net), .I1(n16752[16]), .I2(GND_net), 
            .I3(n51121), .O(n16105[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6257_18_lut (.I0(GND_net), .I1(n16752[15]), .I2(GND_net), 
            .I3(n51120), .O(n16105[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_18 (.CI(n51120), .I0(n16752[15]), .I1(GND_net), 
            .CO(n51121));
    SB_LUT4 add_6257_17_lut (.I0(GND_net), .I1(n16752[14]), .I2(GND_net), 
            .I3(n51119), .O(n16105[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_17 (.CI(n51119), .I0(n16752[14]), .I1(GND_net), 
            .CO(n51120));
    SB_LUT4 add_6257_16_lut (.I0(GND_net), .I1(n16752[13]), .I2(n1111), 
            .I3(n51118), .O(n16105[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_23_lut (.I0(GND_net), .I1(n12157[20]), .I2(GND_net), 
            .I3(n50186), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_16 (.CI(n51118), .I0(n16752[13]), .I1(n1111), .CO(n51119));
    SB_LUT4 add_6257_15_lut (.I0(GND_net), .I1(n16752[12]), .I2(n1038), 
            .I3(n51117), .O(n16105[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6507_5_lut (.I0(GND_net), .I1(n20032[2]), .I2(n338_adj_4592), 
            .I3(n49920), .O(n19905[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51826_4_lut (.I0(n31_adj_4552), .I1(n29_adj_4551), .I2(n27_adj_4558), 
            .I3(n68199), .O(n67554));
    defparam i51826_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_6257_15 (.CI(n51117), .I0(n16752[12]), .I1(n1038), .CO(n51118));
    SB_LUT4 add_6257_14_lut (.I0(GND_net), .I1(n16752[11]), .I2(n965), 
            .I3(n51116), .O(n16105[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_14 (.CI(n51116), .I0(n16752[11]), .I1(n965), .CO(n51117));
    SB_LUT4 i52668_4_lut (.I0(n37_adj_4566), .I1(n35_adj_4565), .I2(n33_adj_4564), 
            .I3(n67554), .O(n68396));
    defparam i52668_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6257_13_lut (.I0(GND_net), .I1(n16752[10]), .I2(n892), 
            .I3(n51115), .O(n16105[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_23 (.CI(n50186), .I0(n12157[20]), .I1(GND_net), 
            .CO(n50187));
    SB_CARRY add_6257_13 (.CI(n51115), .I0(n16752[10]), .I1(n892), .CO(n51116));
    SB_LUT4 add_6257_12_lut (.I0(GND_net), .I1(n16752[9]), .I2(n819), 
            .I3(n51114), .O(n16105[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_22_lut (.I0(GND_net), .I1(n12157[19]), .I2(GND_net), 
            .I3(n50185), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_12 (.CI(n51114), .I0(n16752[9]), .I1(n819), .CO(n51115));
    SB_CARRY add_6507_5 (.CI(n49920), .I0(n20032[2]), .I1(n338_adj_4592), 
            .CO(n49921));
    SB_CARRY mult_16_add_1225_22 (.CI(n50185), .I0(n12157[19]), .I1(GND_net), 
            .CO(n50186));
    SB_LUT4 mult_16_add_1225_21_lut (.I0(GND_net), .I1(n12157[18]), .I2(GND_net), 
            .I3(n50184), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6257_11_lut (.I0(GND_net), .I1(n16752[8]), .I2(n746), 
            .I3(n51113), .O(n16105[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6507_4_lut (.I0(GND_net), .I1(n20032[1]), .I2(n265), .I3(n49919), 
            .O(n19905[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_4 (.CI(n49919), .I0(n20032[1]), .I1(n265), .CO(n49920));
    SB_CARRY mult_16_add_1225_21 (.CI(n50184), .I0(n12157[18]), .I1(GND_net), 
            .CO(n50185));
    SB_LUT4 add_6507_3_lut (.I0(GND_net), .I1(n20032[0]), .I2(n192_adj_4593), 
            .I3(n49918), .O(n19905[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_11 (.CI(n51113), .I0(n16752[8]), .I1(n746), .CO(n51114));
    SB_CARRY add_6507_3 (.CI(n49918), .I0(n20032[0]), .I1(n192_adj_4593), 
            .CO(n49919));
    SB_LUT4 add_6507_2_lut (.I0(GND_net), .I1(n50_adj_4594), .I2(n119_adj_4595), 
            .I3(GND_net), .O(n19905[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6257_10_lut (.I0(GND_net), .I1(n16752[7]), .I2(n673), 
            .I3(n51112), .O(n16105[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43_adj_4550), 
            .I3(GND_net), .O(n16_adj_4596));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4597));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6257_10 (.CI(n51112), .I0(n16752[7]), .I1(n673), .CO(n51113));
    SB_LUT4 add_6257_9_lut (.I0(GND_net), .I1(n16752[6]), .I2(n600), .I3(n51111), 
            .O(n16105[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_9 (.CI(n51111), .I0(n16752[6]), .I1(n600), .CO(n51112));
    SB_LUT4 mult_16_add_1225_20_lut (.I0(GND_net), .I1(n12157[17]), .I2(GND_net), 
            .I3(n50183), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6257_8_lut (.I0(GND_net), .I1(n16752[5]), .I2(n527_adj_4598), 
            .I3(n51110), .O(n16105[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52469_3_lut (.I0(n6_adj_4599), .I1(n182[10]), .I2(n21_adj_4562), 
            .I3(GND_net), .O(n68197));   // verilog/motorControl.v(47[21:44])
    defparam i52469_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_16_add_1225_20 (.CI(n50183), .I0(n12157[17]), .I1(GND_net), 
            .CO(n50184));
    SB_CARRY add_6507_2 (.CI(GND_net), .I0(n50_adj_4594), .I1(n119_adj_4595), 
            .CO(n49918));
    SB_LUT4 mult_16_add_1225_19_lut (.I0(GND_net), .I1(n12157[16]), .I2(GND_net), 
            .I3(n50182), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_16_lut (.I0(GND_net), .I1(n18065[13]), .I2(n1120), 
            .I3(n49917), .O(n17585[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_8 (.CI(n51110), .I0(n16752[5]), .I1(n527_adj_4598), 
            .CO(n51111));
    SB_LUT4 add_6257_7_lut (.I0(GND_net), .I1(n16752[4]), .I2(n454_adj_4600), 
            .I3(n51109), .O(n16105[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_7 (.CI(n51109), .I0(n16752[4]), .I1(n454_adj_4600), 
            .CO(n51110));
    SB_LUT4 add_6338_15_lut (.I0(GND_net), .I1(n18065[12]), .I2(n1047), 
            .I3(n49916), .O(n17585[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_19 (.CI(n50182), .I0(n12157[16]), .I1(GND_net), 
            .CO(n50183));
    SB_LUT4 add_6257_6_lut (.I0(GND_net), .I1(n16752[3]), .I2(n381_adj_4601), 
            .I3(n51108), .O(n16105[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_15 (.CI(n49916), .I0(n18065[12]), .I1(n1047), .CO(n49917));
    SB_LUT4 mult_16_add_1225_18_lut (.I0(GND_net), .I1(n12157[15]), .I2(GND_net), 
            .I3(n50181), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_14_lut (.I0(GND_net), .I1(n18065[11]), .I2(n974), 
            .I3(n49915), .O(n17585[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_6 (.CI(n51108), .I0(n16752[3]), .I1(n381_adj_4601), 
            .CO(n51109));
    SB_LUT4 add_6257_5_lut (.I0(GND_net), .I1(n16752[2]), .I2(n308_adj_4602), 
            .I3(n51107), .O(n16105[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_5 (.CI(n51107), .I0(n16752[2]), .I1(n308_adj_4602), 
            .CO(n51108));
    SB_CARRY mult_16_add_1225_18 (.CI(n50181), .I0(n12157[15]), .I1(GND_net), 
            .CO(n50182));
    SB_LUT4 mult_16_add_1225_17_lut (.I0(GND_net), .I1(n12157[14]), .I2(GND_net), 
            .I3(n50180), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_14 (.CI(n49915), .I0(n18065[11]), .I1(n974), .CO(n49916));
    SB_LUT4 add_6257_4_lut (.I0(GND_net), .I1(n16752[1]), .I2(n235_adj_4603), 
            .I3(n51106), .O(n16105[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_4 (.CI(n51106), .I0(n16752[1]), .I1(n235_adj_4603), 
            .CO(n51107));
    SB_CARRY mult_16_add_1225_17 (.CI(n50180), .I0(n12157[14]), .I1(GND_net), 
            .CO(n50181));
    SB_LUT4 add_6338_13_lut (.I0(GND_net), .I1(n18065[10]), .I2(n901), 
            .I3(n49914), .O(n17585[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_16_lut (.I0(GND_net), .I1(n12157[13]), .I2(n1096_adj_4604), 
            .I3(n50179), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_13 (.CI(n49914), .I0(n18065[10]), .I1(n901), .CO(n49915));
    SB_LUT4 add_6338_12_lut (.I0(GND_net), .I1(n18065[9]), .I2(n828), 
            .I3(n49913), .O(n17585[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6257_3_lut (.I0(GND_net), .I1(n16752[0]), .I2(n162_adj_4605), 
            .I3(n51105), .O(n16105[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_3 (.CI(n51105), .I0(n16752[0]), .I1(n162_adj_4605), 
            .CO(n51106));
    SB_CARRY add_6338_12 (.CI(n49913), .I0(n18065[9]), .I1(n828), .CO(n49914));
    SB_LUT4 add_6257_2_lut (.I0(GND_net), .I1(n20_adj_4606), .I2(n89_adj_4607), 
            .I3(GND_net), .O(n16105[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_11_lut (.I0(GND_net), .I1(n18065[8]), .I2(n755), 
            .I3(n49912), .O(n17585[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_2 (.CI(GND_net), .I0(n20_adj_4606), .I1(n89_adj_4607), 
            .CO(n51105));
    SB_CARRY add_6338_11 (.CI(n49912), .I0(n18065[8]), .I1(n755), .CO(n49913));
    SB_LUT4 add_6291_18_lut (.I0(GND_net), .I1(n17329[15]), .I2(GND_net), 
            .I3(n51104), .O(n16752[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n306[0]), .CO(n49605));
    SB_LUT4 add_6291_17_lut (.I0(GND_net), .I1(n17329[14]), .I2(GND_net), 
            .I3(n51103), .O(n16752[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_16 (.CI(n50179), .I0(n12157[13]), .I1(n1096_adj_4604), 
            .CO(n50180));
    SB_LUT4 add_6338_10_lut (.I0(GND_net), .I1(n18065[7]), .I2(n682), 
            .I3(n49911), .O(n17585[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_15_lut (.I0(GND_net), .I1(n12157[12]), .I2(n1023_adj_4608), 
            .I3(n50178), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_15 (.CI(n50178), .I0(n12157[12]), .I1(n1023_adj_4608), 
            .CO(n50179));
    SB_CARRY add_6291_17 (.CI(n51103), .I0(n17329[14]), .I1(GND_net), 
            .CO(n51104));
    SB_LUT4 add_6291_16_lut (.I0(GND_net), .I1(n17329[13]), .I2(n1114_adj_4609), 
            .I3(n51102), .O(n16752[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_14_lut (.I0(GND_net), .I1(n12157[11]), .I2(n950_adj_4610), 
            .I3(n50177), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_14 (.CI(n50177), .I0(n12157[11]), .I1(n950_adj_4610), 
            .CO(n50178));
    SB_LUT4 i52470_3_lut (.I0(n68197), .I1(n182[11]), .I2(n23_adj_4563), 
            .I3(GND_net), .O(n68198));   // verilog/motorControl.v(47[21:44])
    defparam i52470_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6291_16 (.CI(n51102), .I0(n17329[13]), .I1(n1114_adj_4609), 
            .CO(n51103));
    SB_LUT4 mult_16_add_1225_13_lut (.I0(GND_net), .I1(n12157[10]), .I2(n877_adj_4611), 
            .I3(n50176), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_13 (.CI(n50176), .I0(n12157[10]), .I1(n877_adj_4611), 
            .CO(n50177));
    SB_LUT4 mult_16_add_1225_12_lut (.I0(GND_net), .I1(n12157[9]), .I2(n804_adj_4612), 
            .I3(n50175), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_12 (.CI(n50175), .I0(n12157[9]), .I1(n804_adj_4612), 
            .CO(n50176));
    SB_LUT4 add_6291_15_lut (.I0(GND_net), .I1(n17329[12]), .I2(n1041_adj_4613), 
            .I3(n51101), .O(n16752[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_15 (.CI(n51101), .I0(n17329[12]), .I1(n1041_adj_4613), 
            .CO(n51102));
    SB_LUT4 add_6291_14_lut (.I0(GND_net), .I1(n17329[11]), .I2(n968_adj_4614), 
            .I3(n51100), .O(n16752[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_11_lut (.I0(GND_net), .I1(n12157[8]), .I2(n731_adj_4615), 
            .I3(n50174), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_11 (.CI(n50174), .I0(n12157[8]), .I1(n731_adj_4615), 
            .CO(n50175));
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n1[23]), .I3(n49604), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_10_lut (.I0(GND_net), .I1(n12157[7]), .I2(n658_adj_4616), 
            .I3(n50173), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_10 (.CI(n49911), .I0(n18065[7]), .I1(n682), .CO(n49912));
    SB_CARRY mult_16_add_1225_10 (.CI(n50173), .I0(n12157[7]), .I1(n658_adj_4616), 
            .CO(n50174));
    SB_LUT4 mult_16_add_1225_9_lut (.I0(GND_net), .I1(n12157[6]), .I2(n585_adj_4617), 
            .I3(n50172), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_14 (.CI(n51100), .I0(n17329[11]), .I1(n968_adj_4614), 
            .CO(n51101));
    SB_LUT4 add_6291_13_lut (.I0(GND_net), .I1(n17329[10]), .I2(n895_adj_4618), 
            .I3(n51099), .O(n16752[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_9 (.CI(n50172), .I0(n12157[6]), .I1(n585_adj_4617), 
            .CO(n50173));
    SB_LUT4 mult_16_add_1225_8_lut (.I0(GND_net), .I1(n12157[5]), .I2(n512_adj_4619), 
            .I3(n50171), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_9_lut (.I0(GND_net), .I1(n18065[6]), .I2(n609), .I3(n49910), 
            .O(n17585[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_13 (.CI(n51099), .I0(n17329[10]), .I1(n895_adj_4618), 
            .CO(n51100));
    SB_LUT4 add_6291_12_lut (.I0(GND_net), .I1(n17329[9]), .I2(n822_adj_4620), 
            .I3(n51098), .O(n16752[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_8 (.CI(n50171), .I0(n12157[5]), .I1(n512_adj_4619), 
            .CO(n50172));
    SB_CARRY add_6291_12 (.CI(n51098), .I0(n17329[9]), .I1(n822_adj_4620), 
            .CO(n51099));
    SB_LUT4 add_6291_11_lut (.I0(GND_net), .I1(n17329[8]), .I2(n749_adj_4621), 
            .I3(n51097), .O(n16752[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_11 (.CI(n51097), .I0(n17329[8]), .I1(n749_adj_4621), 
            .CO(n51098));
    SB_CARRY add_6338_9 (.CI(n49910), .I0(n18065[6]), .I1(n609), .CO(n49911));
    SB_LUT4 mult_16_add_1225_7_lut (.I0(GND_net), .I1(n12157[4]), .I2(n439_adj_4622), 
            .I3(n50170), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6291_10_lut (.I0(GND_net), .I1(n17329[7]), .I2(n676_adj_4623), 
            .I3(n51096), .O(n16752[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_10 (.CI(n51096), .I0(n17329[7]), .I1(n676_adj_4623), 
            .CO(n51097));
    SB_LUT4 add_6291_9_lut (.I0(GND_net), .I1(n17329[6]), .I2(n603_adj_4624), 
            .I3(n51095), .O(n16752[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_9 (.CI(n51095), .I0(n17329[6]), .I1(n603_adj_4624), 
            .CO(n51096));
    SB_LUT4 add_6291_8_lut (.I0(GND_net), .I1(n17329[5]), .I2(n530_adj_4625), 
            .I3(n51094), .O(n16752[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_8 (.CI(n51094), .I0(n17329[5]), .I1(n530_adj_4625), 
            .CO(n51095));
    SB_LUT4 add_6291_7_lut (.I0(GND_net), .I1(n17329[4]), .I2(n457_adj_4626), 
            .I3(n51093), .O(n16752[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_7 (.CI(n51093), .I0(n17329[4]), .I1(n457_adj_4626), 
            .CO(n51094));
    SB_CARRY mult_16_add_1225_7 (.CI(n50170), .I0(n12157[4]), .I1(n439_adj_4622), 
            .CO(n50171));
    SB_LUT4 add_6291_6_lut (.I0(GND_net), .I1(n17329[3]), .I2(n384_adj_4627), 
            .I3(n51092), .O(n16752[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_6_lut (.I0(GND_net), .I1(n12157[3]), .I2(n366_adj_4628), 
            .I3(n50169), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_8_lut (.I0(GND_net), .I1(n18065[5]), .I2(n536), .I3(n49909), 
            .O(n17585[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_8 (.CI(n49909), .I0(n18065[5]), .I1(n536), .CO(n49910));
    SB_CARRY mult_16_add_1225_6 (.CI(n50169), .I0(n12157[3]), .I1(n366_adj_4628), 
            .CO(n50170));
    SB_LUT4 mult_16_add_1225_5_lut (.I0(GND_net), .I1(n12157[2]), .I2(n293_adj_4629), 
            .I3(n50168), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_7_lut (.I0(GND_net), .I1(n18065[4]), .I2(n463), .I3(n49908), 
            .O(n17585[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n1[22]), .I3(n49603), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_6 (.CI(n51092), .I0(n17329[3]), .I1(n384_adj_4627), 
            .CO(n51093));
    SB_CARRY mult_16_add_1225_5 (.CI(n50168), .I0(n12157[2]), .I1(n293_adj_4629), 
            .CO(n50169));
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_4560), 
            .I3(GND_net), .O(n8_adj_4630));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_add_1225_4_lut (.I0(GND_net), .I1(n12157[1]), .I2(n220_adj_4631), 
            .I3(n50167), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_4 (.CI(n50167), .I0(n12157[1]), .I1(n220_adj_4631), 
            .CO(n50168));
    SB_LUT4 mult_16_add_1225_3_lut (.I0(GND_net), .I1(n12157[0]), .I2(n147_adj_4632), 
            .I3(n50166), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_3 (.CI(n50166), .I0(n12157[0]), .I1(n147_adj_4632), 
            .CO(n50167));
    SB_LUT4 mult_16_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4633), .I2(n74_adj_4634), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_2 (.CI(GND_net), .I0(n5_adj_4633), .I1(n74_adj_4634), 
            .CO(n50166));
    SB_LUT4 add_6291_5_lut (.I0(GND_net), .I1(n17329[2]), .I2(n311_adj_4635), 
            .I3(n51091), .O(n16752[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_5 (.CI(n51091), .I0(n17329[2]), .I1(n311_adj_4635), 
            .CO(n51092));
    SB_LUT4 add_6291_4_lut (.I0(GND_net), .I1(n17329[1]), .I2(n238_adj_4636), 
            .I3(n51090), .O(n16752[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_4 (.CI(n51090), .I0(n17329[1]), .I1(n238_adj_4636), 
            .CO(n51091));
    SB_LUT4 add_6291_3_lut (.I0(GND_net), .I1(n17329[0]), .I2(n165_adj_4637), 
            .I3(n51089), .O(n16752[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_3 (.CI(n51089), .I0(n17329[0]), .I1(n165_adj_4637), 
            .CO(n51090));
    SB_LUT4 add_6291_2_lut (.I0(GND_net), .I1(n23_adj_4638), .I2(n92_adj_4639), 
            .I3(GND_net), .O(n16752[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_2 (.CI(GND_net), .I0(n23_adj_4638), .I1(n92_adj_4639), 
            .CO(n51089));
    SB_LUT4 add_6499_9_lut (.I0(GND_net), .I1(n19969[6]), .I2(n630_adj_4640), 
            .I3(n51088), .O(n19825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_8_lut (.I0(GND_net), .I1(n19969[5]), .I2(n557_adj_4641), 
            .I3(n51087), .O(n19825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_4596), .I1(n182[22]), .I2(n45_adj_4549), 
            .I3(GND_net), .O(n24_adj_4642));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6499_8 (.CI(n51087), .I0(n19969[5]), .I1(n557_adj_4641), 
            .CO(n51088));
    SB_LUT4 i50142_4_lut (.I0(n43_adj_4550), .I1(n25_adj_4553), .I2(n23_adj_4563), 
            .I3(n66006), .O(n65870));
    defparam i50142_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6499_7_lut (.I0(GND_net), .I1(n19969[4]), .I2(n484_adj_4643), 
            .I3(n51086), .O(n19825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_7 (.CI(n51086), .I0(n19969[4]), .I1(n484_adj_4643), 
            .CO(n51087));
    SB_LUT4 i51852_4_lut (.I0(n24_adj_4642), .I1(n8_adj_4630), .I2(n45_adj_4549), 
            .I3(n65855), .O(n67580));   // verilog/motorControl.v(47[21:44])
    defparam i51852_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_6499_6_lut (.I0(GND_net), .I1(n19969[3]), .I2(n411_adj_4644), 
            .I3(n51085), .O(n19825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_6 (.CI(n51085), .I0(n19969[3]), .I1(n411_adj_4644), 
            .CO(n51086));
    SB_LUT4 add_6499_5_lut (.I0(GND_net), .I1(n19969[2]), .I2(n338_adj_4645), 
            .I3(n51084), .O(n19825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_7 (.CI(n49908), .I0(n18065[4]), .I1(n463), .CO(n49909));
    SB_CARRY add_6499_5 (.CI(n51084), .I0(n19969[2]), .I1(n338_adj_4645), 
            .CO(n51085));
    SB_LUT4 add_6499_4_lut (.I0(GND_net), .I1(n19969[1]), .I2(n265_adj_4646), 
            .I3(n51083), .O(n19825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_4 (.CI(n51083), .I0(n19969[1]), .I1(n265_adj_4646), 
            .CO(n51084));
    SB_LUT4 add_6499_3_lut (.I0(GND_net), .I1(n19969[0]), .I2(n192_adj_4647), 
            .I3(n51082), .O(n19825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_3 (.CI(n51082), .I0(n19969[0]), .I1(n192_adj_4647), 
            .CO(n51083));
    SB_LUT4 add_6499_2_lut (.I0(GND_net), .I1(n50_adj_4648), .I2(n119_adj_4649), 
            .I3(GND_net), .O(n19825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_2 (.CI(GND_net), .I0(n50_adj_4648), .I1(n119_adj_4649), 
            .CO(n51082));
    SB_LUT4 add_6323_17_lut (.I0(GND_net), .I1(n17840[14]), .I2(GND_net), 
            .I3(n51081), .O(n17329[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_16_lut (.I0(GND_net), .I1(n17840[13]), .I2(n1117_adj_4650), 
            .I3(n51080), .O(n17329[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_16 (.CI(n51080), .I0(n17840[13]), .I1(n1117_adj_4650), 
            .CO(n51081));
    SB_LUT4 add_6323_15_lut (.I0(GND_net), .I1(n17840[12]), .I2(n1044_adj_4651), 
            .I3(n51079), .O(n17329[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52169_3_lut (.I0(n68198), .I1(n182[12]), .I2(n25_adj_4553), 
            .I3(GND_net), .O(n67897));   // verilog/motorControl.v(47[21:44])
    defparam i52169_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6323_15 (.CI(n51079), .I0(n17840[12]), .I1(n1044_adj_4651), 
            .CO(n51080));
    SB_LUT4 add_6323_14_lut (.I0(GND_net), .I1(n17840[11]), .I2(n971_adj_4652), 
            .I3(n51078), .O(n17329[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_6_lut (.I0(GND_net), .I1(n18065[3]), .I2(n390_adj_4653), 
            .I3(n49907), .O(n17585[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_4654));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_6323_14 (.CI(n51078), .I0(n17840[11]), .I1(n971_adj_4652), 
            .CO(n51079));
    SB_LUT4 add_6323_13_lut (.I0(GND_net), .I1(n17840[10]), .I2(n898_adj_4655), 
            .I3(n51077), .O(n17329[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_6 (.CI(n49907), .I0(n18065[3]), .I1(n390_adj_4653), 
            .CO(n49908));
    SB_CARRY add_6323_13 (.CI(n51077), .I0(n17840[10]), .I1(n898_adj_4655), 
            .CO(n51078));
    SB_LUT4 add_6323_12_lut (.I0(GND_net), .I1(n17840[9]), .I2(n825_adj_4656), 
            .I3(n51076), .O(n17329[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_12 (.CI(n51076), .I0(n17840[9]), .I1(n825_adj_4656), 
            .CO(n51077));
    SB_LUT4 add_6323_11_lut (.I0(GND_net), .I1(n17840[8]), .I2(n752_adj_4657), 
            .I3(n51075), .O(n17329[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_11 (.CI(n51075), .I0(n17840[8]), .I1(n752_adj_4657), 
            .CO(n51076));
    SB_LUT4 add_6323_10_lut (.I0(GND_net), .I1(n17840[7]), .I2(n679_adj_4658), 
            .I3(n51074), .O(n17329[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_10 (.CI(n51074), .I0(n17840[7]), .I1(n679_adj_4658), 
            .CO(n51075));
    SB_LUT4 i52429_3_lut (.I0(n4_adj_4654), .I1(n182[13]), .I2(n27_adj_4558), 
            .I3(GND_net), .O(n68157));   // verilog/motorControl.v(47[21:44])
    defparam i52429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6323_9_lut (.I0(GND_net), .I1(n17840[6]), .I2(n606_adj_4659), 
            .I3(n51073), .O(n17329[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52430_3_lut (.I0(n68157), .I1(n182[14]), .I2(n29_adj_4551), 
            .I3(GND_net), .O(n68158));   // verilog/motorControl.v(47[21:44])
    defparam i52430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6323_9 (.CI(n51073), .I0(n17840[6]), .I1(n606_adj_4659), 
            .CO(n51074));
    SB_LUT4 add_6323_8_lut (.I0(GND_net), .I1(n17840[5]), .I2(n533_adj_4660), 
            .I3(n51072), .O(n17329[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_8 (.CI(n51072), .I0(n17840[5]), .I1(n533_adj_4660), 
            .CO(n51073));
    SB_LUT4 add_6323_7_lut (.I0(GND_net), .I1(n17840[4]), .I2(n460_adj_4661), 
            .I3(n51071), .O(n17329[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_7 (.CI(n51071), .I0(n17840[4]), .I1(n460_adj_4661), 
            .CO(n51072));
    SB_LUT4 add_6323_6_lut (.I0(GND_net), .I1(n17840[3]), .I2(n387_adj_4662), 
            .I3(n51070), .O(n17329[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_6 (.CI(n51070), .I0(n17840[3]), .I1(n387_adj_4662), 
            .CO(n51071));
    SB_LUT4 add_6338_5_lut (.I0(GND_net), .I1(n18065[2]), .I2(n317), .I3(n49906), 
            .O(n17585[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_5_lut (.I0(GND_net), .I1(n17840[2]), .I2(n314_adj_4663), 
            .I3(n51069), .O(n17329[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_5 (.CI(n51069), .I0(n17840[2]), .I1(n314_adj_4663), 
            .CO(n51070));
    SB_CARRY add_6338_5 (.CI(n49906), .I0(n18065[2]), .I1(n317), .CO(n49907));
    SB_LUT4 add_6323_4_lut (.I0(GND_net), .I1(n17840[1]), .I2(n241_adj_4664), 
            .I3(n51068), .O(n17329[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_4 (.CI(n51068), .I0(n17840[1]), .I1(n241_adj_4664), 
            .CO(n51069));
    SB_LUT4 add_6323_3_lut (.I0(GND_net), .I1(n17840[0]), .I2(n168_adj_4665), 
            .I3(n51067), .O(n17329[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13751_3_lut (.I0(n356[23]), .I1(n436[23]), .I2(n11610), .I3(GND_net), 
            .O(n27817));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13751_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6323_3 (.CI(n51067), .I0(n17840[0]), .I1(n168_adj_4665), 
            .CO(n51068));
    SB_LUT4 i29327_4_lut (.I0(PWMLimit[23]), .I1(n60589), .I2(n27817), 
            .I3(n11608), .O(n49[23]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29327_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6323_2_lut (.I0(GND_net), .I1(n26_adj_4667), .I2(n95_adj_4668), 
            .I3(GND_net), .O(n17329[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_2 (.CI(GND_net), .I0(n26_adj_4667), .I1(n95_adj_4668), 
            .CO(n51067));
    SB_LUT4 add_6353_16_lut (.I0(GND_net), .I1(n18289[13]), .I2(n1120_adj_4669), 
            .I3(n51066), .O(n17840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6353_15_lut (.I0(GND_net), .I1(n18289[12]), .I2(n1047_adj_4670), 
            .I3(n51065), .O(n17840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_15 (.CI(n51065), .I0(n18289[12]), .I1(n1047_adj_4670), 
            .CO(n51066));
    SB_LUT4 add_6353_14_lut (.I0(GND_net), .I1(n18289[11]), .I2(n974_adj_4671), 
            .I3(n51064), .O(n17840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_14 (.CI(n51064), .I0(n18289[11]), .I1(n974_adj_4671), 
            .CO(n51065));
    SB_LUT4 add_6353_13_lut (.I0(GND_net), .I1(n18289[10]), .I2(n901_adj_4672), 
            .I3(n51063), .O(n17840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_13 (.CI(n51063), .I0(n18289[10]), .I1(n901_adj_4672), 
            .CO(n51064));
    SB_LUT4 add_6353_12_lut (.I0(GND_net), .I1(n18289[9]), .I2(n828_adj_4673), 
            .I3(n51062), .O(n17840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_12 (.CI(n51062), .I0(n18289[9]), .I1(n828_adj_4673), 
            .CO(n51063));
    SB_LUT4 add_6353_11_lut (.I0(GND_net), .I1(n18289[8]), .I2(n755_adj_4674), 
            .I3(n51061), .O(n17840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_11 (.CI(n51061), .I0(n18289[8]), .I1(n755_adj_4674), 
            .CO(n51062));
    SB_LUT4 add_6353_10_lut (.I0(GND_net), .I1(n18289[7]), .I2(n682_adj_4675), 
            .I3(n51060), .O(n17840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_10 (.CI(n51060), .I0(n18289[7]), .I1(n682_adj_4675), 
            .CO(n51061));
    SB_LUT4 add_6353_9_lut (.I0(GND_net), .I1(n18289[6]), .I2(n609_adj_4676), 
            .I3(n51059), .O(n17840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_9 (.CI(n51059), .I0(n18289[6]), .I1(n609_adj_4676), 
            .CO(n51060));
    SB_LUT4 add_6353_8_lut (.I0(GND_net), .I1(n18289[5]), .I2(n536_adj_4677), 
            .I3(n51058), .O(n17840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_8 (.CI(n51058), .I0(n18289[5]), .I1(n536_adj_4677), 
            .CO(n51059));
    SB_LUT4 add_6353_7_lut (.I0(GND_net), .I1(n18289[4]), .I2(n463_adj_4678), 
            .I3(n51057), .O(n17840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_7 (.CI(n51057), .I0(n18289[4]), .I1(n463_adj_4678), 
            .CO(n51058));
    SB_LUT4 add_6353_6_lut (.I0(GND_net), .I1(n18289[3]), .I2(n390_adj_4679), 
            .I3(n51056), .O(n17840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_6 (.CI(n51056), .I0(n18289[3]), .I1(n390_adj_4679), 
            .CO(n51057));
    SB_LUT4 add_6338_4_lut (.I0(GND_net), .I1(n18065[1]), .I2(n244), .I3(n49905), 
            .O(n17585[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6353_5_lut (.I0(GND_net), .I1(n18289[2]), .I2(n317_adj_4680), 
            .I3(n51055), .O(n17840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_5 (.CI(n51055), .I0(n18289[2]), .I1(n317_adj_4680), 
            .CO(n51056));
    SB_LUT4 add_6353_4_lut (.I0(GND_net), .I1(n18289[1]), .I2(n244_adj_4681), 
            .I3(n51054), .O(n17840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_4 (.CI(n49905), .I0(n18065[1]), .I1(n244), .CO(n49906));
    SB_CARRY add_6353_4 (.CI(n51054), .I0(n18289[1]), .I1(n244_adj_4681), 
            .CO(n51055));
    SB_LUT4 add_6353_3_lut (.I0(GND_net), .I1(n18289[0]), .I2(n171), .I3(n51053), 
            .O(n17840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_3 (.CI(n51053), .I0(n18289[0]), .I1(n171), .CO(n51054));
    SB_LUT4 add_6353_2_lut (.I0(GND_net), .I1(n29_adj_4682), .I2(n98), 
            .I3(GND_net), .O(n17840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_2 (.CI(GND_net), .I0(n29_adj_4682), .I1(n98), .CO(n51053));
    SB_LUT4 add_6514_8_lut (.I0(GND_net), .I1(n20081[5]), .I2(n560_adj_4683), 
            .I3(n51052), .O(n19969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6514_7_lut (.I0(GND_net), .I1(n20081[4]), .I2(n487_adj_4684), 
            .I3(n51051), .O(n19969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6514_7 (.CI(n51051), .I0(n20081[4]), .I1(n487_adj_4684), 
            .CO(n51052));
    SB_LUT4 i50177_4_lut (.I0(n33_adj_4564), .I1(n31_adj_4552), .I2(n29_adj_4551), 
            .I3(n65918), .O(n65905));
    defparam i50177_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6514_6_lut (.I0(GND_net), .I1(n20081[3]), .I2(n414_adj_4685), 
            .I3(n51050), .O(n19969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52721_4_lut (.I0(n30_adj_4573), .I1(n10_adj_4572), .I2(n35_adj_4565), 
            .I3(n65901), .O(n68449));   // verilog/motorControl.v(47[21:44])
    defparam i52721_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52171_3_lut (.I0(n68158), .I1(n182[15]), .I2(n31_adj_4552), 
            .I3(GND_net), .O(n67899));   // verilog/motorControl.v(47[21:44])
    defparam i52171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52846_4_lut (.I0(n67899), .I1(n68449), .I2(n35_adj_4565), 
            .I3(n65905), .O(n68574));   // verilog/motorControl.v(47[21:44])
    defparam i52846_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52847_3_lut (.I0(n68574), .I1(n182[18]), .I2(n37_adj_4566), 
            .I3(GND_net), .O(n68575));   // verilog/motorControl.v(47[21:44])
    defparam i52847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52814_3_lut (.I0(n68575), .I1(n182[19]), .I2(n39_adj_4548), 
            .I3(GND_net), .O(n68542));   // verilog/motorControl.v(47[21:44])
    defparam i52814_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6514_6 (.CI(n51050), .I0(n20081[3]), .I1(n414_adj_4685), 
            .CO(n51051));
    SB_LUT4 add_6514_5_lut (.I0(GND_net), .I1(n20081[2]), .I2(n341_adj_4686), 
            .I3(n51049), .O(n19969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6514_5 (.CI(n51049), .I0(n20081[2]), .I1(n341_adj_4686), 
            .CO(n51050));
    SB_LUT4 add_6514_4_lut (.I0(GND_net), .I1(n20081[1]), .I2(n268_adj_4687), 
            .I3(n51048), .O(n19969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6514_4 (.CI(n51048), .I0(n20081[1]), .I1(n268_adj_4687), 
            .CO(n51049));
    SB_LUT4 i50144_4_lut (.I0(n43_adj_4550), .I1(n41_adj_4547), .I2(n39_adj_4548), 
            .I3(n68396), .O(n65872));
    defparam i50144_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6514_3_lut (.I0(GND_net), .I1(n20081[0]), .I2(n195_adj_4688), 
            .I3(n51047), .O(n19969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6338_3_lut (.I0(GND_net), .I1(n18065[0]), .I2(n171_adj_4689), 
            .I3(n49904), .O(n17585[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6514_3 (.CI(n51047), .I0(n20081[0]), .I1(n195_adj_4688), 
            .CO(n51048));
    SB_CARRY add_6338_3 (.CI(n49904), .I0(n18065[0]), .I1(n171_adj_4689), 
            .CO(n49905));
    SB_LUT4 add_6514_2_lut (.I0(GND_net), .I1(n53_c), .I2(n122_adj_4690), 
            .I3(GND_net), .O(n19969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6514_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6514_2 (.CI(GND_net), .I0(n53_c), .I1(n122_adj_4690), 
            .CO(n51047));
    SB_LUT4 add_6381_15_lut (.I0(GND_net), .I1(n18680[12]), .I2(n1050_adj_4691), 
            .I3(n51046), .O(n18289[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6381_14_lut (.I0(GND_net), .I1(n18680[11]), .I2(n977_adj_4692), 
            .I3(n51045), .O(n18289[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_14 (.CI(n51045), .I0(n18680[11]), .I1(n977_adj_4692), 
            .CO(n51046));
    SB_LUT4 add_6381_13_lut (.I0(GND_net), .I1(n18680[10]), .I2(n904_adj_4693), 
            .I3(n51044), .O(n18289[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_13 (.CI(n51044), .I0(n18680[10]), .I1(n904_adj_4693), 
            .CO(n51045));
    SB_LUT4 add_6381_12_lut (.I0(GND_net), .I1(n18680[9]), .I2(n831_adj_4694), 
            .I3(n51043), .O(n18289[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52174_4_lut (.I0(n67897), .I1(n67580), .I2(n45_adj_4549), 
            .I3(n65870), .O(n67902));   // verilog/motorControl.v(47[21:44])
    defparam i52174_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52759_3_lut (.I0(n68542), .I1(n182[20]), .I2(n41_adj_4547), 
            .I3(GND_net), .O(n40_adj_4695));   // verilog/motorControl.v(47[21:44])
    defparam i52759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52479_4_lut (.I0(n40_adj_4695), .I1(n67902), .I2(n45_adj_4549), 
            .I3(n65872), .O(n68207));   // verilog/motorControl.v(47[21:44])
    defparam i52479_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_6381_12 (.CI(n51043), .I0(n18680[9]), .I1(n831_adj_4694), 
            .CO(n51044));
    SB_LUT4 i52480_3_lut (.I0(n68207), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(47[21:44])
    defparam i52480_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6381_11_lut (.I0(GND_net), .I1(n18680[8]), .I2(n758), 
            .I3(n51042), .O(n18289[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_11 (.CI(n51042), .I0(n18680[8]), .I1(n758), .CO(n51043));
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[14] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6338_2_lut (.I0(GND_net), .I1(n29_adj_4696), .I2(n98_adj_4697), 
            .I3(GND_net), .O(n17585[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6338_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6381_10_lut (.I0(GND_net), .I1(n18680[7]), .I2(n685), 
            .I3(n51041), .O(n18289[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6338_2 (.CI(GND_net), .I0(n29_adj_4696), .I1(n98_adj_4697), 
            .CO(n49904));
    SB_CARRY add_6381_10 (.CI(n51041), .I0(n18680[7]), .I1(n685), .CO(n51042));
    SB_LUT4 add_6381_9_lut (.I0(GND_net), .I1(n18680[6]), .I2(n612), .I3(n51040), 
            .O(n18289[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_9 (.CI(n51040), .I0(n18680[6]), .I1(n612), .CO(n51041));
    SB_LUT4 add_6381_8_lut (.I0(GND_net), .I1(n18680[5]), .I2(n539), .I3(n51039), 
            .O(n18289[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_8 (.CI(n51039), .I0(n18680[5]), .I1(n539), .CO(n51040));
    SB_LUT4 add_6381_7_lut (.I0(GND_net), .I1(n18680[4]), .I2(n466), .I3(n51038), 
            .O(n18289[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_7 (.CI(n51038), .I0(n18680[4]), .I1(n466), .CO(n51039));
    SB_LUT4 add_6381_6_lut (.I0(GND_net), .I1(n18680[3]), .I2(n393_adj_4698), 
            .I3(n51037), .O(n18289[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_6 (.CI(n51037), .I0(n18680[3]), .I1(n393_adj_4698), 
            .CO(n51038));
    SB_LUT4 add_6381_5_lut (.I0(GND_net), .I1(n18680[2]), .I2(n320), .I3(n51036), 
            .O(n18289[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_5 (.CI(n51036), .I0(n18680[2]), .I1(n320), .CO(n51037));
    SB_CARRY add_9_24 (.CI(n49603), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n1[22]), .CO(n49604));
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n1[21]), .I3(n49602), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6381_4_lut (.I0(GND_net), .I1(n18680[1]), .I2(n247), .I3(n51035), 
            .O(n18289[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_4 (.CI(n51035), .I0(n18680[1]), .I1(n247), .CO(n51036));
    SB_LUT4 add_6381_3_lut (.I0(GND_net), .I1(n18680[0]), .I2(n174), .I3(n51034), 
            .O(n18289[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_3 (.CI(n51034), .I0(n18680[0]), .I1(n174), .CO(n51035));
    SB_LUT4 add_6381_2_lut (.I0(GND_net), .I1(n32_adj_4699), .I2(n101), 
            .I3(GND_net), .O(n18289[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_2 (.CI(GND_net), .I0(n32_adj_4699), .I1(n101), .CO(n51034));
    SB_LUT4 add_6407_14_lut (.I0(GND_net), .I1(n19017[11]), .I2(n980_adj_4700), 
            .I3(n51033), .O(n18680[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_13_lut (.I0(GND_net), .I1(n19017[10]), .I2(n907_adj_4701), 
            .I3(n51032), .O(n18680[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_13 (.CI(n51032), .I0(n19017[10]), .I1(n907_adj_4701), 
            .CO(n51033));
    SB_LUT4 add_6407_12_lut (.I0(GND_net), .I1(n19017[9]), .I2(n834_adj_4702), 
            .I3(n51031), .O(n18680[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_23_lut (.I0(GND_net), .I1(n13220[20]), .I2(GND_net), 
            .I3(n50148), .O(n12157[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_12 (.CI(n51031), .I0(n19017[9]), .I1(n834_adj_4702), 
            .CO(n51032));
    SB_LUT4 add_6407_11_lut (.I0(GND_net), .I1(n19017[8]), .I2(n761_adj_4703), 
            .I3(n51030), .O(n18680[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_11 (.CI(n51030), .I0(n19017[8]), .I1(n761_adj_4703), 
            .CO(n51031));
    SB_LUT4 add_6407_10_lut (.I0(GND_net), .I1(n19017[7]), .I2(n688_adj_4704), 
            .I3(n51029), .O(n18680[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_10 (.CI(n51029), .I0(n19017[7]), .I1(n688_adj_4704), 
            .CO(n51030));
    SB_LUT4 add_6407_9_lut (.I0(GND_net), .I1(n19017[6]), .I2(n615), .I3(n51028), 
            .O(n18680[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_22_lut (.I0(GND_net), .I1(n13220[19]), .I2(GND_net), 
            .I3(n50147), .O(n12157[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_9 (.CI(n51028), .I0(n19017[6]), .I1(n615), .CO(n51029));
    SB_CARRY add_6052_22 (.CI(n50147), .I0(n13220[19]), .I1(GND_net), 
            .CO(n50148));
    SB_LUT4 add_6407_8_lut (.I0(GND_net), .I1(n19017[5]), .I2(n542), .I3(n51027), 
            .O(n18680[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_8 (.CI(n51027), .I0(n19017[5]), .I1(n542), .CO(n51028));
    SB_LUT4 add_6407_7_lut (.I0(GND_net), .I1(n19017[4]), .I2(n469), .I3(n51026), 
            .O(n18680[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_7 (.CI(n51026), .I0(n19017[4]), .I1(n469), .CO(n51027));
    SB_LUT4 add_6052_21_lut (.I0(GND_net), .I1(n13220[18]), .I2(GND_net), 
            .I3(n50146), .O(n12157[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_6_lut (.I0(GND_net), .I1(n19017[3]), .I2(n396_adj_4705), 
            .I3(n51025), .O(n18680[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_21 (.CI(n50146), .I0(n13220[18]), .I1(GND_net), 
            .CO(n50147));
    SB_LUT4 add_6052_20_lut (.I0(GND_net), .I1(n13220[17]), .I2(GND_net), 
            .I3(n50145), .O(n12157[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_20 (.CI(n50145), .I0(n13220[17]), .I1(GND_net), 
            .CO(n50146));
    SB_CARRY add_6407_6 (.CI(n51025), .I0(n19017[3]), .I1(n396_adj_4705), 
            .CO(n51026));
    SB_LUT4 add_6052_19_lut (.I0(GND_net), .I1(n13220[16]), .I2(GND_net), 
            .I3(n50144), .O(n12157[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_5_lut (.I0(GND_net), .I1(n19017[2]), .I2(n323), .I3(n51024), 
            .O(n18680[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_5 (.CI(n51024), .I0(n19017[2]), .I1(n323), .CO(n51025));
    SB_CARRY add_6052_19 (.CI(n50144), .I0(n13220[16]), .I1(GND_net), 
            .CO(n50145));
    SB_LUT4 add_6407_4_lut (.I0(GND_net), .I1(n19017[1]), .I2(n250), .I3(n51023), 
            .O(n18680[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_4 (.CI(n51023), .I0(n19017[1]), .I1(n250), .CO(n51024));
    SB_LUT4 add_6407_3_lut (.I0(GND_net), .I1(n19017[0]), .I2(n177), .I3(n51022), 
            .O(n18680[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_3 (.CI(n51022), .I0(n19017[0]), .I1(n177), .CO(n51023));
    SB_LUT4 add_6052_18_lut (.I0(GND_net), .I1(n13220[15]), .I2(GND_net), 
            .I3(n50143), .O(n12157[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_2_lut (.I0(GND_net), .I1(n35_adj_4706), .I2(n104), 
            .I3(GND_net), .O(n18680[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_2 (.CI(GND_net), .I0(n35_adj_4706), .I1(n104), .CO(n51022));
    SB_CARRY add_6052_18 (.CI(n50143), .I0(n13220[15]), .I1(GND_net), 
            .CO(n50144));
    SB_LUT4 add_6527_7_lut (.I0(GND_net), .I1(n59281), .I2(n490_c), .I3(n51021), 
            .O(n20081[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6527_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_17_lut (.I0(GND_net), .I1(n13220[14]), .I2(GND_net), 
            .I3(n50142), .O(n12157[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6527_6_lut (.I0(GND_net), .I1(n20165[3]), .I2(n417_c), 
            .I3(n51020), .O(n20081[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6527_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6527_6 (.CI(n51020), .I0(n20165[3]), .I1(n417_c), .CO(n51021));
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[10]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6527_5_lut (.I0(GND_net), .I1(n20165[2]), .I2(n344_adj_4707), 
            .I3(n51019), .O(n20081[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6527_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[11]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6527_5 (.CI(n51019), .I0(n20165[2]), .I1(n344_adj_4707), 
            .CO(n51020));
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[12]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6527_4_lut (.I0(GND_net), .I1(n20165[1]), .I2(n271_c), 
            .I3(n51018), .O(n20081[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6527_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6527_4 (.CI(n51018), .I0(n20165[1]), .I1(n271_c), .CO(n51019));
    SB_LUT4 add_6527_3_lut (.I0(GND_net), .I1(n20165[0]), .I2(n198_adj_4708), 
            .I3(n51017), .O(n20081[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6527_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6527_3 (.CI(n51017), .I0(n20165[0]), .I1(n198_adj_4708), 
            .CO(n51018));
    SB_LUT4 add_6527_2_lut (.I0(GND_net), .I1(n56_adj_4709), .I2(n125_adj_4710), 
            .I3(GND_net), .O(n20081[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6527_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6527_2 (.CI(GND_net), .I0(n56_adj_4709), .I1(n125_adj_4710), 
            .CO(n51017));
    SB_LUT4 add_6431_13_lut (.I0(GND_net), .I1(n19304[10]), .I2(n910), 
            .I3(n51016), .O(n19017[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6431_12_lut (.I0(GND_net), .I1(n19304[9]), .I2(n837), 
            .I3(n51015), .O(n19017[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_12 (.CI(n51015), .I0(n19304[9]), .I1(n837), .CO(n51016));
    SB_LUT4 add_6431_11_lut (.I0(GND_net), .I1(n19304[8]), .I2(n764), 
            .I3(n51014), .O(n19017[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_11 (.CI(n51014), .I0(n19304[8]), .I1(n764), .CO(n51015));
    SB_LUT4 add_6431_10_lut (.I0(GND_net), .I1(n19304[7]), .I2(n691), 
            .I3(n51013), .O(n19017[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_10 (.CI(n51013), .I0(n19304[7]), .I1(n691), .CO(n51014));
    SB_LUT4 add_6431_9_lut (.I0(GND_net), .I1(n19304[6]), .I2(n618), .I3(n51012), 
            .O(n19017[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_9 (.CI(n51012), .I0(n19304[6]), .I1(n618), .CO(n51013));
    SB_CARRY add_6052_17 (.CI(n50142), .I0(n13220[14]), .I1(GND_net), 
            .CO(n50143));
    SB_LUT4 add_6431_8_lut (.I0(GND_net), .I1(n19304[5]), .I2(n545), .I3(n51011), 
            .O(n19017[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_16_lut (.I0(GND_net), .I1(n13220[13]), .I2(n1099_adj_4711), 
            .I3(n50141), .O(n12157[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_8 (.CI(n51011), .I0(n19304[5]), .I1(n545), .CO(n51012));
    SB_LUT4 add_6431_7_lut (.I0(GND_net), .I1(n19304[4]), .I2(n472), .I3(n51010), 
            .O(n19017[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n49602), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n1[21]), .CO(n49603));
    SB_CARRY add_6052_16 (.CI(n50141), .I0(n13220[13]), .I1(n1099_adj_4711), 
            .CO(n50142));
    SB_CARRY add_6431_7 (.CI(n51010), .I0(n19304[4]), .I1(n472), .CO(n51011));
    SB_LUT4 add_6052_15_lut (.I0(GND_net), .I1(n13220[12]), .I2(n1026_adj_4712), 
            .I3(n50140), .O(n12157[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6431_6_lut (.I0(GND_net), .I1(n19304[3]), .I2(n399), .I3(n51009), 
            .O(n19017[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_15 (.CI(n50140), .I0(n13220[12]), .I1(n1026_adj_4712), 
            .CO(n50141));
    SB_CARRY add_6431_6 (.CI(n51009), .I0(n19304[3]), .I1(n399), .CO(n51010));
    SB_LUT4 add_6431_5_lut (.I0(GND_net), .I1(n19304[2]), .I2(n326), .I3(n51008), 
            .O(n19017[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_5 (.CI(n51008), .I0(n19304[2]), .I1(n326), .CO(n51009));
    SB_LUT4 add_6431_4_lut (.I0(GND_net), .I1(n19304[1]), .I2(n253), .I3(n51007), 
            .O(n19017[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_14_lut (.I0(GND_net), .I1(n13220[11]), .I2(n953_adj_4713), 
            .I3(n50139), .O(n12157[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_4 (.CI(n51007), .I0(n19304[1]), .I1(n253), .CO(n51008));
    SB_LUT4 add_6431_3_lut (.I0(GND_net), .I1(n19304[0]), .I2(n180), .I3(n51006), 
            .O(n19017[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_3 (.CI(n51006), .I0(n19304[0]), .I1(n180), .CO(n51007));
    SB_LUT4 add_6431_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_4715), 
            .I3(GND_net), .O(n19017[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_4715), .CO(n51006));
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[13]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6453_12_lut (.I0(GND_net), .I1(n19545[9]), .I2(n840), 
            .I3(n51005), .O(n19304[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6453_11_lut (.I0(GND_net), .I1(n19545[8]), .I2(n767_adj_4716), 
            .I3(n51004), .O(n19304[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_11 (.CI(n51004), .I0(n19545[8]), .I1(n767_adj_4716), 
            .CO(n51005));
    SB_LUT4 add_6453_10_lut (.I0(GND_net), .I1(n19545[7]), .I2(n694_adj_4717), 
            .I3(n51003), .O(n19304[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_10 (.CI(n51003), .I0(n19545[7]), .I1(n694_adj_4717), 
            .CO(n51004));
    SB_LUT4 add_6453_9_lut (.I0(GND_net), .I1(n19545[6]), .I2(n621_adj_4718), 
            .I3(n51002), .O(n19304[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_9 (.CI(n51002), .I0(n19545[6]), .I1(n621_adj_4718), 
            .CO(n51003));
    SB_LUT4 add_6453_8_lut (.I0(GND_net), .I1(n19545[5]), .I2(n548_adj_4719), 
            .I3(n51001), .O(n19304[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_8 (.CI(n51001), .I0(n19545[5]), .I1(n548_adj_4719), 
            .CO(n51002));
    SB_LUT4 add_6453_7_lut (.I0(GND_net), .I1(n19545[4]), .I2(n475_adj_4720), 
            .I3(n51000), .O(n19304[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_7 (.CI(n51000), .I0(n19545[4]), .I1(n475_adj_4720), 
            .CO(n51001));
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29669), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_6453_6_lut (.I0(GND_net), .I1(n19545[3]), .I2(n402_adj_4721), 
            .I3(n50999), .O(n19304[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_6 (.CI(n50999), .I0(n19545[3]), .I1(n402_adj_4721), 
            .CO(n51000));
    SB_LUT4 add_6453_5_lut (.I0(GND_net), .I1(n19545[2]), .I2(n329_adj_4722), 
            .I3(n50998), .O(n19304[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_5 (.CI(n50998), .I0(n19545[2]), .I1(n329_adj_4722), 
            .CO(n50999));
    SB_LUT4 add_6453_4_lut (.I0(GND_net), .I1(n19545[1]), .I2(n256_adj_4723), 
            .I3(n50997), .O(n19304[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_4 (.CI(n50997), .I0(n19545[1]), .I1(n256_adj_4723), 
            .CO(n50998));
    SB_LUT4 add_6453_3_lut (.I0(GND_net), .I1(n19545[0]), .I2(n183_adj_4724), 
            .I3(n50996), .O(n19304[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_3 (.CI(n50996), .I0(n19545[0]), .I1(n183_adj_4724), 
            .CO(n50997));
    SB_LUT4 add_6453_2_lut (.I0(GND_net), .I1(n41_adj_4725), .I2(n110), 
            .I3(GND_net), .O(n19304[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_2 (.CI(GND_net), .I0(n41_adj_4725), .I1(n110), .CO(n50996));
    SB_CARRY add_6052_14 (.CI(n50139), .I0(n13220[11]), .I1(n953_adj_4713), 
            .CO(n50140));
    SB_LUT4 add_6052_13_lut (.I0(GND_net), .I1(n13220[10]), .I2(n880_adj_4727), 
            .I3(n50138), .O(n12157[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n1[20]), .I3(n49601), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1943__i0 (.Q(counter[0]), .C(clk16MHz), .D(n51[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i31 (.Q(counter[31]), .C(clk16MHz), .D(n51[31]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i30 (.Q(counter[30]), .C(clk16MHz), .D(n51[30]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i29 (.Q(counter[29]), .C(clk16MHz), .D(n51[29]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i28 (.Q(counter[28]), .C(clk16MHz), .D(n51[28]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i27 (.Q(counter[27]), .C(clk16MHz), .D(n51[27]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i26 (.Q(counter[26]), .C(clk16MHz), .D(n51[26]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i25 (.Q(counter[25]), .C(clk16MHz), .D(n51[25]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i24 (.Q(counter[24]), .C(clk16MHz), .D(n51[24]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i23 (.Q(counter[23]), .C(clk16MHz), .D(n51[23]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i22 (.Q(counter[22]), .C(clk16MHz), .D(n51[22]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i21 (.Q(counter[21]), .C(clk16MHz), .D(n51[21]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i20 (.Q(counter[20]), .C(clk16MHz), .D(n51[20]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i19 (.Q(counter[19]), .C(clk16MHz), .D(n51[19]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i18 (.Q(counter[18]), .C(clk16MHz), .D(n51[18]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i17 (.Q(counter[17]), .C(clk16MHz), .D(n51[17]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i16 (.Q(counter[16]), .C(clk16MHz), .D(n51[16]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i15 (.Q(counter[15]), .C(clk16MHz), .D(n51[15]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i14 (.Q(counter[14]), .C(clk16MHz), .D(n51[14]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i13 (.Q(counter[13]), .C(clk16MHz), .D(n51[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i12 (.Q(counter[12]), .C(clk16MHz), .D(n51[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i11 (.Q(counter[11]), .C(clk16MHz), .D(n51[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i10 (.Q(counter[10]), .C(clk16MHz), .D(n51[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i9 (.Q(counter[9]), .C(clk16MHz), .D(n51[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i8 (.Q(counter[8]), .C(clk16MHz), .D(n51[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i7 (.Q(counter[7]), .C(clk16MHz), .D(n51[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i6 (.Q(counter[6]), .C(clk16MHz), .D(n51[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i5 (.Q(counter[5]), .C(clk16MHz), .D(n51[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i4 (.Q(counter[4]), .C(clk16MHz), .D(n51[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i3 (.Q(counter[3]), .C(clk16MHz), .D(n51[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i2 (.Q(counter[2]), .C(clk16MHz), .D(n51[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i1 (.Q(counter[1]), .C(clk16MHz), .D(n51[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFER result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n49[23]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY add_6052_13 (.CI(n50138), .I0(n13220[10]), .I1(n880_adj_4727), 
            .CO(n50139));
    SB_LUT4 add_6367_15_lut (.I0(GND_net), .I1(n18485[12]), .I2(n1050), 
            .I3(n49893), .O(n18065[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_22 (.CI(n49601), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n1[20]), .CO(n49602));
    SB_LUT4 add_6367_14_lut (.I0(GND_net), .I1(n18485[11]), .I2(n977), 
            .I3(n49892), .O(n18065[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n1[19]), .I3(n49600), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_12_lut (.I0(GND_net), .I1(n13220[9]), .I2(n807_adj_4597), 
            .I3(n50137), .O(n12157[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1943_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n50869), .O(n51[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1943_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n50868), .O(n51[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_32 (.CI(n50868), .I0(GND_net), .I1(counter[30]), 
            .CO(n50869));
    SB_LUT4 counter_1943_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n50867), .O(n51[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_31 (.CI(n50867), .I0(GND_net), .I1(counter[29]), 
            .CO(n50868));
    SB_LUT4 counter_1943_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n50866), .O(n51[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_30 (.CI(n50866), .I0(GND_net), .I1(counter[28]), 
            .CO(n50867));
    SB_DFFER result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n49[22]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 counter_1943_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n50865), .O(n51[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_29 (.CI(n50865), .I0(GND_net), .I1(counter[27]), 
            .CO(n50866));
    SB_LUT4 counter_1943_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n50864), .O(n51[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_28 (.CI(n50864), .I0(GND_net), .I1(counter[26]), 
            .CO(n50865));
    SB_LUT4 counter_1943_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n50863), .O(n51[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_27 (.CI(n50863), .I0(GND_net), .I1(counter[25]), 
            .CO(n50864));
    SB_LUT4 counter_1943_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n50862), .O(n51[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4462));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_1943_add_4_26 (.CI(n50862), .I0(GND_net), .I1(counter[24]), 
            .CO(n50863));
    SB_LUT4 counter_1943_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n50861), .O(n51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_25 (.CI(n50861), .I0(GND_net), .I1(counter[23]), 
            .CO(n50862));
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_1943_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n50860), .O(n51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_24 (.CI(n50860), .I0(GND_net), .I1(counter[22]), 
            .CO(n50861));
    SB_LUT4 counter_1943_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n50859), .O(n51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_23 (.CI(n50859), .I0(GND_net), .I1(counter[21]), 
            .CO(n50860));
    SB_LUT4 counter_1943_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n50858), .O(n51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n49[21]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_CARRY counter_1943_add_4_22 (.CI(n50858), .I0(GND_net), .I1(counter[20]), 
            .CO(n50859));
    SB_LUT4 counter_1943_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n50857), .O(n51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_21 (.CI(n50857), .I0(GND_net), .I1(counter[19]), 
            .CO(n50858));
    SB_DFFER result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n49[20]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n49[19]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 counter_1943_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n50856), .O(n51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_20 (.CI(n50856), .I0(GND_net), .I1(counter[18]), 
            .CO(n50857));
    SB_CARRY add_6367_14 (.CI(n49892), .I0(n18485[11]), .I1(n977), .CO(n49893));
    SB_LUT4 counter_1943_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n50855), .O(n51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_19 (.CI(n50855), .I0(GND_net), .I1(counter[17]), 
            .CO(n50856));
    SB_LUT4 counter_1943_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n50854), .O(n51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_18 (.CI(n50854), .I0(GND_net), .I1(counter[16]), 
            .CO(n50855));
    SB_LUT4 counter_1943_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n50853), .O(n51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_17 (.CI(n50853), .I0(GND_net), .I1(counter[15]), 
            .CO(n50854));
    SB_LUT4 counter_1943_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n50852), .O(n51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_16 (.CI(n50852), .I0(GND_net), .I1(counter[14]), 
            .CO(n50853));
    SB_LUT4 counter_1943_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n50851), .O(n51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_15 (.CI(n50851), .I0(GND_net), .I1(counter[13]), 
            .CO(n50852));
    SB_LUT4 counter_1943_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n50850), .O(n51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_14 (.CI(n50850), .I0(GND_net), .I1(counter[12]), 
            .CO(n50851));
    SB_LUT4 counter_1943_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n50849), .O(n51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_13 (.CI(n50849), .I0(GND_net), .I1(counter[11]), 
            .CO(n50850));
    SB_LUT4 counter_1943_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n50848), .O(n51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_12 (.CI(n50848), .I0(GND_net), .I1(counter[10]), 
            .CO(n50849));
    SB_LUT4 counter_1943_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n50847), .O(n51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_11 (.CI(n50847), .I0(GND_net), .I1(counter[9]), 
            .CO(n50848));
    SB_LUT4 counter_1943_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n50846), .O(n51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_10 (.CI(n50846), .I0(GND_net), .I1(counter[8]), 
            .CO(n50847));
    SB_LUT4 counter_1943_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n50845), .O(n51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_9 (.CI(n50845), .I0(GND_net), .I1(counter[7]), 
            .CO(n50846));
    SB_LUT4 counter_1943_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n50844), .O(n51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_8 (.CI(n50844), .I0(GND_net), .I1(counter[6]), 
            .CO(n50845));
    SB_LUT4 counter_1943_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n50843), .O(n51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_7 (.CI(n50843), .I0(GND_net), .I1(counter[5]), 
            .CO(n50844));
    SB_LUT4 counter_1943_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n50842), .O(n51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_6 (.CI(n50842), .I0(GND_net), .I1(counter[4]), 
            .CO(n50843));
    SB_DFFER result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n49[18]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 counter_1943_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n50841), .O(n51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_5 (.CI(n50841), .I0(GND_net), .I1(counter[3]), 
            .CO(n50842));
    SB_DFFER result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n49[17]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 counter_1943_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n50840), .O(n51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_4 (.CI(n50840), .I0(GND_net), .I1(counter[2]), 
            .CO(n50841));
    SB_LUT4 counter_1943_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n50839), .O(n51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_3 (.CI(n50839), .I0(GND_net), .I1(counter[1]), 
            .CO(n50840));
    SB_LUT4 counter_1943_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n50839));
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[14]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_DFFER result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n49[16]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n49[15]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n49[14]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n49[13]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n49[12]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n49[11]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n49[10]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4727));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n49[9]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n49[8]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n49[7]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n49[6]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n49[5]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n49[4]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n49[3]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n49[2]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30497), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n30496), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n30495), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n30494), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n30493), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n30491), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n49[1]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n30489), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n30488), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n30487), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n30486), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30485), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30484), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30483), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30482), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30481), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30480), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30479), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30478), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30477), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30476), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30475), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30474), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30473), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 add_6367_13_lut (.I0(GND_net), .I1(n18485[10]), .I2(n904), 
            .I3(n49891), .O(n18065[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6367_13 (.CI(n49891), .I0(n18485[10]), .I1(n904), .CO(n49892));
    SB_LUT4 add_6367_12_lut (.I0(GND_net), .I1(n18485[9]), .I2(n831), 
            .I3(n49890), .O(n18065[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6367_12 (.CI(n49890), .I0(n18485[9]), .I1(n831), .CO(n49891));
    SB_CARRY add_6052_12 (.CI(n50137), .I0(n13220[9]), .I1(n807_adj_4597), 
            .CO(n50138));
    SB_LUT4 add_6052_11_lut (.I0(GND_net), .I1(n13220[8]), .I2(n734), 
            .I3(n50136), .O(n12157[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_11 (.CI(n50136), .I0(n13220[8]), .I1(n734), .CO(n50137));
    SB_LUT4 add_6367_11_lut (.I0(GND_net), .I1(n18485[8]), .I2(n758_adj_4753), 
            .I3(n49889), .O(n18065[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_10_lut (.I0(GND_net), .I1(n13220[7]), .I2(n661_adj_4754), 
            .I3(n50135), .O(n12157[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_10 (.CI(n50135), .I0(n13220[7]), .I1(n661_adj_4754), 
            .CO(n50136));
    SB_LUT4 add_6052_9_lut (.I0(GND_net), .I1(n13220[6]), .I2(n588_adj_4755), 
            .I3(n50134), .O(n12157[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_21 (.CI(n49600), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n1[19]), .CO(n49601));
    SB_CARRY add_6052_9 (.CI(n50134), .I0(n13220[6]), .I1(n588_adj_4755), 
            .CO(n50135));
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[15]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6052_8_lut (.I0(GND_net), .I1(n13220[5]), .I2(n515_adj_4756), 
            .I3(n50133), .O(n12157[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[23]), 
            .I3(n49743), .O(n436[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_8 (.CI(n50133), .I0(n13220[5]), .I1(n515_adj_4756), 
            .CO(n50134));
    SB_LUT4 add_6052_7_lut (.I0(GND_net), .I1(n13220[4]), .I2(n442_adj_4757), 
            .I3(n50132), .O(n12157[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_7 (.CI(n50132), .I0(n13220[4]), .I1(n442_adj_4757), 
            .CO(n50133));
    SB_CARRY add_6367_11 (.CI(n49889), .I0(n18485[8]), .I1(n758_adj_4753), 
            .CO(n49890));
    SB_LUT4 add_6367_10_lut (.I0(GND_net), .I1(n18485[7]), .I2(n685_adj_4758), 
            .I3(n49888), .O(n18065[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6367_10 (.CI(n49888), .I0(n18485[7]), .I1(n685_adj_4758), 
            .CO(n49889));
    SB_LUT4 add_6052_6_lut (.I0(GND_net), .I1(n13220[3]), .I2(n369_adj_4759), 
            .I3(n50131), .O(n12157[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[22]), 
            .I3(n49742), .O(n436[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_6 (.CI(n50131), .I0(n13220[3]), .I1(n369_adj_4759), 
            .CO(n50132));
    SB_LUT4 add_6367_9_lut (.I0(GND_net), .I1(n18485[6]), .I2(n612_adj_4760), 
            .I3(n49887), .O(n18065[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6052_5_lut (.I0(GND_net), .I1(n13220[2]), .I2(n296_adj_4761), 
            .I3(n50130), .O(n12157[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_5 (.CI(n50130), .I0(n13220[2]), .I1(n296_adj_4761), 
            .CO(n50131));
    SB_CARRY unary_minus_26_add_3_24 (.CI(n49742), .I0(GND_net), .I1(n1_adj_4985[22]), 
            .CO(n49743));
    SB_CARRY add_6367_9 (.CI(n49887), .I0(n18485[6]), .I1(n612_adj_4760), 
            .CO(n49888));
    SB_LUT4 add_6052_4_lut (.I0(GND_net), .I1(n13220[1]), .I2(n223_adj_4762), 
            .I3(n50129), .O(n12157[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n1[18]), .I3(n49599), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_4 (.CI(n50129), .I0(n13220[1]), .I1(n223_adj_4762), 
            .CO(n50130));
    SB_LUT4 add_6052_3_lut (.I0(GND_net), .I1(n13220[0]), .I2(n150_adj_4763), 
            .I3(n50128), .O(n12157[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_3 (.CI(n50128), .I0(n13220[0]), .I1(n150_adj_4763), 
            .CO(n50129));
    SB_LUT4 add_6052_2_lut (.I0(GND_net), .I1(n8_adj_4764), .I2(n77_adj_4765), 
            .I3(GND_net), .O(n12157[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6052_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[21]), 
            .I3(n49741), .O(n436[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_23 (.CI(n49741), .I0(GND_net), .I1(n1_adj_4985[21]), 
            .CO(n49742));
    SB_LUT4 add_6367_8_lut (.I0(GND_net), .I1(n18485[5]), .I2(n539_adj_4767), 
            .I3(n49886), .O(n18065[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6052_2 (.CI(GND_net), .I0(n8_adj_4764), .I1(n77_adj_4765), 
            .CO(n50128));
    SB_LUT4 add_6121_22_lut (.I0(GND_net), .I1(n14145[19]), .I2(GND_net), 
            .I3(n50127), .O(n13220[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6367_8 (.CI(n49886), .I0(n18485[5]), .I1(n539_adj_4767), 
            .CO(n49887));
    SB_LUT4 add_6367_7_lut (.I0(GND_net), .I1(n18485[4]), .I2(n466_adj_4768), 
            .I3(n49885), .O(n18065[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_21_lut (.I0(GND_net), .I1(n14145[18]), .I2(GND_net), 
            .I3(n50126), .O(n13220[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_21 (.CI(n50126), .I0(n14145[18]), .I1(GND_net), 
            .CO(n50127));
    SB_CARRY add_6367_7 (.CI(n49885), .I0(n18485[4]), .I1(n466_adj_4768), 
            .CO(n49886));
    SB_LUT4 add_6121_20_lut (.I0(GND_net), .I1(n14145[17]), .I2(GND_net), 
            .I3(n50125), .O(n13220[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6367_6_lut (.I0(GND_net), .I1(n18485[3]), .I2(n393_adj_4769), 
            .I3(n49884), .O(n18065[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_20 (.CI(n50125), .I0(n14145[17]), .I1(GND_net), 
            .CO(n50126));
    SB_LUT4 add_6121_19_lut (.I0(GND_net), .I1(n14145[16]), .I2(GND_net), 
            .I3(n50124), .O(n13220[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[16]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6121_19 (.CI(n50124), .I0(n14145[16]), .I1(GND_net), 
            .CO(n50125));
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[20]), 
            .I3(n49740), .O(n436[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_22 (.CI(n49740), .I0(GND_net), .I1(n1_adj_4985[20]), 
            .CO(n49741));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[19]), 
            .I3(n49739), .O(n436[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_18_lut (.I0(GND_net), .I1(n14145[15]), .I2(GND_net), 
            .I3(n50123), .O(n13220[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_18 (.CI(n50123), .I0(n14145[15]), .I1(GND_net), 
            .CO(n50124));
    SB_LUT4 add_6121_17_lut (.I0(GND_net), .I1(n14145[14]), .I2(GND_net), 
            .I3(n50122), .O(n13220[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[13] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6121_17 (.CI(n50122), .I0(n14145[14]), .I1(GND_net), 
            .CO(n50123));
    SB_LUT4 add_6121_16_lut (.I0(GND_net), .I1(n14145[13]), .I2(n1102_adj_4772), 
            .I3(n50121), .O(n13220[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_21 (.CI(n49739), .I0(GND_net), .I1(n1_adj_4985[19]), 
            .CO(n49740));
    SB_CARRY add_6121_16 (.CI(n50121), .I0(n14145[13]), .I1(n1102_adj_4772), 
            .CO(n50122));
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4725));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4724));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6121_15_lut (.I0(GND_net), .I1(n14145[12]), .I2(n1029_adj_4773), 
            .I3(n50120), .O(n13220[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_20 (.CI(n49599), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n1[18]), .CO(n49600));
    SB_CARRY add_6121_15 (.CI(n50120), .I0(n14145[12]), .I1(n1029_adj_4773), 
            .CO(n50121));
    SB_CARRY add_6367_6 (.CI(n49884), .I0(n18485[3]), .I1(n393_adj_4769), 
            .CO(n49885));
    SB_LUT4 add_6121_14_lut (.I0(GND_net), .I1(n14145[11]), .I2(n956_adj_4774), 
            .I3(n50119), .O(n13220[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_14 (.CI(n50119), .I0(n14145[11]), .I1(n956_adj_4774), 
            .CO(n50120));
    SB_LUT4 i28890_4_lut (.I0(PWMLimit[0]), .I1(n60589), .I2(n27722), 
            .I3(n11608), .O(n49[0]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i28890_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6121_13_lut (.I0(GND_net), .I1(n14145[10]), .I2(n883_adj_4775), 
            .I3(n50118), .O(n13220[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_13 (.CI(n50118), .I0(n14145[10]), .I1(n883_adj_4775), 
            .CO(n50119));
    SB_LUT4 add_6121_12_lut (.I0(GND_net), .I1(n14145[9]), .I2(n810_adj_4776), 
            .I3(n50117), .O(n13220[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6367_5_lut (.I0(GND_net), .I1(n18485[2]), .I2(n320_adj_4777), 
            .I3(n49883), .O(n18065[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_12 (.CI(n50117), .I0(n14145[9]), .I1(n810_adj_4776), 
            .CO(n50118));
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[18]), 
            .I3(n49738), .O(n436[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_11_lut (.I0(GND_net), .I1(n14145[8]), .I2(n737_adj_4779), 
            .I3(n50116), .O(n13220[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_11 (.CI(n50116), .I0(n14145[8]), .I1(n737_adj_4779), 
            .CO(n50117));
    SB_CARRY unary_minus_26_add_3_20 (.CI(n49738), .I0(GND_net), .I1(n1_adj_4985[18]), 
            .CO(n49739));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n1[17]), .I3(n49598), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_10_lut (.I0(GND_net), .I1(n14145[7]), .I2(n664_adj_4780), 
            .I3(n50115), .O(n13220[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_10 (.CI(n50115), .I0(n14145[7]), .I1(n664_adj_4780), 
            .CO(n50116));
    SB_LUT4 add_6121_9_lut (.I0(GND_net), .I1(n14145[6]), .I2(n591_adj_4781), 
            .I3(n50114), .O(n13220[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[17]), 
            .I3(n49737), .O(n436[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_9 (.CI(n50114), .I0(n14145[6]), .I1(n591_adj_4781), 
            .CO(n50115));
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4723));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4722));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6121_8_lut (.I0(GND_net), .I1(n14145[5]), .I2(n518_adj_4783), 
            .I3(n50113), .O(n13220[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_8 (.CI(n50113), .I0(n14145[5]), .I1(n518_adj_4783), 
            .CO(n50114));
    SB_CARRY add_6367_5 (.CI(n49883), .I0(n18485[2]), .I1(n320_adj_4777), 
            .CO(n49884));
    SB_LUT4 add_6121_7_lut (.I0(GND_net), .I1(n14145[4]), .I2(n445_adj_4784), 
            .I3(n50112), .O(n13220[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n49598), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n1[17]), .CO(n49599));
    SB_LUT4 add_6367_4_lut (.I0(GND_net), .I1(n18485[1]), .I2(n247_adj_4785), 
            .I3(n49882), .O(n18065[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_7 (.CI(n50112), .I0(n14145[4]), .I1(n445_adj_4784), 
            .CO(n50113));
    SB_CARRY add_6367_4 (.CI(n49882), .I0(n18485[1]), .I1(n247_adj_4785), 
            .CO(n49883));
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4721));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_19 (.CI(n49737), .I0(GND_net), .I1(n1_adj_4985[17]), 
            .CO(n49738));
    SB_LUT4 add_6367_3_lut (.I0(GND_net), .I1(n18485[0]), .I2(n174_adj_4786), 
            .I3(n49881), .O(n18065[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_6_lut (.I0(GND_net), .I1(n14145[3]), .I2(n372_adj_4787), 
            .I3(n50111), .O(n13220[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6367_3 (.CI(n49881), .I0(n18485[0]), .I1(n174_adj_4786), 
            .CO(n49882));
    SB_CARRY add_6121_6 (.CI(n50111), .I0(n14145[3]), .I1(n372_adj_4787), 
            .CO(n50112));
    SB_LUT4 add_6367_2_lut (.I0(GND_net), .I1(n32_adj_4788), .I2(n101_adj_4789), 
            .I3(GND_net), .O(n18065[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6367_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_5_lut (.I0(GND_net), .I1(n14145[2]), .I2(n299_adj_4790), 
            .I3(n50110), .O(n13220[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_5 (.CI(n50110), .I0(n14145[2]), .I1(n299_adj_4790), 
            .CO(n50111));
    SB_LUT4 add_6121_4_lut (.I0(GND_net), .I1(n14145[1]), .I2(n226_adj_4791), 
            .I3(n50109), .O(n13220[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n1[16]), .I3(n49597), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_4 (.CI(n50109), .I0(n14145[1]), .I1(n226_adj_4791), 
            .CO(n50110));
    SB_CARRY add_6367_2 (.CI(GND_net), .I0(n32_adj_4788), .I1(n101_adj_4789), 
            .CO(n49881));
    SB_LUT4 add_6121_3_lut (.I0(GND_net), .I1(n14145[0]), .I2(n153_adj_4792), 
            .I3(n50108), .O(n13220[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_3 (.CI(n50108), .I0(n14145[0]), .I1(n153_adj_4792), 
            .CO(n50109));
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[16]), 
            .I3(n49736), .O(n436[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6121_2_lut (.I0(GND_net), .I1(n11_adj_4794), .I2(n80_adj_4795), 
            .I3(GND_net), .O(n13220[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6121_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6121_2 (.CI(GND_net), .I0(n11_adj_4794), .I1(n80_adj_4795), 
            .CO(n50108));
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4720));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_18 (.CI(n49597), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n1[16]), .CO(n49598));
    SB_CARRY unary_minus_26_add_3_18 (.CI(n49736), .I0(GND_net), .I1(n1_adj_4985[16]), 
            .CO(n49737));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[15]), 
            .I3(n49735), .O(n436[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n1[15]), .I3(n49596), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_17 (.CI(n49735), .I0(GND_net), .I1(n1_adj_4985[15]), 
            .CO(n49736));
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[14]), 
            .I3(n49734), .O(n436[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_17 (.CI(n49596), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n1[15]), .CO(n49597));
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n1[14]), .I3(n49595), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_16 (.CI(n49734), .I0(GND_net), .I1(n1_adj_4985[14]), 
            .CO(n49735));
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[13]), 
            .I3(n49733), .O(n436[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_16 (.CI(n49595), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n1[14]), .CO(n49596));
    SB_LUT4 add_6163_21_lut (.I0(GND_net), .I1(n14985[18]), .I2(GND_net), 
            .I3(n50091), .O(n14145[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n1[13]), .I3(n49594), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_15 (.CI(n49594), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n1[13]), .CO(n49595));
    SB_LUT4 add_6521_8_lut (.I0(GND_net), .I1(n20129[5]), .I2(n560), .I3(n49871), 
            .O(n20032[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n1[12]), .I3(n49593), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_14 (.CI(n49593), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n1[12]), .CO(n49594));
    SB_LUT4 add_6163_20_lut (.I0(GND_net), .I1(n14985[17]), .I2(GND_net), 
            .I3(n50090), .O(n14145[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_15 (.CI(n49733), .I0(GND_net), .I1(n1_adj_4985[13]), 
            .CO(n49734));
    SB_LUT4 add_6521_7_lut (.I0(GND_net), .I1(n20129[4]), .I2(n487), .I3(n49870), 
            .O(n20032[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[12]), 
            .I3(n49732), .O(n436[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_20 (.CI(n50090), .I0(n14985[17]), .I1(GND_net), 
            .CO(n50091));
    SB_LUT4 add_6163_19_lut (.I0(GND_net), .I1(n14985[16]), .I2(GND_net), 
            .I3(n50089), .O(n14145[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_19 (.CI(n50089), .I0(n14985[16]), .I1(GND_net), 
            .CO(n50090));
    SB_CARRY add_6521_7 (.CI(n49870), .I0(n20129[4]), .I1(n487), .CO(n49871));
    SB_LUT4 add_6163_18_lut (.I0(GND_net), .I1(n14985[15]), .I2(GND_net), 
            .I3(n50088), .O(n14145[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n1[11]), .I3(n49592), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_13 (.CI(n49592), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n1[11]), .CO(n49593));
    SB_CARRY add_6163_18 (.CI(n50088), .I0(n14985[15]), .I1(GND_net), 
            .CO(n50089));
    SB_LUT4 add_6163_17_lut (.I0(GND_net), .I1(n14985[14]), .I2(GND_net), 
            .I3(n50087), .O(n14145[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_6_lut (.I0(GND_net), .I1(n20129[3]), .I2(n414), .I3(n49869), 
            .O(n20032[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_6 (.CI(n49869), .I0(n20129[3]), .I1(n414), .CO(n49870));
    SB_CARRY add_6163_17 (.CI(n50087), .I0(n14985[14]), .I1(GND_net), 
            .CO(n50088));
    SB_LUT4 add_6163_16_lut (.I0(GND_net), .I1(n14985[13]), .I2(n1105), 
            .I3(n50086), .O(n14145[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_5_lut (.I0(GND_net), .I1(n20129[2]), .I2(n341), .I3(n49868), 
            .O(n20032[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_16 (.CI(n50086), .I0(n14985[13]), .I1(n1105), .CO(n50087));
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n1[10]), .I3(n49591), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_12 (.CI(n49591), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n1[10]), .CO(n49592));
    SB_CARRY add_6521_5 (.CI(n49868), .I0(n20129[2]), .I1(n341), .CO(n49869));
    SB_LUT4 add_6163_15_lut (.I0(GND_net), .I1(n14985[12]), .I2(n1032), 
            .I3(n50085), .O(n14145[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_14 (.CI(n49732), .I0(GND_net), .I1(n1_adj_4985[12]), 
            .CO(n49733));
    SB_CARRY add_6163_15 (.CI(n50085), .I0(n14985[12]), .I1(n1032), .CO(n50086));
    SB_LUT4 add_6163_14_lut (.I0(GND_net), .I1(n14985[11]), .I2(n959), 
            .I3(n50084), .O(n14145[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_14 (.CI(n50084), .I0(n14985[11]), .I1(n959), .CO(n50085));
    SB_LUT4 add_6163_13_lut (.I0(GND_net), .I1(n14985[10]), .I2(n886), 
            .I3(n50083), .O(n14145[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_13 (.CI(n50083), .I0(n14985[10]), .I1(n886), .CO(n50084));
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n1[9]), .I3(n49590), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[11]), 
            .I3(n49731), .O(n436[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_12_lut (.I0(GND_net), .I1(n14985[9]), .I2(n813), 
            .I3(n50082), .O(n14145[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_12 (.CI(n50082), .I0(n14985[9]), .I1(n813), .CO(n50083));
    SB_CARRY add_9_11 (.CI(n49590), .I0(\PID_CONTROLLER.integral [9]), .I1(n1[9]), 
            .CO(n49591));
    SB_LUT4 add_6163_11_lut (.I0(GND_net), .I1(n14985[8]), .I2(n740), 
            .I3(n50081), .O(n14145[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_4_lut (.I0(GND_net), .I1(n20129[1]), .I2(n268), .I3(n49867), 
            .O(n20032[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_4 (.CI(n49867), .I0(n20129[1]), .I1(n268), .CO(n49868));
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4719));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n49731), .I0(GND_net), .I1(n1_adj_4985[11]), 
            .CO(n49732));
    SB_LUT4 add_6521_3_lut (.I0(GND_net), .I1(n20129[0]), .I2(n195), .I3(n49866), 
            .O(n20032[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[10]), 
            .I3(n49730), .O(n436[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_11 (.CI(n50081), .I0(n14985[8]), .I1(n740), .CO(n50082));
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n1[8]), .I3(n49589), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_10_lut (.I0(GND_net), .I1(n14985[7]), .I2(n667), 
            .I3(n50080), .O(n14145[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_3 (.CI(n49866), .I0(n20129[0]), .I1(n195), .CO(n49867));
    SB_CARRY add_9_10 (.CI(n49589), .I0(\PID_CONTROLLER.integral [8]), .I1(n1[8]), 
            .CO(n49590));
    SB_LUT4 add_6521_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20032[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n49866));
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4718));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_12 (.CI(n49730), .I0(GND_net), .I1(n1_adj_4985[10]), 
            .CO(n49731));
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n1[7]), .I3(n49588), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_14_lut (.I0(GND_net), .I1(n18849[11]), .I2(n980), 
            .I3(n49865), .O(n18485[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_10 (.CI(n50080), .I0(n14985[7]), .I1(n667), .CO(n50081));
    SB_LUT4 add_6163_9_lut (.I0(GND_net), .I1(n14985[6]), .I2(n594), .I3(n50079), 
            .O(n14145[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4717));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6163_9 (.CI(n50079), .I0(n14985[6]), .I1(n594), .CO(n50080));
    SB_LUT4 add_6394_13_lut (.I0(GND_net), .I1(n18849[10]), .I2(n907), 
            .I3(n49864), .O(n18485[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_13 (.CI(n49864), .I0(n18849[10]), .I1(n907), .CO(n49865));
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[9]), 
            .I3(n49729), .O(n436[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_9 (.CI(n49588), .I0(\PID_CONTROLLER.integral [7]), .I1(n1[7]), 
            .CO(n49589));
    SB_LUT4 add_6163_8_lut (.I0(GND_net), .I1(n14985[5]), .I2(n521), .I3(n50078), 
            .O(n14145[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_8 (.CI(n50078), .I0(n14985[5]), .I1(n521), .CO(n50079));
    SB_LUT4 add_6394_12_lut (.I0(GND_net), .I1(n18849[9]), .I2(n834), 
            .I3(n49863), .O(n18485[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_12 (.CI(n49863), .I0(n18849[9]), .I1(n834), .CO(n49864));
    SB_LUT4 add_6394_11_lut (.I0(GND_net), .I1(n18849[8]), .I2(n761), 
            .I3(n49862), .O(n18485[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_11 (.CI(n49862), .I0(n18849[8]), .I1(n761), .CO(n49863));
    SB_LUT4 add_6394_10_lut (.I0(GND_net), .I1(n18849[7]), .I2(n688), 
            .I3(n49861), .O(n18485[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_11 (.CI(n49729), .I0(GND_net), .I1(n1_adj_4985[9]), 
            .CO(n49730));
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4716));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6394_10 (.CI(n49861), .I0(n18849[7]), .I1(n688), .CO(n49862));
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[8]), 
            .I3(n49728), .O(n436[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n49728), .I0(GND_net), .I1(n1_adj_4985[8]), 
            .CO(n49729));
    SB_LUT4 add_6163_7_lut (.I0(GND_net), .I1(n14985[4]), .I2(n448), .I3(n50077), 
            .O(n14145[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_7 (.CI(n50077), .I0(n14985[4]), .I1(n448), .CO(n50078));
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[7]), 
            .I3(n49727), .O(n436[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_6_lut (.I0(GND_net), .I1(n14985[3]), .I2(n375), .I3(n50076), 
            .O(n14145[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_6 (.CI(n50076), .I0(n14985[3]), .I1(n375), .CO(n50077));
    SB_CARRY unary_minus_26_add_3_9 (.CI(n49727), .I0(GND_net), .I1(n1_adj_4985[7]), 
            .CO(n49728));
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[6]), 
            .I3(n49726), .O(n436[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_9_lut (.I0(GND_net), .I1(n18849[6]), .I2(n615_adj_4799), 
            .I3(n49860), .O(n18485[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_9 (.CI(n49860), .I0(n18849[6]), .I1(n615_adj_4799), 
            .CO(n49861));
    SB_CARRY unary_minus_26_add_3_8 (.CI(n49726), .I0(GND_net), .I1(n1_adj_4985[6]), 
            .CO(n49727));
    SB_LUT4 add_6394_8_lut (.I0(GND_net), .I1(n18849[5]), .I2(n542_adj_4800), 
            .I3(n49859), .O(n18485[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_5_lut (.I0(GND_net), .I1(n14985[2]), .I2(n302_adj_4801), 
            .I3(n50075), .O(n14145[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_8 (.CI(n49859), .I0(n18849[5]), .I1(n542_adj_4800), 
            .CO(n49860));
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n1[6]), .I3(n49587), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_5 (.CI(n50075), .I0(n14985[2]), .I1(n302_adj_4801), 
            .CO(n50076));
    SB_LUT4 add_6394_7_lut (.I0(GND_net), .I1(n18849[4]), .I2(n469_adj_4802), 
            .I3(n49858), .O(n18485[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_4_lut (.I0(GND_net), .I1(n14985[1]), .I2(n229_adj_4803), 
            .I3(n50074), .O(n14145[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_7 (.CI(n49858), .I0(n18849[4]), .I1(n469_adj_4802), 
            .CO(n49859));
    SB_CARRY add_6163_4 (.CI(n50074), .I0(n14985[1]), .I1(n229_adj_4803), 
            .CO(n50075));
    SB_CARRY add_9_8 (.CI(n49587), .I0(\PID_CONTROLLER.integral [6]), .I1(n1[6]), 
            .CO(n49588));
    SB_LUT4 add_6394_6_lut (.I0(GND_net), .I1(n18849[3]), .I2(n396_adj_4804), 
            .I3(n49857), .O(n18485[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_3_lut (.I0(GND_net), .I1(n14985[0]), .I2(n156_adj_4805), 
            .I3(n50073), .O(n14145[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_6 (.CI(n49857), .I0(n18849[3]), .I1(n396_adj_4804), 
            .CO(n49858));
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[5]), 
            .I3(n49725), .O(n436[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_5_lut (.I0(GND_net), .I1(n18849[2]), .I2(n323_adj_4807), 
            .I3(n49856), .O(n18485[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_5 (.CI(n49856), .I0(n18849[2]), .I1(n323_adj_4807), 
            .CO(n49857));
    SB_LUT4 add_6394_4_lut (.I0(GND_net), .I1(n18849[1]), .I2(n250_adj_4808), 
            .I3(n49855), .O(n18485[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n49725), .I0(GND_net), .I1(n1_adj_4985[5]), 
            .CO(n49726));
    SB_CARRY add_6163_3 (.CI(n50073), .I0(n14985[0]), .I1(n156_adj_4805), 
            .CO(n50074));
    SB_CARRY add_6394_4 (.CI(n49855), .I0(n18849[1]), .I1(n250_adj_4808), 
            .CO(n49856));
    SB_LUT4 add_6394_3_lut (.I0(GND_net), .I1(n18849[0]), .I2(n177_adj_4809), 
            .I3(n49854), .O(n18485[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[4]), 
            .I3(n49724), .O(n436[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6163_2_lut (.I0(GND_net), .I1(n14_adj_4811), .I2(n83_adj_4812), 
            .I3(GND_net), .O(n14145[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6163_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6163_2 (.CI(GND_net), .I0(n14_adj_4811), .I1(n83_adj_4812), 
            .CO(n50073));
    SB_CARRY add_6394_3 (.CI(n49854), .I0(n18849[0]), .I1(n177_adj_4809), 
            .CO(n49855));
    SB_CARRY unary_minus_26_add_3_6 (.CI(n49724), .I0(GND_net), .I1(n1_adj_4985[4]), 
            .CO(n49725));
    SB_LUT4 add_6394_2_lut (.I0(GND_net), .I1(n35_adj_4813), .I2(n104_adj_4814), 
            .I3(GND_net), .O(n18485[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_2 (.CI(GND_net), .I0(n35_adj_4813), .I1(n104_adj_4814), 
            .CO(n49854));
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n1[5]), .I3(n49586), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_7 (.CI(n49586), .I0(\PID_CONTROLLER.integral [5]), .I1(n1[5]), 
            .CO(n49587));
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[3]), 
            .I3(n49723), .O(n436[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_5 (.CI(n49723), .I0(GND_net), .I1(n1_adj_4985[3]), 
            .CO(n49724));
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[2]), 
            .I3(n49722), .O(n436[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_4 (.CI(n49722), .I0(GND_net), .I1(n1_adj_4985[2]), 
            .CO(n49723));
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n1[4]), .I3(n49585), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_6 (.CI(n49585), .I0(\PID_CONTROLLER.integral [4]), .I1(n1[4]), 
            .CO(n49586));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n1[3]), .I3(n49584), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_5 (.CI(n49584), .I0(\PID_CONTROLLER.integral [3]), .I1(n1[3]), 
            .CO(n49585));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[1]), 
            .I3(n49721), .O(n459)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n1[2]), .I3(n49583), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n49721), .I0(GND_net), .I1(n1_adj_4985[1]), 
            .CO(n49722));
    SB_LUT4 add_6419_13_lut (.I0(GND_net), .I1(n19161[10]), .I2(n910_adj_4820), 
            .I3(n49845), .O(n18849[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4985[0]), 
            .I3(VCC_net), .O(n460)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6419_12_lut (.I0(GND_net), .I1(n19161[9]), .I2(n837_adj_4823), 
            .I3(n49844), .O(n18849[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_12 (.CI(n49844), .I0(n19161[9]), .I1(n837_adj_4823), 
            .CO(n49845));
    SB_LUT4 add_6419_11_lut (.I0(GND_net), .I1(n19161[8]), .I2(n764_adj_4824), 
            .I3(n49843), .O(n18849[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_11 (.CI(n49843), .I0(n19161[8]), .I1(n764_adj_4824), 
            .CO(n49844));
    SB_LUT4 add_6419_10_lut (.I0(GND_net), .I1(n19161[7]), .I2(n691_adj_4825), 
            .I3(n49842), .O(n18849[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4985[0]), 
            .CO(n49721));
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n356[23]), .I1(GND_net), .I2(n1_adj_4986[23]), 
            .I3(n49720), .O(n47_adj_4498)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6419_10 (.CI(n49842), .I0(n19161[7]), .I1(n691_adj_4825), 
            .CO(n49843));
    SB_CARRY add_9_4 (.CI(n49583), .I0(\PID_CONTROLLER.integral [2]), .I1(n1[2]), 
            .CO(n49584));
    SB_LUT4 add_6473_11_lut (.I0(GND_net), .I1(n19744[8]), .I2(n770_adj_4827), 
            .I3(n50057), .O(n19545[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6473_10_lut (.I0(GND_net), .I1(n19744[7]), .I2(n697_adj_4828), 
            .I3(n50056), .O(n19545[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_10 (.CI(n50056), .I0(n19744[7]), .I1(n697_adj_4828), 
            .CO(n50057));
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[22]), 
            .I3(n49719), .O(n382[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n1[1]), .I3(n49582), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6419_9_lut (.I0(GND_net), .I1(n19161[6]), .I2(n618_adj_4830), 
            .I3(n49841), .O(n18849[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n49719), .I0(GND_net), .I1(n1_adj_4986[22]), 
            .CO(n49720));
    SB_LUT4 add_6473_9_lut (.I0(GND_net), .I1(n19744[6]), .I2(n624_adj_4831), 
            .I3(n50055), .O(n19545[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[21]), 
            .I3(n49718), .O(n382[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_9 (.CI(n49841), .I0(n19161[6]), .I1(n618_adj_4830), 
            .CO(n49842));
    SB_LUT4 add_6419_8_lut (.I0(GND_net), .I1(n19161[5]), .I2(n545_adj_4833), 
            .I3(n49840), .O(n18849[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_9 (.CI(n50055), .I0(n19744[6]), .I1(n624_adj_4831), 
            .CO(n50056));
    SB_LUT4 add_6473_8_lut (.I0(GND_net), .I1(n19744[5]), .I2(n551_adj_4834), 
            .I3(n50054), .O(n19545[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_8 (.CI(n50054), .I0(n19744[5]), .I1(n551_adj_4834), 
            .CO(n50055));
    SB_LUT4 add_6473_7_lut (.I0(GND_net), .I1(n19744[4]), .I2(n478_adj_4835), 
            .I3(n50053), .O(n19545[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_7 (.CI(n50053), .I0(n19744[4]), .I1(n478_adj_4835), 
            .CO(n50054));
    SB_CARRY add_6419_8 (.CI(n49840), .I0(n19161[5]), .I1(n545_adj_4833), 
            .CO(n49841));
    SB_LUT4 add_6473_6_lut (.I0(GND_net), .I1(n19744[3]), .I2(n405_adj_4836), 
            .I3(n50052), .O(n19545[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_6 (.CI(n50052), .I0(n19744[3]), .I1(n405_adj_4836), 
            .CO(n50053));
    SB_LUT4 add_6473_5_lut (.I0(GND_net), .I1(n19744[2]), .I2(n332_adj_4837), 
            .I3(n50051), .O(n19545[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_5 (.CI(n50051), .I0(n19744[2]), .I1(n332_adj_4837), 
            .CO(n50052));
    SB_LUT4 add_6473_4_lut (.I0(GND_net), .I1(n19744[1]), .I2(n259_adj_4838), 
            .I3(n50050), .O(n19545[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6419_7_lut (.I0(GND_net), .I1(n19161[4]), .I2(n472_adj_4839), 
            .I3(n49839), .O(n18849[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_4 (.CI(n50050), .I0(n19744[1]), .I1(n259_adj_4838), 
            .CO(n50051));
    SB_LUT4 add_6473_3_lut (.I0(GND_net), .I1(n19744[0]), .I2(n186_adj_4840), 
            .I3(n50049), .O(n19545[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_7 (.CI(n49839), .I0(n19161[4]), .I1(n472_adj_4839), 
            .CO(n49840));
    SB_LUT4 add_6419_6_lut (.I0(GND_net), .I1(n19161[3]), .I2(n399_adj_4841), 
            .I3(n49838), .O(n18849[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_3 (.CI(n49582), .I0(\PID_CONTROLLER.integral [1]), .I1(n1[1]), 
            .CO(n49583));
    SB_CARRY add_6473_3 (.CI(n50049), .I0(n19744[0]), .I1(n186_adj_4840), 
            .CO(n50050));
    SB_LUT4 add_6473_2_lut (.I0(GND_net), .I1(n44_adj_4842), .I2(n113_adj_4843), 
            .I3(GND_net), .O(n19545[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_6 (.CI(n49838), .I0(n19161[3]), .I1(n399_adj_4841), 
            .CO(n49839));
    SB_LUT4 add_6419_5_lut (.I0(GND_net), .I1(n19161[2]), .I2(n326_adj_4844), 
            .I3(n49837), .O(n18849[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n49718), .I0(GND_net), .I1(n1_adj_4986[21]), 
            .CO(n49719));
    SB_CARRY add_6473_2 (.CI(GND_net), .I0(n44_adj_4842), .I1(n113_adj_4843), 
            .CO(n50049));
    SB_LUT4 add_6202_20_lut (.I0(GND_net), .I1(n15745[17]), .I2(GND_net), 
            .I3(n50048), .O(n14985[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[20]), 
            .I3(n49717), .O(n382[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_5 (.CI(n49837), .I0(n19161[2]), .I1(n326_adj_4844), 
            .CO(n49838));
    SB_CARRY unary_minus_20_add_3_22 (.CI(n49717), .I0(GND_net), .I1(n1_adj_4986[20]), 
            .CO(n49718));
    SB_LUT4 add_6202_19_lut (.I0(GND_net), .I1(n15745[16]), .I2(GND_net), 
            .I3(n50047), .O(n14985[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6419_4_lut (.I0(GND_net), .I1(n19161[1]), .I2(n253_adj_4846), 
            .I3(n49836), .O(n18849[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_19 (.CI(n50047), .I0(n15745[16]), .I1(GND_net), 
            .CO(n50048));
    SB_LUT4 add_6202_18_lut (.I0(GND_net), .I1(n15745[15]), .I2(GND_net), 
            .I3(n50046), .O(n14985[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_18 (.CI(n50046), .I0(n15745[15]), .I1(GND_net), 
            .CO(n50047));
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n1[0]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n1[0]), 
            .CO(n49582));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[19]), 
            .I3(n49716), .O(n382[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6202_17_lut (.I0(GND_net), .I1(n15745[14]), .I2(GND_net), 
            .I3(n50045), .O(n14985[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n49716), .I0(GND_net), .I1(n1_adj_4986[19]), 
            .CO(n49717));
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n49581), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_4 (.CI(n49836), .I0(n19161[1]), .I1(n253_adj_4846), 
            .CO(n49837));
    SB_CARRY add_6202_17 (.CI(n50045), .I0(n15745[14]), .I1(GND_net), 
            .CO(n50046));
    SB_LUT4 add_6202_16_lut (.I0(GND_net), .I1(n15745[13]), .I2(n1108_adj_4848), 
            .I3(n50044), .O(n14985[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_16 (.CI(n50044), .I0(n15745[13]), .I1(n1108_adj_4848), 
            .CO(n50045));
    SB_LUT4 add_6202_15_lut (.I0(GND_net), .I1(n15745[12]), .I2(n1035_adj_4849), 
            .I3(n50043), .O(n14985[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[18]), 
            .I3(n49715), .O(n382[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_15 (.CI(n50043), .I0(n15745[12]), .I1(n1035_adj_4849), 
            .CO(n50044));
    SB_LUT4 add_6202_14_lut (.I0(GND_net), .I1(n15745[11]), .I2(n962_adj_4851), 
            .I3(n50042), .O(n14985[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6419_3_lut (.I0(GND_net), .I1(n19161[0]), .I2(n180_adj_4852), 
            .I3(n49835), .O(n18849[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_14 (.CI(n50042), .I0(n15745[11]), .I1(n962_adj_4851), 
            .CO(n50043));
    SB_LUT4 add_6202_13_lut (.I0(GND_net), .I1(n15745[10]), .I2(n889_adj_4853), 
            .I3(n50041), .O(n14985[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_13 (.CI(n50041), .I0(n15745[10]), .I1(n889_adj_4853), 
            .CO(n50042));
    SB_LUT4 add_6202_12_lut (.I0(GND_net), .I1(n15745[9]), .I2(n816_adj_4854), 
            .I3(n50040), .O(n14985[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_12 (.CI(n50040), .I0(n15745[9]), .I1(n816_adj_4854), 
            .CO(n50041));
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n49580), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_3 (.CI(n49835), .I0(n19161[0]), .I1(n180_adj_4852), 
            .CO(n49836));
    SB_LUT4 add_6419_2_lut (.I0(GND_net), .I1(n38_adj_4855), .I2(n107_adj_4856), 
            .I3(GND_net), .O(n18849[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_2 (.CI(GND_net), .I0(n38_adj_4855), .I1(n107_adj_4856), 
            .CO(n49835));
    SB_LUT4 add_6202_11_lut (.I0(GND_net), .I1(n15745[8]), .I2(n743_adj_4857), 
            .I3(n50039), .O(n14985[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_11 (.CI(n50039), .I0(n15745[8]), .I1(n743_adj_4857), 
            .CO(n50040));
    SB_LUT4 add_6202_10_lut (.I0(GND_net), .I1(n15745[7]), .I2(n670_adj_4858), 
            .I3(n50038), .O(n14985[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_10 (.CI(n50038), .I0(n15745[7]), .I1(n670_adj_4858), 
            .CO(n50039));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n49715), .I0(GND_net), .I1(n1_adj_4986[18]), 
            .CO(n49716));
    SB_LUT4 add_6202_9_lut (.I0(GND_net), .I1(n15745[6]), .I2(n597_adj_4859), 
            .I3(n50037), .O(n14985[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[17]), 
            .I3(n49714), .O(n382[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n49714), .I0(GND_net), .I1(n1_adj_4986[17]), 
            .CO(n49715));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[16]), 
            .I3(n49713), .O(n382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_9 (.CI(n50037), .I0(n15745[6]), .I1(n597_adj_4859), 
            .CO(n50038));
    SB_LUT4 add_6202_8_lut (.I0(GND_net), .I1(n15745[5]), .I2(n524_adj_4862), 
            .I3(n50036), .O(n14985[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_24 (.CI(n49580), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n49581));
    SB_CARRY add_6202_8 (.CI(n50036), .I0(n15745[5]), .I1(n524_adj_4862), 
            .CO(n50037));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n49713), .I0(GND_net), .I1(n1_adj_4986[16]), 
            .CO(n49714));
    SB_LUT4 add_6202_7_lut (.I0(GND_net), .I1(n15745[4]), .I2(n451_adj_4863), 
            .I3(n50035), .O(n14985[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_7 (.CI(n50035), .I0(n15745[4]), .I1(n451_adj_4863), 
            .CO(n50036));
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n49579), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6202_6_lut (.I0(GND_net), .I1(n15745[3]), .I2(n378_adj_4864), 
            .I3(n50034), .O(n14985[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_6 (.CI(n50034), .I0(n15745[3]), .I1(n378_adj_4864), 
            .CO(n50035));
    SB_LUT4 add_6202_5_lut (.I0(GND_net), .I1(n15745[2]), .I2(n305_adj_4865), 
            .I3(n50033), .O(n14985[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[15]), 
            .I3(n49712), .O(n382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_5 (.CI(n50033), .I0(n15745[2]), .I1(n305_adj_4865), 
            .CO(n50034));
    SB_LUT4 add_6202_4_lut (.I0(GND_net), .I1(n15745[1]), .I2(n232_adj_4867), 
            .I3(n50032), .O(n14985[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n49712), .I0(GND_net), .I1(n1_adj_4986[15]), 
            .CO(n49713));
    SB_CARRY add_6202_4 (.CI(n50032), .I0(n15745[1]), .I1(n232_adj_4867), 
            .CO(n50033));
    SB_CARRY sub_8_add_2_23 (.CI(n49579), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n49580));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[14]), 
            .I3(n49711), .O(n382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6202_3_lut (.I0(GND_net), .I1(n15745[0]), .I2(n159_adj_4869), 
            .I3(n50031), .O(n14985[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n219));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6202_3 (.CI(n50031), .I0(n15745[0]), .I1(n159_adj_4869), 
            .CO(n50032));
    SB_LUT4 add_6202_2_lut (.I0(GND_net), .I1(n17_adj_4870), .I2(n86_adj_4871), 
            .I3(GND_net), .O(n14985[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6202_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6202_2 (.CI(GND_net), .I0(n17_adj_4870), .I1(n86_adj_4871), 
            .CO(n50031));
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n49578), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4715));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_22 (.CI(n49578), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n49579));
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n49577), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n49711), .I0(GND_net), .I1(n1_adj_4986[14]), 
            .CO(n49712));
    SB_LUT4 add_6533_7_lut (.I0(GND_net), .I1(n60309), .I2(n490), .I3(n49827), 
            .O(n20129[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6533_6_lut (.I0(GND_net), .I1(n20200[3]), .I2(n417), .I3(n49826), 
            .O(n20129[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6533_6 (.CI(n49826), .I0(n20200[3]), .I1(n417), .CO(n49827));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[13]), 
            .I3(n49710), .O(n382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_21 (.CI(n49577), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n49578));
    SB_CARRY unary_minus_20_add_3_15 (.CI(n49710), .I0(GND_net), .I1(n1_adj_4986[13]), 
            .CO(n49711));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[12]), 
            .I3(n49709), .O(n382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n49576), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6533_5_lut (.I0(GND_net), .I1(n20203), .I2(n344), .I3(n49825), 
            .O(n20129[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_20 (.CI(n49576), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n49577));
    SB_CARRY add_6533_5 (.CI(n49825), .I0(n20203), .I1(n344), .CO(n49826));
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n49575), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n49709), .I0(GND_net), .I1(n1_adj_4986[12]), 
            .CO(n49710));
    SB_LUT4 add_6533_4_lut (.I0(GND_net), .I1(n20204), .I2(n271), .I3(n49824), 
            .O(n20129[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6533_4 (.CI(n49824), .I0(n20204), .I1(n271), .CO(n49825));
    SB_LUT4 add_6533_3_lut (.I0(GND_net), .I1(n20205), .I2(n198), .I3(n49823), 
            .O(n20129[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[11]), 
            .I3(n49708), .O(n382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6533_3 (.CI(n49823), .I0(n20205), .I1(n198), .CO(n49824));
    SB_CARRY unary_minus_20_add_3_13 (.CI(n49708), .I0(GND_net), .I1(n1_adj_4986[11]), 
            .CO(n49709));
    SB_LUT4 add_6533_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20129[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6533_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n49823));
    SB_CARRY sub_8_add_2_19 (.CI(n49575), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n49576));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[10]), 
            .I3(n49707), .O(n382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n49707), .I0(GND_net), .I1(n1_adj_4986[10]), 
            .CO(n49708));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[9]), 
            .I3(n49706), .O(n382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n49706), .I0(GND_net), .I1(n1_adj_4986[9]), 
            .CO(n49707));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[8]), 
            .I3(n49705), .O(n382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(n20), 
            .I3(n49574), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4713));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_18 (.CI(n49574), .I0(setpoint[16]), .I1(n20), 
            .CO(n49575));
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n49573), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_17 (.CI(n49573), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n49574));
    SB_CARRY unary_minus_20_add_3_10 (.CI(n49705), .I0(GND_net), .I1(n1_adj_4986[8]), 
            .CO(n49706));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[7]), 
            .I3(n49704), .O(n382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n49704), .I0(GND_net), .I1(n1_adj_4986[7]), 
            .CO(n49705));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[6]), 
            .I3(n49703), .O(n382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n49703), .I0(GND_net), .I1(n1_adj_4986[6]), 
            .CO(n49704));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[5]), 
            .I3(n49702), .O(n382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n11650[0]), .I2(n12229[0]), 
            .I3(n49627), .O(n356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n49702), .I0(GND_net), .I1(n1_adj_4986[5]), 
            .CO(n49703));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[4]), 
            .I3(n49701), .O(n382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n49572), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n49701), .I0(GND_net), .I1(n1_adj_4986[4]), 
            .CO(n49702));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[3]), 
            .I3(n49700), .O(n382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n49700), .I0(GND_net), .I1(n1_adj_4986[3]), 
            .CO(n49701));
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n306[22]), 
            .I3(n49626), .O(n356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_16 (.CI(n49572), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n49573));
    SB_LUT4 add_6239_19_lut (.I0(GND_net), .I1(n16429[16]), .I2(GND_net), 
            .I3(n50016), .O(n15745[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6239_18_lut (.I0(GND_net), .I1(n16429[15]), .I2(GND_net), 
            .I3(n50015), .O(n15745[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[2]), 
            .I3(n49699), .O(n382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_24 (.CI(n49626), .I0(n257[22]), .I1(n306[22]), .CO(n49627));
    SB_CARRY add_6239_18 (.CI(n50015), .I0(n16429[15]), .I1(GND_net), 
            .CO(n50016));
    SB_CARRY unary_minus_20_add_3_4 (.CI(n49699), .I0(GND_net), .I1(n1_adj_4986[2]), 
            .CO(n49700));
    SB_LUT4 add_6239_17_lut (.I0(GND_net), .I1(n16429[14]), .I2(GND_net), 
            .I3(n50014), .O(n15745[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4986[1]), 
            .I3(n49698), .O(n405)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_17 (.CI(n50014), .I0(n16429[14]), .I1(GND_net), 
            .CO(n50015));
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n306[21]), 
            .I3(n49625), .O(n356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n49571), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_15 (.CI(n49571), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n49572));
    SB_CARRY unary_minus_20_add_3_3 (.CI(n49698), .I0(GND_net), .I1(n1_adj_4986[1]), 
            .CO(n49699));
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n49570), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_23 (.CI(n49625), .I0(n257[21]), .I1(n306[21]), .CO(n49626));
    SB_LUT4 add_6239_16_lut (.I0(GND_net), .I1(n16429[13]), .I2(n1111_adj_4896), 
            .I3(n50013), .O(n15745[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_16 (.CI(n50013), .I0(n16429[13]), .I1(n1111_adj_4896), 
            .CO(n50014));
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4712));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6239_15_lut (.I0(GND_net), .I1(n16429[12]), .I2(n1038_adj_4897), 
            .I3(n50012), .O(n15745[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_14 (.CI(n49570), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n49571));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n37293), .I1(GND_net), .I2(n1_adj_4986[0]), 
            .I3(VCC_net), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n306[20]), 
            .I3(n49624), .O(n356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4711));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n49569), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_13 (.CI(n49569), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n49570));
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4900));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4710));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4709));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4708));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4901));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4902));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4903));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4707));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4904));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4905));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4906));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_966 (.I0(n20225[2]), .I1(n6_adj_4907), .I2(\Kp[4] ), 
            .I3(n1[18]), .O(n20165[3]));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_966.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_23_i7_2_lut (.I0(PWMLimit[3]), .I1(n356[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4908));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4909));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4795));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35508_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n20289[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35508_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_18_22 (.CI(n49624), .I0(n257[20]), .I1(n306[20]), .CO(n49625));
    SB_LUT4 mult_16_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4794));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6239_15 (.CI(n50012), .I0(n16429[12]), .I1(n1038_adj_4897), 
            .CO(n50013));
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4910));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[16]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_23_i5_2_lut (.I0(PWMLimit[2]), .I1(n356[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4911));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i5_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4986[0]), 
            .CO(n49698));
    SB_LUT4 add_6239_14_lut (.I0(GND_net), .I1(n16429[11]), .I2(n965_adj_4912), 
            .I3(n50011), .O(n15745[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50877_4_lut (.I0(n11_adj_4910), .I1(n9_adj_4909), .I2(n7_adj_4908), 
            .I3(n5_adj_4911), .O(n66605));
    defparam i50877_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6239_14 (.CI(n50011), .I0(n16429[11]), .I1(n965_adj_4912), 
            .CO(n50012));
    SB_LUT4 i50873_4_lut (.I0(n17_adj_4906), .I1(n15_adj_4905), .I2(n13_adj_4904), 
            .I3(n66605), .O(n66601));
    defparam i50873_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4792));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6239_13_lut (.I0(GND_net), .I1(n16429[10]), .I2(n892_adj_4913), 
            .I3(n50010), .O(n15745[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_4904), 
            .I3(GND_net), .O(n10_adj_4914));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_967 (.I0(\Kp[4] ), .I1(\Kp[5] ), .I2(n1[19]), 
            .I3(n1[18]), .O(n62242));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_967.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4791));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\Kp[3] ), .I1(n62242), .I2(n1[20]), .I3(GND_net), 
            .O(n62244));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4790));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i142_2_lut (.I0(\Kp[2] ), .I1(n1[21]), .I2(GND_net), 
            .I3(GND_net), .O(n210_adj_4915));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_968 (.I0(\Kp[1] ), .I1(n210_adj_4915), .I2(n1[22]), 
            .I3(n62244), .O(n62248));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_968.LUT_INIT = 16'h936c;
    SB_LUT4 i35510_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n49454));   // verilog/motorControl.v(50[18:24])
    defparam i35510_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[23]), 
            .I3(n49697), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4789));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4788));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4787));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4786));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_969 (.I0(n49454), .I1(\Kp[0] ), .I2(n62248), 
            .I3(n1[23]), .O(n62252));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_969.LUT_INIT = 16'h695a;
    SB_LUT4 i35430_4_lut (.I0(n20225[2]), .I1(\Kp[4] ), .I2(n6_adj_4907), 
            .I3(n1[18]), .O(n8_adj_4917));   // verilog/motorControl.v(50[18:24])
    defparam i35430_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_970 (.I0(n6_c), .I1(n8_adj_4917), .I2(n4_adj_4918), 
            .I3(n62252), .O(n59281));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[22]), 
            .I3(n49696), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n10_adj_4914), .I1(n356[7]), .I2(n15_adj_4905), 
            .I3(GND_net), .O(n12_adj_4920));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6239_13 (.CI(n50010), .I0(n16429[10]), .I1(n892_adj_4913), 
            .CO(n50011));
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_4906), 
            .I3(GND_net), .O(n8_adj_4921));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[11] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6239_12_lut (.I0(GND_net), .I1(n16429[9]), .I2(n819_adj_4923), 
            .I3(n50009), .O(n15745[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_12 (.CI(n50009), .I0(n16429[9]), .I1(n819_adj_4923), 
            .CO(n50010));
    SB_LUT4 add_6239_11_lut (.I0(GND_net), .I1(n16429[8]), .I2(n746_adj_4924), 
            .I3(n50008), .O(n15745[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_11 (.CI(n50008), .I0(n16429[8]), .I1(n746_adj_4924), 
            .CO(n50009));
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4706));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6239_10_lut (.I0(GND_net), .I1(n16429[7]), .I2(n673_adj_4925), 
            .I3(n50007), .O(n15745[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i6_3_lut (.I0(n356[2]), .I1(n356[3]), .I2(n7_adj_4908), 
            .I3(GND_net), .O(n6_adj_4926));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n8_adj_4921), .I1(n356[9]), .I2(n19_adj_4903), 
            .I3(GND_net), .O(n16_adj_4927));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52625_4_lut (.I0(n16_adj_4927), .I1(n6_adj_4926), .I2(n19_adj_4903), 
            .I3(n66599), .O(n68353));   // verilog/motorControl.v(52[14:29])
    defparam i52625_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52626_3_lut (.I0(n68353), .I1(n356[10]), .I2(n21_adj_4902), 
            .I3(GND_net), .O(n68354));   // verilog/motorControl.v(52[14:29])
    defparam i52626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52520_3_lut (.I0(n68354), .I1(n356[11]), .I2(n23_adj_4901), 
            .I3(GND_net), .O(n68248));   // verilog/motorControl.v(52[14:29])
    defparam i52520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52373_4_lut (.I0(n23_adj_4901), .I1(n21_adj_4902), .I2(n19_adj_4903), 
            .I3(n66601), .O(n68101));
    defparam i52373_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52423_4_lut (.I0(n12_adj_4920), .I1(n4_adj_7), .I2(n15_adj_4905), 
            .I3(n66603), .O(n68151));   // verilog/motorControl.v(52[14:29])
    defparam i52423_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6239_10 (.CI(n50007), .I0(n16429[7]), .I1(n673_adj_4925), 
            .CO(n50008));
    SB_LUT4 i51154_3_lut (.I0(n68248), .I1(n356[12]), .I2(n25_adj_4900), 
            .I3(GND_net), .O(n66882));   // verilog/motorControl.v(52[14:29])
    defparam i51154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52635_4_lut (.I0(n66882), .I1(n68151), .I2(n25_adj_4900), 
            .I3(n68101), .O(n68363));   // verilog/motorControl.v(52[14:29])
    defparam i52635_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n306[19]), 
            .I3(n49623), .O(n356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6239_9_lut (.I0(GND_net), .I1(n16429[6]), .I2(n600_adj_4929), 
            .I3(n50006), .O(n15745[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6239_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_24 (.CI(n49696), .I0(GND_net), .I1(n1_adj_4984[22]), 
            .CO(n49697));
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4984[21]), 
            .I3(n49695), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n49568), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6239_9 (.CI(n50006), .I0(n16429[6]), .I1(n600_adj_4929), 
            .CO(n50007));
    SB_LUT4 i52636_3_lut (.I0(n68363), .I1(n356[13]), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n68364));   // verilog/motorControl.v(52[14:29])
    defparam i52636_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52486_3_lut (.I0(n68364), .I1(n356[14]), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(52[14:29])
    defparam i52486_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6442_12_lut (.I0(GND_net), .I1(n19425[9]), .I2(n840_adj_4931), 
            .I3(n49811), .O(n19161[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4705));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4704));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4785));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4784));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4783));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4703));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[17]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4781));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4702));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4701));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4700));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4780));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[10] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4699));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4779));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[18]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4777));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4776));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4775));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4774));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4773));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4698));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4772));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4697));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4696));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4694));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4693));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4692));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4691));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4690));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4689));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4688));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4687));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4686));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4685));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4684));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50871_2_lut_4_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(PWMLimit[4]), 
            .I3(n356[4]), .O(n66599));
    defparam i50871_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4683));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50875_2_lut_4_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(PWMLimit[5]), 
            .I3(n356[5]), .O(n66603));
    defparam i50875_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i35342_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n20225[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35342_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(GND_net), .O(n6_adj_4932));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i50814_3_lut_4_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(n356[2]), .O(n66542));   // verilog/motorControl.v(54[23:39])
    defparam i50814_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[9] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4682));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4681));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4680));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4679));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4678));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4677));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4676));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4675));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4674));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4673));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4672));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4671));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4669));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[17]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[8] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4668));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4667));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4931));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4929));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4925));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4924));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4923));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[22]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[23]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4913));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4912));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4665));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23266_1_lut (.I0(n380), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37293));   // verilog/motorControl.v(50[18:38])
    defparam i23266_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4664));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4663));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[0]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4897));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4896));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[1]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[2]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[3]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[19]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[20]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[4]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[5]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[6]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[7]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4769));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4768));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4767));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[21]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4765));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4764));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4763));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4762));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4760));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[8]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[22]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[9]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4759));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4758));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[10]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4662));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[11]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4757));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4661));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4660));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4659));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[23]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50294_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n66022));   // verilog/motorControl.v(47[21:44])
    defparam i50294_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4657));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4756));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4656));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4655));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4653));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4652));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_adj_4599));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4651));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4650));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4649));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4648));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4647));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4646));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4645));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[12]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4644));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4643));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[13]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4641));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4640));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[7] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4639));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_971 (.I0(n20249[2]), .I1(n6), .I2(n36852), .I3(\Ki[4] ), 
            .O(n20200[3]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_971.LUT_INIT = 16'h9666;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4638));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4637));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4636));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4635));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4634));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4633));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4632));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4631));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50393_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n66121));   // verilog/motorControl.v(45[12:34])
    defparam i50393_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_4542));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i35327_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n20297[0]));   // verilog/motorControl.v(50[27:38])
    defparam i35327_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4629));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4628));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4627));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4626));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_972 (.I0(n20280[1]), .I1(n4_adj_8), .I2(n36823), 
            .I3(\Ki[3] ), .O(n20249[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h9666;
    SB_LUT4 i1_4_lut_adj_973 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[23] ), .O(n62200));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_973.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_974 (.I0(n36852), .I1(\Ki[2] ), .I2(\Ki[5] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n62202));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_974.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4625));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4624));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4623));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4622));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35552_4_lut (.I0(n20249[2]), .I1(n36852), .I2(n6), .I3(\Ki[4] ), 
            .O(n8_adj_4936));   // verilog/motorControl.v(50[27:38])
    defparam i35552_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4621));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4620));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35498_4_lut (.I0(n20280[1]), .I1(n36823), .I2(n4_adj_8), 
            .I3(\Ki[3] ), .O(n6_adj_4937));   // verilog/motorControl.v(50[27:38])
    defparam i35498_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4619));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4618));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4617));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4616));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_975 (.I0(n36823), .I1(\Ki[3] ), .I2(\Ki[4] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[20] ), .O(n62208));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_975.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[18]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4615));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4614));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4613));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4612));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4611));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35329_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n49260));   // verilog/motorControl.v(50[27:38])
    defparam i35329_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4610));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4609));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4608));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_976 (.I0(n6_adj_4937), .I1(n8_adj_4936), .I2(n62202), 
            .I3(n62200), .O(n60055));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[6] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4607));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4606));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4605));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(counter[17]), .I1(counter[22]), .I2(counter[21]), 
            .I3(counter[18]), .O(n60322));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_977 (.I0(n4_adj_4938), .I1(n60055), .I2(n49260), 
            .I3(n62208), .O(n60309));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4604));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4603));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4602));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_2_lut (.I0(counter[20]), .I1(counter[27]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4939));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4601));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11_4_lut (.I0(counter[19]), .I1(counter[26]), .I2(n60322), 
            .I3(counter[15]), .O(n26_adj_4940));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12_adj_4941));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4600));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(counter[5]), .I1(n12_adj_4941), .I2(counter[2]), 
            .I3(counter[0]), .O(n59546));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4598));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_4942));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i50127_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n65855));
    defparam i50127_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i3_4_lut_adj_978 (.I0(counter[12]), .I1(n59546), .I2(counter[8]), 
            .I3(counter[7]), .O(n9_adj_4943));
    defparam i3_4_lut_adj_978.LUT_INIT = 16'ha8a0;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut (.I0(counter[24]), .I1(counter[16]), .I2(counter[29]), 
            .I3(counter[14]), .O(n24_adj_4944));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(counter[28]), .I1(n26_adj_4940), .I2(n20_adj_4939), 
            .I3(counter[30]), .O(n28_adj_4945));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut (.I0(counter[25]), .I1(counter[23]), .I2(n9_adj_4943), 
            .I3(n10_adj_4942), .O(n23_adj_4946));
    defparam i8_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[16] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4595));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4594));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4593));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28977_4_lut (.I0(n23_adj_4946), .I1(counter[31]), .I2(n28_adj_4945), 
            .I3(n24_adj_4944), .O(counter_31__N_3714));   // verilog/motorControl.v(26[8:41])
    defparam i28977_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[19]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50173_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n65901));
    defparam i50173_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4871));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4870));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4592));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4869));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[14]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50296_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n66024));
    defparam i50296_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[20]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4591));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4590));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4589));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4867));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[15]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50329_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n66057));
    defparam i50329_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4587));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4865));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4586));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4585));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4584));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4583));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4582));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4864));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4578));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n306[0]));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[5] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4576));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4863));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4862));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[16]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[17]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4575));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4859));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4574));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4858));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4857));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4856));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4855));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[4] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4854));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4853));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4571));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4852));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4570));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4569));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4851));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4568));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4540));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4539));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4538));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[18]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4537));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4536));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4535));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4849));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4848));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[19]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4846));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4534));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4533));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[20]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4532));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4844));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4843));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4530));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4528));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4527));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_c));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4842));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4841));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[3] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4524));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4840));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4839));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4838));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4837));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4836));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4523));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4522));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4835));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4834));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4833));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[21]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4831));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4830));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[22]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[2] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4518));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4828));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4515));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4514));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4827));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4512));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4986[23]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4825));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4824));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4823));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[0]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4820));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[1]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[2]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[3]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[1] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4508));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29479_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43450));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29479_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4814));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4506));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4505));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4813));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4812));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4811));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[4]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4809));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4808));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4807));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[5]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4805));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4804));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4803));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4802));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4801));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4800));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4799));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4755));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4754));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4753));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50968_2_lut_4_lut (.I0(deadband[17]), .I1(n356[17]), .I2(deadband[8]), 
            .I3(n356[8]), .O(n66696));
    defparam i50968_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i35477_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(\Ki[1] ), .I3(n36823), .O(n20253));   // verilog/motorControl.v(50[27:38])
    defparam i35477_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i35479_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(\Ki[1] ), .I3(n36823), .O(n49420));   // verilog/motorControl.v(50[27:38])
    defparam i35479_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i35460_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(n49388), .I3(n20297[0]), .O(n4_adj_4938));   // verilog/motorControl.v(50[27:38])
    defparam i35460_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_979 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(n49388), .I3(n20297[0]), .O(n20280[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_979.LUT_INIT = 16'h8778;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35449_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), .I3(\Ki[1] ), 
            .O(n49388));   // verilog/motorControl.v(50[27:38])
    defparam i35449_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4984[21]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35447_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), .I3(\Ki[1] ), 
            .O(n20283));   // verilog/motorControl.v(50[27:38])
    defparam i35447_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i50068_2_lut_4_lut (.I0(deadband[9]), .I1(n356[9]), .I2(deadband[5]), 
            .I3(n356[5]), .O(n65796));
    defparam i50068_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n356[20]), .I1(n436[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4949));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n356[19]), .I1(n436[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4950));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n356[22]), .I1(n436[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4951));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n356[21]), .I1(n436[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4952));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n356[18]), .I1(n436[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4953));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n356[14]), .I1(n436[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4954));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n365), .I1(n436[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4955));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n356[11]), .I1(n436[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4956));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_3_lut (.I0(n380), .I1(PWMLimit[0]), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(50[18:38])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n356[12]), .I1(n436[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4958));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n356[17]), .I1(n436[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4959));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n356[16]), .I1(n436[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4960));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n356[4]), .I1(n436[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4961));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n356[8]), .I1(n436[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4962));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n356[9]), .I1(n436[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4963));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n356[10]), .I1(n436[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4964));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n356[5]), .I1(n436[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4965));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n356[6]), .I1(n436[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4966));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n356[7]), .I1(n436[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4967));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n356[13]), .I1(n436[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4968));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50798_4_lut (.I0(n21_adj_4964), .I1(n19_adj_4963), .I2(n17_adj_4962), 
            .I3(n9_adj_4961), .O(n66526));
    defparam i50798_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50786_4_lut (.I0(n27_adj_4968), .I1(n15_adj_4967), .I2(n13_adj_4966), 
            .I3(n11_adj_4965), .O(n66514));
    defparam i50786_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n436[7]), .I1(n436[16]), .I2(n33_adj_4960), 
            .I3(GND_net), .O(n12_adj_4969));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n436[5]), .I1(n436[6]), .I2(n13_adj_4966), 
            .I3(GND_net), .O(n10_adj_4970));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12_adj_4969), .I1(n436[17]), .I2(n35_adj_4959), 
            .I3(GND_net), .O(n30_adj_4971));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51692_4_lut (.I0(n13_adj_4966), .I1(n11_adj_4965), .I2(n9_adj_4961), 
            .I3(n66542), .O(n67420));
    defparam i51692_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51682_4_lut (.I0(n19_adj_4963), .I1(n17_adj_4962), .I2(n15_adj_4967), 
            .I3(n67420), .O(n67410));
    defparam i51682_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52593_4_lut (.I0(n25_adj_4958), .I1(n23_adj_4956), .I2(n21_adj_4964), 
            .I3(n67410), .O(n68321));
    defparam i52593_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52068_4_lut (.I0(n31_adj_4955), .I1(n29_adj_4954), .I2(n27_adj_4968), 
            .I3(n68321), .O(n67796));
    defparam i52068_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52710_4_lut (.I0(n37_adj_4953), .I1(n35_adj_4959), .I2(n33_adj_4960), 
            .I3(n67796), .O(n68438));
    defparam i52710_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52232_3_lut (.I0(n6_adj_4932), .I1(n436[10]), .I2(n21_adj_4964), 
            .I3(GND_net), .O(n67960));   // verilog/motorControl.v(54[23:39])
    defparam i52232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n436[9]), .I1(n436[21]), .I2(n43_adj_4952), 
            .I3(GND_net), .O(n16_adj_4972));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n436[4]), .I1(n436[8]), .I2(n17_adj_4962), 
            .I3(GND_net), .O(n8_adj_4973));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_4972), .I1(n436[22]), .I2(n45_adj_4951), 
            .I3(GND_net), .O(n24_adj_4974));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52233_3_lut (.I0(n67960), .I1(n436[11]), .I2(n23_adj_4956), 
            .I3(GND_net), .O(n67961));   // verilog/motorControl.v(54[23:39])
    defparam i52233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50759_4_lut (.I0(n43_adj_4952), .I1(n25_adj_4958), .I2(n23_adj_4956), 
            .I3(n66526), .O(n66487));
    defparam i50759_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51860_4_lut (.I0(n24_adj_4974), .I1(n8_adj_4973), .I2(n45_adj_4951), 
            .I3(n66485), .O(n67588));   // verilog/motorControl.v(54[23:39])
    defparam i51860_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51159_3_lut (.I0(n67961), .I1(n436[12]), .I2(n25_adj_4958), 
            .I3(GND_net), .O(n66887));   // verilog/motorControl.v(54[23:39])
    defparam i51159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52230_3_lut (.I0(n4_adj_9), .I1(n436[13]), .I2(n27_adj_4968), 
            .I3(GND_net), .O(n67958));   // verilog/motorControl.v(54[23:39])
    defparam i52230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52231_3_lut (.I0(n67958), .I1(n436[14]), .I2(n29_adj_4954), 
            .I3(GND_net), .O(n67959));   // verilog/motorControl.v(54[23:39])
    defparam i52231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50778_4_lut (.I0(n33_adj_4960), .I1(n31_adj_4955), .I2(n29_adj_4954), 
            .I3(n66514), .O(n66506));
    defparam i50778_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52627_4_lut (.I0(n30_adj_4971), .I1(n10_adj_4970), .I2(n35_adj_4959), 
            .I3(n66502), .O(n68355));   // verilog/motorControl.v(54[23:39])
    defparam i52627_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51161_3_lut (.I0(n67959), .I1(n436[15]), .I2(n31_adj_4955), 
            .I3(GND_net), .O(n66889));   // verilog/motorControl.v(54[23:39])
    defparam i51161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52811_4_lut (.I0(n66889), .I1(n68355), .I2(n35_adj_4959), 
            .I3(n66506), .O(n68539));   // verilog/motorControl.v(54[23:39])
    defparam i52811_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52812_3_lut (.I0(n68539), .I1(n436[18]), .I2(n37_adj_4953), 
            .I3(GND_net), .O(n68540));   // verilog/motorControl.v(54[23:39])
    defparam i52812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52767_3_lut (.I0(n68540), .I1(n436[19]), .I2(n39_adj_4950), 
            .I3(GND_net), .O(n68495));   // verilog/motorControl.v(54[23:39])
    defparam i52767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50761_4_lut (.I0(n43_adj_4952), .I1(n41_adj_4949), .I2(n39_adj_4950), 
            .I3(n68438), .O(n66489));
    defparam i50761_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52487_4_lut (.I0(n66887), .I1(n67588), .I2(n45_adj_4951), 
            .I3(n66487), .O(n68215));   // verilog/motorControl.v(54[23:39])
    defparam i52487_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51167_3_lut (.I0(n68495), .I1(n436[20]), .I2(n41_adj_4949), 
            .I3(GND_net), .O(n66895));   // verilog/motorControl.v(54[23:39])
    defparam i51167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52680_4_lut (.I0(n66895), .I1(n68215), .I2(n45_adj_4951), 
            .I3(n66489), .O(n68408));   // verilog/motorControl.v(54[23:39])
    defparam i52680_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52681_3_lut (.I0(n68408), .I1(n356[23]), .I2(n436[23]), .I3(GND_net), 
            .O(n68409));   // verilog/motorControl.v(54[23:39])
    defparam i52681_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5969_3_lut (.I0(control_update), .I1(n409), .I2(n68409), 
            .I3(GND_net), .O(n11610));   // verilog/motorControl.v(20[7:21])
    defparam i5969_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n365), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4985[6]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4452));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4451));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4450));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4976));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4977));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4978));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4979));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52236_3_lut (.I0(n32), .I1(n356[19]), .I2(n39_adj_4978), 
            .I3(GND_net), .O(n67964));   // verilog/motorControl.v(52[14:29])
    defparam i52236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52237_3_lut (.I0(n67964), .I1(n356[20]), .I2(n41_adj_4979), 
            .I3(GND_net), .O(n67965));   // verilog/motorControl.v(52[14:29])
    defparam i52237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51702_4_lut (.I0(n41_adj_4979), .I1(n39_adj_4978), .I2(n37_adj_4977), 
            .I3(n66569), .O(n67430));
    defparam i51702_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52180_3_lut (.I0(n34), .I1(n356[18]), .I2(n37_adj_4977), 
            .I3(GND_net), .O(n67908));   // verilog/motorControl.v(52[14:29])
    defparam i52180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51156_3_lut (.I0(n67965), .I1(n356[21]), .I2(n43_adj_4976), 
            .I3(GND_net), .O(n66884));   // verilog/motorControl.v(52[14:29])
    defparam i51156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52234_4_lut (.I0(n66884), .I1(n67908), .I2(n43_adj_4976), 
            .I3(n67430), .O(n67962));   // verilog/motorControl.v(52[14:29])
    defparam i52234_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52235_3_lut (.I0(n67962), .I1(n356[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n67963));   // verilog/motorControl.v(52[14:29])
    defparam i52235_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_23_i48_3_lut (.I0(n67963), .I1(PWMLimit[23]), .I2(n356[23]), 
            .I3(GND_net), .O(n409));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50952_4_lut (.I0(n356[6]), .I1(n356[5]), .I2(n382[6]), .I3(n382[5]), 
            .O(n66680));
    defparam i50952_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i51760_3_lut (.I0(n356[7]), .I1(n66680), .I2(n382[7]), .I3(GND_net), 
            .O(n67488));
    defparam i51760_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i27_rep_81_2_lut (.I0(n356[13]), .I1(n382[13]), 
            .I2(GND_net), .I3(GND_net), .O(n69904));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i27_rep_81_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51748_4_lut (.I0(n356[14]), .I1(n69904), .I2(n382[14]), .I3(n67488), 
            .O(n67476));
    defparam i51748_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i31_rep_75_2_lut (.I0(n365), .I1(n382[15]), .I2(GND_net), 
            .I3(GND_net), .O(n69898));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i31_rep_75_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35317_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n49235), 
            .I3(n20289[0]), .O(n4_adj_4918));   // verilog/motorControl.v(50[18:24])
    defparam i35317_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_980 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n20289[0]), 
            .I3(n49235), .O(n20265[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_980.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n382[7]), .I1(n382[16]), .I2(n356[16]), 
            .I3(GND_net), .O(n12_adj_4981));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50909_4_lut (.I0(n356[16]), .I1(n356[7]), .I2(n382[16]), 
            .I3(n382[7]), .O(n66637));
    defparam i50909_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n382[5]), .I1(n382[6]), .I2(n356[6]), 
            .I3(GND_net), .O(n10_adj_4486));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_4981), .I1(n382[17]), .I2(n356[17]), 
            .I3(GND_net), .O(n30_c));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50937_4_lut (.I0(n356[8]), .I1(n356[4]), .I2(n382[8]), .I3(n382[4]), 
            .O(n66665));
    defparam i50937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i35304_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n20265[0]));   // verilog/motorControl.v(50[18:24])
    defparam i35304_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i51756_3_lut (.I0(n356[9]), .I1(n66665), .I2(n382[9]), .I3(GND_net), 
            .O(n67484));
    defparam i51756_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i35306_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n49235));   // verilog/motorControl.v(50[18:24])
    defparam i35306_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_21_i21_rep_94_2_lut (.I0(n356[10]), .I1(n382[10]), 
            .I2(GND_net), .I3(GND_net), .O(n69917));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i21_rep_94_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51754_4_lut (.I0(n356[11]), .I1(n69917), .I2(n382[11]), .I3(n67484), 
            .O(n67482));
    defparam i51754_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i25_rep_89_2_lut (.I0(n356[12]), .I1(n382[12]), 
            .I2(GND_net), .I3(GND_net), .O(n69912));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i25_rep_89_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n382[9]), .I1(n382[21]), .I2(n356[21]), 
            .I3(GND_net), .O(n16_adj_4982));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50883_4_lut (.I0(n356[21]), .I1(n356[9]), .I2(n382[21]), 
            .I3(n382[9]), .O(n66611));
    defparam i50883_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n382[4]), .I1(n382[8]), .I2(n356[8]), 
            .I3(GND_net), .O(n8_adj_4489));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_4982), .I1(n382[22]), .I2(n356[22]), 
            .I3(GND_net), .O(n24_adj_4488));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50956_4_lut (.I0(n356[3]), .I1(n356[2]), .I2(n382[3]), .I3(n382[2]), 
            .O(n66684));
    defparam i50956_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i35422_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4983), 
            .I3(n20225[1]), .O(n6_adj_4907));   // verilog/motorControl.v(50[18:24])
    defparam i35422_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 LessThan_21_i9_rep_120_2_lut (.I0(n356[4]), .I1(n382[4]), .I2(GND_net), 
            .I3(GND_net), .O(n69943));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i9_rep_120_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50954_4_lut (.I0(n356[5]), .I1(n69943), .I2(n382[5]), .I3(n66684), 
            .O(n66682));
    defparam i50954_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i13_rep_113_2_lut (.I0(n356[6]), .I1(n382[6]), .I2(GND_net), 
            .I3(GND_net), .O(n69936));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i13_rep_113_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52108_4_lut (.I0(n356[7]), .I1(n69936), .I2(n382[7]), .I3(n66682), 
            .O(n67836));
    defparam i52108_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i17_rep_116_2_lut (.I0(n356[8]), .I1(n382[8]), .I2(GND_net), 
            .I3(GND_net), .O(n69939));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i17_rep_116_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_981 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n20225[1]), 
            .I3(n4_adj_4983), .O(n20165[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_981.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_982 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n20225[0]), 
            .I3(n49338), .O(n20165[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_982.LUT_INIT = 16'h8778;
    SB_LUT4 i51758_4_lut (.I0(n356[9]), .I1(n69939), .I2(n382[9]), .I3(n67836), 
            .O(n67486));
    defparam i51758_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i52379_4_lut (.I0(n356[11]), .I1(n69917), .I2(n382[11]), .I3(n67486), 
            .O(n68107));
    defparam i52379_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i50931_4_lut (.I0(n356[13]), .I1(n69912), .I2(n382[13]), .I3(n68107), 
            .O(n66659));
    defparam i50931_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35414_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n49338), 
            .I3(n20225[0]), .O(n4_adj_4983));   // verilog/motorControl.v(50[18:24])
    defparam i35414_3_lut_4_lut.LUT_INIT = 16'hf880;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2873, pwm_out, clk32MHz, GND_net, \pwm_counter[21] , 
            \pwm_counter[22] , pwm_setpoint, reset, n45, n43, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input n2873;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    output \pwm_counter[21] ;
    output \pwm_counter[22] ;
    input [23:0]pwm_setpoint;
    input reset;
    input n45;
    input n43;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_577;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n59301, n22, n15, n20, n24, n19, n48, n39, n41, n29, 
        n31, n37, n23, n25, n35, n11, n13, n15_adj_4445, n27, 
        n33, n9, n17, n19_adj_4446, n21, n66227, n66208, n56822, 
        n12, n30, n66262, n67176, n67166, n68293, n67694, n68422, 
        n55824, n55852, n55874, n55902, n55930, n55958, n55982, 
        n56020, n56064, n56102, n56142, n56186, n56224, n56264, 
        n56304, n56332, n56364, n56426, n56544, n56694, n56824, 
        n56826, n56828, n6, n68051, n68052, n16, n24_adj_4447, 
        n66136, n8, n66127, n67570, n66832, n4, n67688, n67689, 
        n66187, n10, n66176, n68287, n66834, n68442, n68443, n68433, 
        n66144, n68193, n66840, n68402, n50800, n50799, n50798, 
        n50797, n50796, n50795, n50794, n50793, n50792, n50791, 
        n50790, n50789, n50788, n50787, n50786, n50785, n50784, 
        n50783, n50782, n50781, n50780, n50779, n50778;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2873), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n59301));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(\pwm_counter[21] ), .I1(pwm_counter[15]), .I2(pwm_counter[18]), 
            .I3(pwm_counter[16]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n59301), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[17]), .I1(\pwm_counter[22] ), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22), .I2(pwm_counter[20]), .I3(pwm_counter[13]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[19]), .I1(pwm_counter[14]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4445));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4446));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50499_4_lut (.I0(n21), .I1(n19_adj_4446), .I2(n17), .I3(n9), 
            .O(n66227));
    defparam i50499_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50480_4_lut (.I0(n27), .I1(n15_adj_4445), .I2(n13), .I3(n11), 
            .O(n66208));
    defparam i50480_4_lut.LUT_INIT = 16'haaab;
    SB_DFFR pwm_counter_1939__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n56822), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51448_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n66262), 
            .O(n67176));
    defparam i51448_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51438_4_lut (.I0(n19_adj_4446), .I1(n17), .I2(n15_adj_4445), 
            .I3(n67176), .O(n67166));
    defparam i51438_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52565_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n67166), 
            .O(n68293));
    defparam i52565_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51966_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n68293), 
            .O(n67694));
    defparam i51966_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52694_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67694), 
            .O(n68422));
    defparam i52694_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFR pwm_counter_1939__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n55824), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i22 (.Q(\pwm_counter[22] ), .C(clk32MHz), 
            .D(n55852), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i21 (.Q(\pwm_counter[21] ), .C(clk32MHz), 
            .D(n55874), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n55902), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n55930), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n55958), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n55982), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n56020), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n56064), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n56102), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n56142), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n56186), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n56224), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n56264), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n56304), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n56332), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n56364), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n56426), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n56544), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n56694), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n56824), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n56826), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n56828), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i52323_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n68051));   // verilog/pwm.v(21[8:24])
    defparam i52323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52324_3_lut (.I0(n68051), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n68052));   // verilog/pwm.v(21[8:24])
    defparam i52324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4447));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50408_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n66227), 
            .O(n66136));
    defparam i50408_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51842_4_lut (.I0(n24_adj_4447), .I1(n8), .I2(n45), .I3(n66127), 
            .O(n67570));   // verilog/pwm.v(21[8:24])
    defparam i51842_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51104_3_lut (.I0(n68052), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n66832));   // verilog/pwm.v(21[8:24])
    defparam i51104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51960_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n67688));   // verilog/pwm.v(21[8:24])
    defparam i51960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51961_3_lut (.I0(n67688), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n67689));   // verilog/pwm.v(21[8:24])
    defparam i51961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50459_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n66208), 
            .O(n66187));
    defparam i50459_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52559_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n66176), 
            .O(n68287));   // verilog/pwm.v(21[8:24])
    defparam i52559_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51106_3_lut (.I0(n67689), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n66834));   // verilog/pwm.v(21[8:24])
    defparam i51106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52714_4_lut (.I0(n66834), .I1(n68287), .I2(n35), .I3(n66187), 
            .O(n68442));   // verilog/pwm.v(21[8:24])
    defparam i52714_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52715_3_lut (.I0(n68442), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n68443));   // verilog/pwm.v(21[8:24])
    defparam i52715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52705_3_lut (.I0(n68443), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n68433));   // verilog/pwm.v(21[8:24])
    defparam i52705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50416_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n68422), 
            .O(n66144));
    defparam i50416_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52465_4_lut (.I0(n66832), .I1(n67570), .I2(n45), .I3(n66136), 
            .O(n68193));   // verilog/pwm.v(21[8:24])
    defparam i52465_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51112_3_lut (.I0(n68433), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n66840));   // verilog/pwm.v(21[8:24])
    defparam i51112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52674_4_lut (.I0(n66840), .I1(n68193), .I2(n45), .I3(n66144), 
            .O(n68402));   // verilog/pwm.v(21[8:24])
    defparam i52674_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52675_3_lut (.I0(n68402), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i52675_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 pwm_counter_1939_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n50800), .O(n55824)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1939_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[22] ), 
            .I3(n50799), .O(n55852)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_24 (.CI(n50799), .I0(GND_net), .I1(\pwm_counter[22] ), 
            .CO(n50800));
    SB_LUT4 pwm_counter_1939_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[21] ), 
            .I3(n50798), .O(n55874)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_23 (.CI(n50798), .I0(GND_net), .I1(\pwm_counter[21] ), 
            .CO(n50799));
    SB_LUT4 pwm_counter_1939_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n50797), .O(n55902)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_22 (.CI(n50797), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n50798));
    SB_LUT4 pwm_counter_1939_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n50796), .O(n55930)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_21 (.CI(n50796), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n50797));
    SB_LUT4 pwm_counter_1939_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n50795), .O(n55958)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_20 (.CI(n50795), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n50796));
    SB_LUT4 pwm_counter_1939_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n50794), .O(n55982)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_19 (.CI(n50794), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n50795));
    SB_LUT4 pwm_counter_1939_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n50793), .O(n56020)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_18 (.CI(n50793), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n50794));
    SB_LUT4 pwm_counter_1939_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n50792), .O(n56064)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_17 (.CI(n50792), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n50793));
    SB_LUT4 pwm_counter_1939_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n50791), .O(n56102)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_16 (.CI(n50791), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n50792));
    SB_LUT4 pwm_counter_1939_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n50790), .O(n56142)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_15 (.CI(n50790), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n50791));
    SB_LUT4 pwm_counter_1939_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n50789), .O(n56186)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_14 (.CI(n50789), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n50790));
    SB_LUT4 pwm_counter_1939_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n50788), .O(n56224)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_13 (.CI(n50788), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n50789));
    SB_LUT4 pwm_counter_1939_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n50787), .O(n56264)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_12 (.CI(n50787), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n50788));
    SB_LUT4 pwm_counter_1939_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n50786), .O(n56304)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_11 (.CI(n50786), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n50787));
    SB_LUT4 pwm_counter_1939_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n50785), .O(n56332)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_10 (.CI(n50785), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n50786));
    SB_LUT4 pwm_counter_1939_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n50784), .O(n56364)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_9 (.CI(n50784), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n50785));
    SB_LUT4 pwm_counter_1939_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n50783), .O(n56426)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_8 (.CI(n50783), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n50784));
    SB_LUT4 pwm_counter_1939_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n50782), .O(n56544)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_7 (.CI(n50782), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n50783));
    SB_LUT4 pwm_counter_1939_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n50781), .O(n56694)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_6 (.CI(n50781), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n50782));
    SB_LUT4 pwm_counter_1939_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n50780), .O(n56824)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_5 (.CI(n50780), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n50781));
    SB_LUT4 pwm_counter_1939_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n50779), .O(n56826)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_4 (.CI(n50779), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n50780));
    SB_LUT4 pwm_counter_1939_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n50778), .O(n56828)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_3 (.CI(n50778), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n50779));
    SB_LUT4 pwm_counter_1939_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n56822)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n50778));
    SB_LUT4 i50534_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n66262));   // verilog/pwm.v(21[8:24])
    defparam i50534_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50399_2_lut_4_lut (.I0(pwm_setpoint[21]), .I1(\pwm_counter[21] ), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n66127));
    defparam i50399_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(\pwm_counter[21] ), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50448_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n66176));
    defparam i50448_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (enable_slow_N_4211, ready_prev, clk16MHz, n5773, \state[2] , 
            \state[0] , n57392, GND_net, n3, \state[1] , \state[0]_adj_4 , 
            data, ID, n25471, n28027, n29676, rw, n56774, data_ready, 
            n56368, n56570, baudrate, n30440, n30438, n30437, n30436, 
            n30435, n30434, n30433, n30432, n42792, n25612, \state_7__N_3916[0] , 
            scl_enable, VCC_net, \state_7__N_4108[0] , \saved_addr[0] , 
            \state_7__N_4124[3] , n10, n6428, n10_adj_5, n29683, n30523, 
            n8, n30246, n30245, n30244, n30243, n30242, n30241, 
            n30240, scl, sda_enable, n65775, n25595, n25600, sda_out, 
            n4, n4_adj_6, n42890) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output enable_slow_N_4211;
    output ready_prev;
    input clk16MHz;
    output [0:0]n5773;
    output \state[2] ;
    output \state[0] ;
    output n57392;
    input GND_net;
    output n3;
    output \state[1] ;
    output \state[0]_adj_4 ;
    output [7:0]data;
    output [7:0]ID;
    output n25471;
    output n28027;
    input n29676;
    output rw;
    input n56774;
    output data_ready;
    input n56368;
    input n56570;
    output [31:0]baudrate;
    input n30440;
    input n30438;
    input n30437;
    input n30436;
    input n30435;
    input n30434;
    input n30433;
    input n30432;
    output n42792;
    output n25612;
    input \state_7__N_3916[0] ;
    output scl_enable;
    input VCC_net;
    output \state_7__N_4108[0] ;
    output \saved_addr[0] ;
    input \state_7__N_4124[3] ;
    output n10;
    output n6428;
    output n10_adj_5;
    input n29683;
    input n30523;
    input n8;
    input n30246;
    input n30245;
    input n30244;
    input n30243;
    input n30242;
    input n30241;
    input n30240;
    output scl;
    output sda_enable;
    output n65775;
    output n25595;
    output n25600;
    output sda_out;
    output n4;
    output n4_adj_6;
    output n42890;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire enable;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    wire [15:0]delay_counter_15__N_3954;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    wire [15:0]n5113;
    
    wire n49794, n49793;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n51243, n47670, n49792, n49791, n49790, n6687, n49789, 
        n47643, n6686, n49788, n6685, n49787, n6684, n49786, n6683, 
        n49785, n49784, n6681, n49783, n49782, n49781, n49780, 
        n47662, n15, n30465, n30467, n30468, n30469, n30470, n30471, 
        n30472, n29670;
    wire [2:0]n17;
    
    wire n27799, n29186, n52217, n30464, n30463, n30462, n30461, 
        n30460, n30459, n30458, n30457, n30456, n30455, n30454, 
        n30453, n56640, n56656, n56638, n56642, n30448, n30447, 
        n30446, n30445, n30444, n30443, n30442, n30441;
    wire [7:0]state_7__N_3883;
    
    wire n60233, n6, n27727, n47640, n62678, n4_c, n4_adj_4441, 
        n65784, n28, n26, n27, n25;
    
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4211));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5773[0]), .R(\state[2] ));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(state[3]), .I2(state[2]), 
            .I3(state[1]), .O(n57392));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_1103_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5113[11]), 
            .I3(n49794), .O(delay_counter_15__N_3954[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1103_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5113[11]), 
            .I3(n49793), .O(delay_counter_15__N_3954[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_16 (.CI(n49793), .I0(delay_counter[14]), .I1(n5113[11]), 
            .CO(n49794));
    SB_LUT4 i2_3_lut (.I0(byte_counter[2]), .I1(n51243), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n47670));
    defparam i2_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 add_1103_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5113[11]), 
            .I3(n49792), .O(delay_counter_15__N_3954[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_15 (.CI(n49792), .I0(delay_counter[13]), .I1(n5113[11]), 
            .CO(n49793));
    SB_LUT4 add_1103_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5113[11]), 
            .I3(n49791), .O(delay_counter_15__N_3954[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_14 (.CI(n49791), .I0(delay_counter[12]), .I1(n5113[11]), 
            .CO(n49792));
    SB_LUT4 add_1103_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5113[11]), 
            .I3(n49790), .O(delay_counter_15__N_3954[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_13 (.CI(n49790), .I0(delay_counter[11]), .I1(n5113[11]), 
            .CO(n49791));
    SB_LUT4 add_1103_12_lut (.I0(n47643), .I1(delay_counter[10]), .I2(n5113[11]), 
            .I3(n49789), .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_12 (.CI(n49789), .I0(delay_counter[10]), .I1(n5113[11]), 
            .CO(n49790));
    SB_LUT4 add_1103_11_lut (.I0(n47643), .I1(delay_counter[9]), .I2(n5113[11]), 
            .I3(n49788), .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_11 (.CI(n49788), .I0(delay_counter[9]), .I1(n5113[11]), 
            .CO(n49789));
    SB_LUT4 add_1103_10_lut (.I0(n47643), .I1(delay_counter[8]), .I2(n5113[11]), 
            .I3(n49787), .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_10 (.CI(n49787), .I0(delay_counter[8]), .I1(n5113[11]), 
            .CO(n49788));
    SB_LUT4 add_1103_9_lut (.I0(n47643), .I1(delay_counter[7]), .I2(n5113[11]), 
            .I3(n49786), .O(n6684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_9 (.CI(n49786), .I0(delay_counter[7]), .I1(n5113[11]), 
            .CO(n49787));
    SB_LUT4 add_1103_8_lut (.I0(n47643), .I1(delay_counter[6]), .I2(n5113[11]), 
            .I3(n49785), .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_8 (.CI(n49785), .I0(delay_counter[6]), .I1(n5113[11]), 
            .CO(n49786));
    SB_LUT4 add_1103_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5113[11]), 
            .I3(n49784), .O(delay_counter_15__N_3954[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_7 (.CI(n49784), .I0(delay_counter[5]), .I1(n5113[11]), 
            .CO(n49785));
    SB_LUT4 add_1103_6_lut (.I0(n47643), .I1(delay_counter[4]), .I2(n5113[11]), 
            .I3(n49783), .O(n6681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_6 (.CI(n49783), .I0(delay_counter[4]), .I1(n5113[11]), 
            .CO(n49784));
    SB_LUT4 add_1103_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5113[11]), 
            .I3(n49782), .O(delay_counter_15__N_3954[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_5 (.CI(n49782), .I0(delay_counter[3]), .I1(n5113[11]), 
            .CO(n49783));
    SB_LUT4 add_1103_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5113[11]), 
            .I3(n49781), .O(delay_counter_15__N_3954[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_4 (.CI(n49781), .I0(delay_counter[2]), .I1(n5113[11]), 
            .CO(n49782));
    SB_LUT4 i1_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n3));   // verilog/eeprom.v(30[11:23])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13_2_lut (.I0(\state[2] ), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n47643));
    defparam i13_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 add_1103_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5113[11]), 
            .I3(n49780), .O(delay_counter_15__N_3954[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_3 (.CI(n49780), .I0(delay_counter[1]), .I1(n5113[11]), 
            .CO(n49781));
    SB_LUT4 add_1103_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5113[11]), 
            .I3(GND_net), .O(delay_counter_15__N_3954[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5113[11]), 
            .CO(n49780));
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(\state[0]_adj_4 ), .I2(n3), 
            .I3(\state[2] ), .O(n47662));
    defparam i1_4_lut.LUT_INIT = 16'h0144;
    SB_LUT4 i16389_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(ID[7]), .O(n30465));
    defparam i16389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i52959_2_lut (.I0(n25471), .I1(enable_slow_N_4211), .I2(GND_net), 
            .I3(GND_net), .O(n5113[11]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i52959_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16391_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(ID[6]), .O(n30467));
    defparam i16391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16392_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(ID[5]), .O(n30468));
    defparam i16392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16393_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(ID[4]), .O(n30469));
    defparam i16393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16394_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(ID[3]), .O(n30470));
    defparam i16394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16395_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(ID[2]), .O(n30471));
    defparam i16395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16396_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(ID[1]), .O(n30472));
    defparam i16396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15594_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(ID[0]), .O(n29670));
    defparam i15594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_954 (.I0(byte_counter[1]), .I1(n51243), .I2(byte_counter[2]), 
            .I3(byte_counter[0]), .O(n28027));
    defparam i2_3_lut_4_lut_adj_954.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut (.I0(byte_counter[1]), .I1(n51243), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n15));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n29676));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n56774));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29670));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i2 (.Q(\state[2] ), .C(clk16MHz), .D(n56368));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_1945__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27799), .D(n17[1]), .R(n29186));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1945__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27799), .D(n17[2]), .R(n29186));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1945__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27799), .D(n52217), .R(n29186));   // verilog/eeprom.v(68[25:39])
    SB_DFF state_i0 (.Q(\state[0]_adj_4 ), .C(clk16MHz), .D(n56570));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30472));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30471));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30470));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30469));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30468));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30467));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30465));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30464));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30463));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30462));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30461));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30460));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30459));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30458));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30457));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30456));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30455));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30454));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30453));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n56640));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n56656));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n56638));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n56642));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30448));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30447));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30446));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30445));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30444));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30443));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30442));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30441));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30440));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30438));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30437));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30436));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30435));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30434));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30433));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30432));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i28824_2_lut (.I0(enable_slow_N_4211), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n42792));
    defparam i28824_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(n60233), .D(state_7__N_3883[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut (.I0(\state[0]_adj_4 ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(ready_prev), .I1(n57392), .I2(\state[2] ), .I3(n6), 
            .O(n51243));
    defparam i4_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\state[0]_adj_4 ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n25612));   // verilog/eeprom.v(38[3] 80[10])
    defparam i1_2_lut_adj_955.LUT_INIT = 16'heeee;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27727), .D(delay_counter_15__N_3954[15]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27727), .D(delay_counter_15__N_3954[14]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27727), .D(delay_counter_15__N_3954[13]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27727), .D(delay_counter_15__N_3954[12]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27727), .D(delay_counter_15__N_3954[11]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27727), .D(n6687), .S(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27727), 
            .D(n6686), .S(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27727), 
            .D(n6685), .S(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27727), 
            .D(n6684), .S(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27727), 
            .D(n6683), .S(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27727), 
            .D(delay_counter_15__N_3954[5]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27727), 
            .D(n6681), .S(n47640));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27727), 
            .D(delay_counter_15__N_3954[3]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27727), 
            .D(delay_counter_15__N_3954[2]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27727), 
            .D(delay_counter_15__N_3954[1]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27727), 
            .D(delay_counter_15__N_3954[0]), .R(n47662));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i46960_2_lut_3_lut (.I0(state[1]), .I1(state[2]), .I2(\state[0] ), 
            .I3(GND_net), .O(n62678));   // verilog/eeprom.v(55[12:28])
    defparam i46960_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_4_lut (.I0(state[1]), .I1(state[2]), .I2(\state[0] ), 
            .I3(state[3]), .O(n4_c));   // verilog/eeprom.v(55[12:28])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hffc1;
    SB_LUT4 i1_4_lut_adj_956 (.I0(\state[2] ), .I1(\state[1] ), .I2(\state_7__N_3916[0] ), 
            .I3(\state[0]_adj_4 ), .O(n4_adj_4441));
    defparam i1_4_lut_adj_956.LUT_INIT = 16'hbbba;
    SB_LUT4 i50939_4_lut (.I0(n62678), .I1(n25471), .I2(\state[1] ), .I3(state[3]), 
            .O(n65784));
    defparam i50939_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n65784), .I1(n4_adj_4441), .I2(n42792), .I3(\state[0]_adj_4 ), 
            .O(n60233));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i1_4_lut_adj_957 (.I0(n3), .I1(\state[0]_adj_4 ), .I2(\state[2] ), 
            .I3(\state[1] ), .O(state_7__N_3883[1]));
    defparam i1_4_lut_adj_957.LUT_INIT = 16'hf31c;
    SB_LUT4 i2_3_lut_4_lut_adj_958 (.I0(\state[1] ), .I1(\state_7__N_3916[0] ), 
            .I2(\state[0]_adj_4 ), .I3(\state[2] ), .O(n29186));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut_adj_958.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_4_lut_adj_959 (.I0(\state[1] ), .I1(\state_7__N_3916[0] ), 
            .I2(\state[0]_adj_4 ), .I3(\state[2] ), .O(n27799));   // verilog/eeprom.v(68[25:39])
    defparam i1_4_lut_4_lut_adj_959.LUT_INIT = 16'h00a4;
    SB_LUT4 i35388_2_lut_3_lut_4_lut (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i35388_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i35395_3_lut_4_lut (.I0(n42792), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i35395_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i33688_4_lut_4_lut (.I0(\state[1] ), .I1(n3), .I2(\state[2] ), 
            .I3(\state[0]_adj_4 ), .O(n47640));
    defparam i33688_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 i25_4_lut_4_lut (.I0(\state[1] ), .I1(n3), .I2(\state[0]_adj_4 ), 
            .I3(\state[2] ), .O(n27727));
    defparam i25_4_lut_4_lut.LUT_INIT = 16'h015a;
    SB_LUT4 i1_2_lut_3_lut_adj_960 (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n52217));
    defparam i1_2_lut_3_lut_adj_960.LUT_INIT = 16'hd2d2;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n25471));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1450_Mux_0_i3_4_lut (.I0(\state[0]_adj_4 ), .I1(enable_slow_N_4211), 
            .I2(\state[1] ), .I3(n25471), .O(n5773[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1450_Mux_0_i3_4_lut.LUT_INIT = 16'h0a4a;
    SB_LUT4 i16388_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(baudrate[0]), .O(n30464));   // verilog/eeprom.v(68[25:39])
    defparam i16388_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16381_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(baudrate[7]), .O(n30457));   // verilog/eeprom.v(68[25:39])
    defparam i16381_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16382_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(baudrate[6]), .O(n30458));   // verilog/eeprom.v(68[25:39])
    defparam i16382_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16383_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(baudrate[5]), .O(n30459));   // verilog/eeprom.v(68[25:39])
    defparam i16383_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16384_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(baudrate[4]), .O(n30460));   // verilog/eeprom.v(68[25:39])
    defparam i16384_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16385_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(baudrate[3]), .O(n30461));   // verilog/eeprom.v(68[25:39])
    defparam i16385_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16386_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(baudrate[2]), .O(n30462));   // verilog/eeprom.v(68[25:39])
    defparam i16386_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16387_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(baudrate[1]), .O(n30463));   // verilog/eeprom.v(68[25:39])
    defparam i16387_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16377_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[3]), 
            .I3(baudrate[11]), .O(n30453));   // verilog/eeprom.v(68[25:39])
    defparam i16377_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[7]), 
            .I3(baudrate[15]), .O(n56642));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_961 (.I0(byte_counter[0]), .I1(n47670), 
            .I2(data[6]), .I3(baudrate[14]), .O(n56638));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_961.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_962 (.I0(byte_counter[0]), .I1(n47670), 
            .I2(data[5]), .I3(baudrate[13]), .O(n56656));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_962.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_963 (.I0(byte_counter[0]), .I1(n47670), 
            .I2(data[4]), .I3(baudrate[12]), .O(n56640));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_963.LUT_INIT = 16'hfb40;
    SB_LUT4 i16379_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[1]), 
            .I3(baudrate[9]), .O(n30455));   // verilog/eeprom.v(68[25:39])
    defparam i16379_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16378_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[2]), 
            .I3(baudrate[10]), .O(n30454));   // verilog/eeprom.v(68[25:39])
    defparam i16378_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16380_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[0]), 
            .I3(baudrate[8]), .O(n30456));   // verilog/eeprom.v(68[25:39])
    defparam i16380_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16372_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[0]), 
            .I3(baudrate[16]), .O(n30448));   // verilog/eeprom.v(68[25:39])
    defparam i16372_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16365_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[7]), 
            .I3(baudrate[23]), .O(n30441));   // verilog/eeprom.v(68[25:39])
    defparam i16365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16366_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[6]), 
            .I3(baudrate[22]), .O(n30442));   // verilog/eeprom.v(68[25:39])
    defparam i16366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16367_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[5]), 
            .I3(baudrate[21]), .O(n30443));   // verilog/eeprom.v(68[25:39])
    defparam i16367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16368_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[4]), 
            .I3(baudrate[20]), .O(n30444));   // verilog/eeprom.v(68[25:39])
    defparam i16368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16369_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[3]), 
            .I3(baudrate[19]), .O(n30445));   // verilog/eeprom.v(68[25:39])
    defparam i16369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16370_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[2]), 
            .I3(baudrate[18]), .O(n30446));   // verilog/eeprom.v(68[25:39])
    defparam i16370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16371_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47670), .I2(data[1]), 
            .I3(baudrate[17]), .O(n30447));   // verilog/eeprom.v(68[25:39])
    defparam i16371_3_lut_4_lut.LUT_INIT = 16'hf780;
    i2c_controller i2c (.clk16MHz(clk16MHz), .scl_enable(scl_enable), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\state_7__N_4108[0] (\state_7__N_4108[0] ), 
            .\state[3] (state[3]), .\state[1] (state[1]), .\state[0] (\state[0] ), 
            .\state[2] (state[2]), .\saved_addr[0] (\saved_addr[0] ), .enable_slow_N_4211(enable_slow_N_4211), 
            .\state_7__N_4124[3] (\state_7__N_4124[3] ), .enable(enable), 
            .n10(n10), .n6428(n6428), .n10_adj_1(n10_adj_5), .n29683(n29683), 
            .n4(n4_c), .n30523(n30523), .data({data}), .n8(n8), .n30246(n30246), 
            .n30245(n30245), .n30244(n30244), .n30243(n30243), .n30242(n30242), 
            .n30241(n30241), .n30240(n30240), .scl(scl), .sda_enable(sda_enable), 
            .n65775(n65775), .n25595(n25595), .n25600(n25600), .sda_out(sda_out), 
            .n4_adj_2(n4), .n4_adj_3(n4_adj_6), .n42890(n42890)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (clk16MHz, scl_enable, VCC_net, GND_net, \state_7__N_4108[0] , 
            \state[3] , \state[1] , \state[0] , \state[2] , \saved_addr[0] , 
            enable_slow_N_4211, \state_7__N_4124[3] , enable, n10, n6428, 
            n10_adj_1, n29683, n4, n30523, data, n8, n30246, n30245, 
            n30244, n30243, n30242, n30241, n30240, scl, sda_enable, 
            n65775, n25595, n25600, sda_out, n4_adj_2, n4_adj_3, 
            n42890) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output scl_enable;
    input VCC_net;
    input GND_net;
    output \state_7__N_4108[0] ;
    output \state[3] ;
    output \state[1] ;
    output \state[0] ;
    output \state[2] ;
    output \saved_addr[0] ;
    output enable_slow_N_4211;
    input \state_7__N_4124[3] ;
    input enable;
    output n10;
    output n6428;
    output n10_adj_1;
    input n29683;
    input n4;
    input n30523;
    output [7:0]data;
    input n8;
    input n30246;
    input n30245;
    input n30244;
    input n30243;
    input n30242;
    input n30241;
    input n30240;
    output scl;
    output sda_enable;
    output n65775;
    output n25595;
    output n25600;
    output sda_out;
    output n4_adj_2;
    output n4_adj_3;
    output n42890;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire i2c_clk_N_4197, scl_enable_N_4198;
    wire [7:0]n119;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n49801, n49800, n49799, n49798, n49797, n49796, n49795, 
        enable_slow_N_4210, n27787, n28, n68643, n11, n58282, n27780;
    wire [1:0]n6491;
    
    wire n56624, n27782, n11_adj_4428, n11_adj_4429, n11_adj_4430, 
        n4_c, n43046, n9, state_7__N_4107, n6421, n42942, n5, 
        n12, n15, n65786, n6758, n27982;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n29169, n50933, n50932, n50931, n50930, n50929, n28927, 
        n43552, n43334, n60458, n60061, n59245, n59989, sda_out_adj_4433, 
        n11_adj_4434, n10_adj_4435;
    
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4197));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4198));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n49801), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n49800), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n49800), .I0(counter[6]), .I1(VCC_net), 
            .CO(n49801));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n49799), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n49799), .I0(counter[5]), .I1(VCC_net), 
            .CO(n49800));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n49798), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n49798), .I0(counter[4]), .I1(VCC_net), 
            .CO(n49799));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n49797), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n49797), .I0(counter[3]), .I1(VCC_net), 
            .CO(n49798));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n49796), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n49796), .I0(counter[2]), .I1(VCC_net), 
            .CO(n49797));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n49795), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4108[0] ), .C(clk16MHz), .E(n27787), 
            .D(enable_slow_N_4210));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_CARRY sub_39_add_2_3 (.CI(n49795), .I0(counter[1]), .I1(VCC_net), 
            .CO(n49796));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n49795));
    SB_LUT4 i1_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i52915_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n68643));
    defparam i52915_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_945 (.I0(n11), .I1(n68643), .I2(n28), .I3(n58282), 
            .O(n27780));
    defparam i1_4_lut_adj_945.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1730_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6491[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1730_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i29574_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n58282));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i29574_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n11), .I1(n58282), .I2(\state[3] ), .I3(\state[1] ), 
            .O(n56624));
    defparam i3_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_946 (.I0(n11), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n58282), .O(n27782));
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h0a22;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4428));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4429));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52952_2_lut (.I0(\state_7__N_4108[0] ), .I1(enable_slow_N_4211), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4210));   // verilog/i2c_controller.v(62[6:32])
    defparam i52952_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_947 (.I0(\state_7__N_4124[3] ), .I1(n11_adj_4430), 
            .I2(n11), .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h2a2f;
    SB_LUT4 i53438_2_lut (.I0(\state_7__N_4124[3] ), .I1(n11_adj_4430), 
            .I2(GND_net), .I3(GND_net), .O(n43046));
    defparam i53438_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_141_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_141_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i52934_4_lut (.I0(state_7__N_4107), .I1(n6421), .I2(n11_adj_4429), 
            .I3(n42942), .O(n6428));
    defparam i52934_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n11_adj_4428), .I1(n11_adj_4430), .I2(\state_7__N_4124[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h5755;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_1));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_1), 
            .O(n6421));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29683));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i50070_2_lut (.I0(n15), .I1(\state_7__N_4124[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n65786));
    defparam i50070_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14_4_lut (.I0(n6421), .I1(n65786), .I2(n6758), .I3(n4), 
            .O(n27982));
    defparam i14_4_lut.LUT_INIT = 16'h303a;
    SB_DFFSR counter2_1954_1955__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29169));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29169));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29169));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29169));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29169));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 counter2_1954_1955_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n50933), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1954_1955_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n50932), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_6 (.CI(n50932), .I0(GND_net), .I1(counter2[4]), 
            .CO(n50933));
    SB_LUT4 counter2_1954_1955_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n50931), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_5 (.CI(n50931), .I0(GND_net), .I1(counter2[3]), 
            .CO(n50932));
    SB_LUT4 counter2_1954_1955_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n50930), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_4 (.CI(n50930), .I0(GND_net), .I1(counter2[2]), 
            .CO(n50931));
    SB_LUT4 counter2_1954_1955_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n50929), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_3 (.CI(n50929), .I0(GND_net), .I1(counter2[1]), 
            .CO(n50930));
    SB_LUT4 counter2_1954_1955_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n50929));
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27982), .D(n119[1]), 
            .S(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27982), .D(n119[2]), 
            .S(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27982), .D(n119[3]), 
            .R(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27982), .D(n119[4]), 
            .R(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27982), .D(n119[5]), 
            .R(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27982), .D(n119[6]), 
            .R(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27982), .D(n119[7]), 
            .R(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6428), .D(n5), 
            .S(n43552));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6428), .D(n43046), 
            .S(n43334));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6428), .D(n60458), 
            .S(n60061));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1954_1955__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29169));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30523));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n30246));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n30245));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n30244));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n30243));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n30242));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n30241));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n30240));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i28846_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i28846_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27782), 
            .D(n59245), .S(n56624));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4433), .C(i2c_clk), .E(n27780), 
            .D(n59989), .S(n56624));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27982), .D(n119[0]), 
            .S(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i50189_3_lut_4_lut (.I0(n11_adj_4429), .I1(n11_adj_4434), .I2(enable_slow_N_4211), 
            .I3(\state_7__N_4108[0] ), .O(n65775));
    defparam i50189_3_lut_4_lut.LUT_INIT = 16'h0888;
    SB_LUT4 i53513_3_lut_4_lut (.I0(n11_adj_4429), .I1(n11_adj_4434), .I2(n15), 
            .I3(n6428), .O(n43552));
    defparam i53513_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i29436_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_4107));
    defparam i29436_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9), .O(n60458));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf0f4;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n25595));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_949 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n25600));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_949.LUT_INIT = 16'hfefe;
    SB_LUT4 i53511_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4434), 
            .I3(n6428), .O(n43334));   // verilog/i2c_controller.v(151[5:14])
    defparam i53511_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4435));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4435), .I2(counter2[0]), 
            .I3(GND_net), .O(n29169));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_1517_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));
    defparam equal_1517_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29169), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4197));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2431_2_lut (.I0(sda_out_adj_4433), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2431_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14851_2_lut_4_lut (.I0(n27982), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n28927));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14851_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i28973_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n42942));
    defparam i28973_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i53503_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6428), .O(n60061));
    defparam i53503_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_950 (.I0(enable), .I1(\state_7__N_4108[0] ), 
            .I2(enable_slow_N_4211), .I3(GND_net), .O(n27787));
    defparam i1_2_lut_3_lut_adj_950.LUT_INIT = 16'haeae;
    SB_LUT4 equal_351_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_351_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_349_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_349_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28922_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n42890));
    defparam i28922_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_951 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n59245));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_951.LUT_INIT = 16'h1110;
    SB_LUT4 i29467_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4198));   // verilog/i2c_controller.v(44[32:47])
    defparam i29467_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i52967_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(enable_slow_N_4211));   // verilog/i2c_controller.v(44[32:47])
    defparam i52967_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_4430));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut_adj_952 (.I0(\state[2] ), .I1(\state[3] ), .I2(n6491[1]), 
            .I3(\state[1] ), .O(n59989));   // verilog/i2c_controller.v(44[32:47])
    defparam i2_3_lut_4_lut_adj_952.LUT_INIT = 16'h1000;
    SB_LUT4 equal_272_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n15));   // verilog/i2c_controller.v(44[32:47])
    defparam equal_272_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_953 (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n6758));   // verilog/i2c_controller.v(44[32:47])
    defparam i1_2_lut_3_lut_adj_953.LUT_INIT = 16'h1010;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n11_adj_4434));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    
endmodule
