// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Jan 23 17:00:06 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    output SCL;   // verilog/TinyFPGA_B.v(21[10:13])
    input SDA /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, CLK_c, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c_0;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(42[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(88[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(89[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(125[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(126[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(127[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(128[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(129[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(131[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(132[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(133[22:35])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(163[22:33])
    wire [22:0]pwm_setpoint_22__N_3;
    
    wire RX_N_2;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n1929;
    wire [23:0]displacement_23__N_26;
    
    wire n6, n31239, n7, n31238, n15763, n31237;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n26561, n2649, n4774, n4, n15762, n15619, n4772, n15761, 
        n15760, n15759, n15758, n15757;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n5, n4_adj_4763, n15756, n15755, n15754, n15753, n15752, 
        n3, n4_adj_4764, n5_adj_4765, n6_adj_4766, n7_adj_4767, n8, 
        n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
        n19, n20, n21, n22, n23, n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n122, n123, n4_adj_4768, n25997, n771, n5_adj_4769, n27965, 
        n29876, n29875, n29874, n29873, n29872, n29871, n29870, 
        n29869, n29868, n29867, n29866, n14291, n29865, n29864, 
        n29863, n29862, n29861, n29860, n14259, n29859, n29858, 
        n22558, n22557, n22556, n29857, n29856, n30633, n29855, 
        n22340, n22339, n22555, n29854, n22338, n22337, n22554;
    wire [31:0]\FRAME_MATCHER.state_31__N_2672 ;
    
    wire n22336, n22553, n22552, n25861, n22551, n18753, n29839, 
        n22335, n22550, n22334, n22333, n10_adj_4770, n4452, n22332, 
        n22331, n22330, n22329, n22549, n22328, n22548, n22327, 
        n22547, n22326, n22546, n19323, n22545, n22544, n22543, 
        n22542, n14279, n14288, n22325, n22324, n22541, n22540, 
        n22539, n22538, n22537, n22536, n22323, n26611, n16227, 
        n16226, n16225, n16224, n16223, n16222, n16221, n16220, 
        n16219, n16218, n16217, n16216, n16215, n16214, n16213, 
        n16212, n16211, n16210, n16209, n16208, n16207, n16206, 
        n16205, n16204, n16203, n16202, n16201, n16200, n16199, 
        n16198, n16197, n16196, n16195, n16194, n16193, n16192, 
        n16191, n16190, n16189, n16185, n16183, n16178, n16177, 
        n16176, n16175, n16174, n16173, n16172, n16171, n16170, 
        n16169, n16168, n16167, n16166, n16165, n16164, n16163, 
        n16162, n16161, n16160, n16159, n16158, n16157, n16156, 
        n16155, n16154, n16153, n16152, n16151, n16150, n16149, 
        n22322, n63, n28987, n66, n22321, n22320, n15751, n15750, 
        n15749, n15508, n15460, n6_adj_4771, n7_adj_4772, n8_adj_4773, 
        n9_adj_4774, n10_adj_4775, n11_adj_4776, n12_adj_4777, n13_adj_4778, 
        n14_adj_4779, n15_adj_4780, n16_adj_4781, n17_adj_4782, n18_adj_4783, 
        n19_adj_4784, n20_adj_4785, n21_adj_4786, n22_adj_4787, n23_adj_4788, 
        n24_adj_4789, n25_adj_4790, n15748, n15747, n15446, n15973, 
        n15972, n15971, n15970, n15969, n15968, n15967, n15966, 
        n15965, n15964, n15963, n15962, n15961, n15960, n15959, 
        n15958, n15957, n15956, n15955, n15954, n15953, n15952, 
        n15951, n15746, n15745, n15744, n15743, n15742, n15741, 
        n15740, n15739, n15738, n15737, n15736, n15735, n15734, 
        n15733, n15732, n15731, n15730, n15729, n15728, n15727, 
        n15726, n15725, n15724, n15723, n15950, n15949, n15948, 
        n15947, n63_adj_4791, n15946, n15945, n15944, n15943, n15942, 
        n15941, n15940, n15939, n15722, n15938, n15937, n15936, 
        n15935, n15721, n15934, n15720, n15933, n15932, n15931, 
        n15930, n15929, n15719, n15928, n15927, n15926, n15925, 
        n15924, n15923, n15922, n15921, n15920, n15919, n15918, 
        n15917, n15916, n15915, n15914, n15913, n15718, quadA_debounced, 
        quadB_debounced, n15717, n15912, n15716, n15715, n15911, 
        n15910, quadA_debounced_adj_4792, quadB_debounced_adj_4793, n22319, 
        n15909, n27464, n15908, n15907, n15906, n15905, n15904, 
        n15903, n15902, n15901, n15900, n15899, n15898, n15897, 
        n15896, n15895, n15894, n15893, n15892, n15891, n15890, 
        n15889, n15888, n15887, n15886, n15885, n15884, n4609, 
        n15883, n15882, n15881, n15880, n15879, n15878, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n4_adj_4794, n4677, n15877, n15876, n15875, n15874, n15873, 
        n15872, n15871, n3_adj_4795, n15870;
    wire [2:0]r_SM_Main_2__N_3426;
    
    wire n15869, n15868, n15867, n15866, n15865, n15864, n15863, 
        n15862, n15861, n15860, n15859, n15858, n15857, n15856, 
        n15855, n15854;
    wire [2:0]r_SM_Main_adj_4871;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_4873;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3497;
    
    wire n2, n15853, n15852, n15851, n15850, n15849, n15848, n15847, 
        n15846, n15845, n15844, n15843, n15842, n15841, n15840, 
        n15839, n15838, n15837, n15836, n15835, n15834;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15833, n15832;
    wire [1:0]reg_B_adj_4883;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15831, n15830, n4_adj_4802, n7_adj_4803, n8_adj_4804, n27374, 
        n27362, n27476, n15711, n15707, n15704, n15829, n15828, 
        n15827, n15826, n15825, n15824, n15823, n15822, n15821, 
        n15820, n15819, n15818, n15817, n15816, n15815, n15814, 
        n15813, n15812, n15811, n15810, n15809, n15808, n15807, 
        n15806, n15805, n15804, n15803, n15802, n15801, n15800, 
        n15799, n15798, n15797, n15796, n15795, n15701, n15700, 
        n15699, n15698, n15697, n15695, n15794, n15793, n15792, 
        n15791, n15790, n15789, n15788, n15787, n15694, n15692, 
        n15691, n15690, n15689, n15686, n15786, n15785, n15784, 
        n15783, n15782, n15781, n15780, n15779, n15778, n15777, 
        n15776, n15775, n15774, n15773, n15772, n15771, n15770, 
        n15769, n15768, n15767, n15766, n15765, n15764, n4_adj_4805, 
        n9520, n14254, n14253, n26557, n8595, n15685, n15684, 
        n1, n15683, n15682, n15681, n15680, n28904, n26153, n25291, 
        n1_adj_4806, n1_adj_4807, n1_adj_4808, n1_adj_4809, n1_adj_4810, 
        n1_adj_4811, n1_adj_4812, n1_adj_4813, n1_adj_4814, n1_adj_4815, 
        n1_adj_4816, n1_adj_4817, n1_adj_4818, n1_adj_4819, n1_adj_4820, 
        n1_adj_4821, n1_adj_4822, n1_adj_4823, n1_adj_4824, n1_adj_4825, 
        n1_adj_4826, n1_adj_4827, n1_adj_4828, n7_adj_4829, n28888, 
        n14264, n28359, n11648, n8439, n29784;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced, 
            quadB_debounced}), .n28904(n28904), .reg_B({reg_B}), .VCC_net(VCC_net), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n16183(n16183), .n15697(n15697), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(187[15] 192[4])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_40 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF h2_39 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.timer({timer}), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .GND_net(GND_net), .VCC_net(VCC_net), 
            .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), .start(start), 
            .n4(n4_adj_4802), .\state[0] (state[0]), .n66(n66), .LED_c(LED_c), 
            .\state[1] (state[1]), .n1929(n1929), .n19323(n19323), .neopxl_color({neopxl_color}), 
            .n16226(n16226), .n16225(n16225), .n16224(n16224), .n16223(n16223), 
            .n16222(n16222), .n16221(n16221), .n16220(n16220), .n16219(n16219), 
            .n16218(n16218), .n16217(n16217), .n16216(n16216), .n16215(n16215), 
            .n16214(n16214), .n16213(n16213), .n16212(n16212), .n16211(n16211), 
            .n16210(n16210), .n16209(n16209), .n16208(n16208), .n16207(n16207), 
            .n16206(n16206), .n16205(n16205), .n16204(n16204), .n16203(n16203), 
            .n16202(n16202), .n16201(n16201), .n16200(n16200), .n16199(n16199), 
            .n16198(n16198), .n16197(n16197), .n16196(n16196), .n25291(n25291), 
            .NEOPXL_c(NEOPXL_c), .n15701(n15701)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(44[10] 50[2])
    SB_CARRY add_541_8 (.CI(n22324), .I0(n30633), .I1(n19), .CO(n22325));
    SB_DFF dir_44 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n22545), .I0(encoder1_position[10]), 
            .I1(n15_adj_4780), .CO(n22546));
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4781), .I3(n22544), .O(displacement_23__N_26[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n22544), .I0(encoder1_position[9]), 
            .I1(n16_adj_4781), .CO(n22545));
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4782), .I3(n22543), .O(displacement_23__N_26[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n22543), .I0(encoder1_position[8]), 
            .I1(n17_adj_4782), .CO(n22544));
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4783), .I3(n22542), .O(displacement_23__N_26[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n22542), .I0(encoder1_position[7]), 
            .I1(n18_adj_4783), .CO(n22543));
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4784), .I3(n22541), .O(displacement_23__N_26[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n22541), .I0(encoder1_position[6]), 
            .I1(n19_adj_4784), .CO(n22542));
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4785), .I3(n22540), .O(displacement_23__N_26[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n22540), .I0(encoder1_position[5]), 
            .I1(n20_adj_4785), .CO(n22541));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4786), .I3(n22539), .O(displacement_23__N_26[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n22539), .I0(encoder1_position[4]), 
            .I1(n21_adj_4786), .CO(n22540));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4787), .I3(n22538), .O(displacement_23__N_26[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n22538), .I0(encoder1_position[3]), 
            .I1(n22_adj_4787), .CO(n22539));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4788), .I3(n22537), .O(displacement_23__N_26[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4767));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n22537), .I0(encoder1_position[2]), 
            .I1(n23_adj_4788), .CO(n22538));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4789), .I3(n22536), .O(displacement_23__N_26[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n22536), .I0(encoder1_position[1]), 
            .I1(n24_adj_4789), .CO(n22537));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4790), .I3(VCC_net), .O(displacement_23__N_26[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4790), .CO(n22536));
    SB_LUT4 i11167_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15742));   // verilog/coms.v(127[12] 300[6])
    defparam i11167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4787));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11168_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15743));   // verilog/coms.v(127[12] 300[6])
    defparam i11168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4766));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11169_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15744));   // verilog/coms.v(127[12] 300[6])
    defparam i11169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_13_lut (.I0(duty[11]), .I1(n30633), .I2(n14), .I3(n22329), 
            .O(pwm_setpoint_22__N_3[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_13 (.CI(n22329), .I0(n30633), .I1(n14), .CO(n22330));
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4765));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11170_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15745));   // verilog/coms.v(127[12] 300[6])
    defparam i11170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11171_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15746));   // verilog/coms.v(127[12] 300[6])
    defparam i11171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4764));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11166_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15741));   // verilog/coms.v(127[12] 300[6])
    defparam i11166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24034_2_lut (.I0(displacement[0]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29839));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24034_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_0_i1_3_lut (.I0(encoder0_position[0]), .I1(encoder1_position[0]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14154_4_lut (.I0(n1), .I1(n28359), .I2(n29839), .I3(control_mode[1]), 
            .O(motor_state[0]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14154_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i21516_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n14254), .I2(GND_net), 
            .I3(GND_net), .O(n27362));
    defparam i21516_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24129_2_lut (.I0(displacement[1]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29854));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24129_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_1_i1_3_lut (.I0(encoder0_position[1]), .I1(encoder1_position[1]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4806));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14400_4_lut (.I0(n1_adj_4806), .I1(n28359), .I2(n29854), 
            .I3(control_mode[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14400_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11172_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15747));   // verilog/coms.v(127[12] 300[6])
    defparam i11172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24253_2_lut (.I0(displacement[2]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29855));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24253_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_2_i1_3_lut (.I0(encoder0_position[2]), .I1(encoder1_position[2]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4807));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_2_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14401_4_lut (.I0(n1_adj_4807), .I1(n28359), .I2(n29855), 
            .I3(control_mode[1]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14401_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11173_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15748));   // verilog/coms.v(127[12] 300[6])
    defparam i11173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11174_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15749));   // verilog/coms.v(127[12] 300[6])
    defparam i11174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24254_2_lut (.I0(displacement[3]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29856));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24254_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24268_2_lut (.I0(displacement[17]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29870));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24268_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_3_i1_3_lut (.I0(encoder0_position[3]), .I1(encoder1_position[3]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4808));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_675_Mux_17_i1_3_lut (.I0(encoder0_position[17]), .I1(encoder1_position[17]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4822));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14416_4_lut (.I0(n1_adj_4822), .I1(n28359), .I2(n29870), 
            .I3(control_mode[1]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14416_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i14402_4_lut (.I0(n1_adj_4808), .I1(n28359), .I2(n29856), 
            .I3(control_mode[1]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14402_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24255_2_lut (.I0(displacement[4]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29857));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24255_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_4_i1_3_lut (.I0(encoder0_position[4]), .I1(encoder1_position[4]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4809));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_4_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14403_4_lut (.I0(n1_adj_4809), .I1(n28359), .I2(n29857), 
            .I3(control_mode[1]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14403_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24256_2_lut (.I0(displacement[5]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29858));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24256_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_5_i1_3_lut (.I0(encoder0_position[5]), .I1(encoder1_position[5]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4810));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_5_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_12_lut (.I0(duty[10]), .I1(n30633), .I2(n15), .I3(n22328), 
            .O(pwm_setpoint_22__N_3[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4785));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4784));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11175_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15750));   // verilog/coms.v(127[12] 300[6])
    defparam i11175_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_541_12 (.CI(n22328), .I0(n30633), .I1(n15), .CO(n22329));
    SB_LUT4 add_541_11_lut (.I0(duty[9]), .I1(n30633), .I2(n16), .I3(n22327), 
            .O(pwm_setpoint_22__N_3[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_9 (.CI(n22325), .I0(n30633), .I1(n18), .CO(n22326));
    SB_LUT4 add_541_7_lut (.I0(duty[5]), .I1(n30633), .I2(n20), .I3(n22323), 
            .O(pwm_setpoint_22__N_3[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_541_10_lut (.I0(duty[8]), .I1(n30633), .I2(n17), .I3(n22326), 
            .O(pwm_setpoint_22__N_3[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_10 (.CI(n22326), .I0(n30633), .I1(n17), .CO(n22327));
    SB_CARRY add_541_7 (.CI(n22323), .I0(n30633), .I1(n20), .CO(n22324));
    SB_LUT4 add_541_6_lut (.I0(duty[4]), .I1(n30633), .I2(n21), .I3(n22322), 
            .O(pwm_setpoint_22__N_3[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_6 (.CI(n22322), .I0(n30633), .I1(n21), .CO(n22323));
    SB_LUT4 add_541_5_lut (.I0(duty[3]), .I1(n30633), .I2(n22), .I3(n22321), 
            .O(pwm_setpoint_22__N_3[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_5 (.CI(n22321), .I0(n30633), .I1(n22), .CO(n22322));
    SB_LUT4 add_541_9_lut (.I0(duty[7]), .I1(n30633), .I2(n18), .I3(n22325), 
            .O(pwm_setpoint_22__N_3[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_541_4_lut (.I0(duty[2]), .I1(n30633), .I2(n23), .I3(n22320), 
            .O(pwm_setpoint_22__N_3[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_4 (.CI(n22320), .I0(n30633), .I1(n23), .CO(n22321));
    SB_LUT4 add_541_3_lut (.I0(duty[1]), .I1(n30633), .I2(n24), .I3(n22319), 
            .O(pwm_setpoint_22__N_3[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_3 (.CI(n22319), .I0(n30633), .I1(n24), .CO(n22320));
    SB_LUT4 add_541_2_lut (.I0(duty[0]), .I1(n30633), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_3[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_2 (.CI(VCC_net), .I0(n30633), .I1(n25), .CO(n22319));
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(144[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_541_8_lut (.I0(duty[6]), .I1(n30633), .I2(n19), .I3(n22324), 
            .O(pwm_setpoint_22__N_3[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_8_lut.LUT_INIT = 16'h8BB8;
    SB_DFF h1_38 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_IO SCL_pad (.PACKAGE_PIN(SCL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCL_pad.PIN_TYPE = 6'b011001;
    defparam SCL_pad.PULLUP = 1'b0;
    defparam SCL_pad.NEG_TRIGGER = 1'b0;
    defparam SCL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i24257_2_lut (.I0(displacement[6]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29859));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24257_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4783));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4782));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4781));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24269_2_lut (.I0(displacement[18]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29871));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24269_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_18_i1_3_lut (.I0(encoder0_position[18]), .I1(encoder1_position[18]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4823));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_18_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14417_4_lut (.I0(n1_adj_4823), .I1(n28359), .I2(n29871), 
            .I3(control_mode[1]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14417_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i4_4_lut (.I0(control_mode[5]), .I1(control_mode[7]), .I2(control_mode[4]), 
            .I3(control_mode[6]), .O(n10_adj_4770));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[3]), .I1(n10_adj_4770), .I2(control_mode[2]), 
            .I3(GND_net), .O(n28359));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24270_2_lut (.I0(displacement[19]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29872));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24270_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_19_i1_3_lut (.I0(encoder0_position[19]), .I1(encoder1_position[19]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4824));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_19_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14418_4_lut (.I0(n1_adj_4824), .I1(n28359), .I2(n29872), 
            .I3(control_mode[1]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14418_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4780));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_675_Mux_6_i1_3_lut (.I0(encoder0_position[6]), .I1(encoder1_position[6]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4811));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i14405_4_lut (.I0(n1_adj_4811), .I1(n28359), .I2(n29859), 
            .I3(control_mode[1]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14405_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4786));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[0]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14404_4_lut (.I0(n1_adj_4810), .I1(n28359), .I2(n29858), 
            .I3(control_mode[1]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14404_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11574_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4772), .I3(GND_net), .O(n16149));   // verilog/coms.v(127[12] 300[6])
    defparam i11574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11575_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4772), .I3(GND_net), .O(n16150));   // verilog/coms.v(127[12] 300[6])
    defparam i11575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11576_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4772), .I3(GND_net), .O(n16151));   // verilog/coms.v(127[12] 300[6])
    defparam i11576_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_26[23]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_LUT4 i11577_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4772), .I3(GND_net), .O(n16152));   // verilog/coms.v(127[12] 300[6])
    defparam i11577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11578_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4772), .I3(GND_net), .O(n16153));   // verilog/coms.v(127[12] 300[6])
    defparam i11578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24258_2_lut (.I0(displacement[7]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29860));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24258_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_7_i1_3_lut (.I0(encoder0_position[7]), .I1(encoder1_position[7]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4812));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_7_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11579_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4772), .I3(GND_net), .O(n16154));   // verilog/coms.v(127[12] 300[6])
    defparam i11579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11580_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4772), .I3(GND_net), .O(n16155));   // verilog/coms.v(127[12] 300[6])
    defparam i11580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14406_4_lut (.I0(n1_adj_4812), .I1(n28359), .I2(n29860), 
            .I3(control_mode[1]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14406_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11581_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n4772), .I3(GND_net), .O(n16156));   // verilog/coms.v(127[12] 300[6])
    defparam i11581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11582_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n4772), .I3(GND_net), .O(n16157));   // verilog/coms.v(127[12] 300[6])
    defparam i11582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11583_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n4772), .I3(GND_net), .O(n16158));   // verilog/coms.v(127[12] 300[6])
    defparam i11583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11584_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n4772), .I3(GND_net), .O(n16159));   // verilog/coms.v(127[12] 300[6])
    defparam i11584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11585_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n4772), .I3(GND_net), .O(n16160));   // verilog/coms.v(127[12] 300[6])
    defparam i11585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11586_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n4772), .I3(GND_net), .O(n16161));   // verilog/coms.v(127[12] 300[6])
    defparam i11586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11176_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15751));   // verilog/coms.v(127[12] 300[6])
    defparam i11176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11177_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15752));   // verilog/coms.v(127[12] 300[6])
    defparam i11177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11587_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n4772), .I3(GND_net), .O(n16162));   // verilog/coms.v(127[12] 300[6])
    defparam i11587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11588_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n4772), .I3(GND_net), .O(n16163));   // verilog/coms.v(127[12] 300[6])
    defparam i11588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11589_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n4772), .I3(GND_net), .O(n16164));   // verilog/coms.v(127[12] 300[6])
    defparam i11589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_24_lut (.I0(duty[22]), .I1(n30633), .I2(n3), .I3(n22340), 
            .O(pwm_setpoint_22__N_3[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11178_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15753));   // verilog/coms.v(127[12] 300[6])
    defparam i11178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11182_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15757));   // verilog/coms.v(127[12] 300[6])
    defparam i11182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11179_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15754));   // verilog/coms.v(127[12] 300[6])
    defparam i11179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11183_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15758));   // verilog/coms.v(127[12] 300[6])
    defparam i11183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11590_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n4772), .I3(GND_net), .O(n16165));   // verilog/coms.v(127[12] 300[6])
    defparam i11590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11591_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n4772), .I3(GND_net), .O(n16166));   // verilog/coms.v(127[12] 300[6])
    defparam i11591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11592_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n4772), .I3(GND_net), .O(n16167));   // verilog/coms.v(127[12] 300[6])
    defparam i11592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11593_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n4772), .I3(GND_net), .O(n16168));   // verilog/coms.v(127[12] 300[6])
    defparam i11593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11594_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n4772), .I3(GND_net), .O(n16169));   // verilog/coms.v(127[12] 300[6])
    defparam i11594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11595_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n4772), .I3(GND_net), .O(n16170));   // verilog/coms.v(127[12] 300[6])
    defparam i11595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11596_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n4772), .I3(GND_net), .O(n16171));   // verilog/coms.v(127[12] 300[6])
    defparam i11596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11597_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n4772), .I3(GND_net), .O(n16172));   // verilog/coms.v(127[12] 300[6])
    defparam i11597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11598_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n4772), .I3(GND_net), .O(n16173));   // verilog/coms.v(127[12] 300[6])
    defparam i11598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11599_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n4772), .I3(GND_net), .O(n16174));   // verilog/coms.v(127[12] 300[6])
    defparam i11599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11184_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15759));   // verilog/coms.v(127[12] 300[6])
    defparam i11184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_23_lut (.I0(duty[21]), .I1(n30633), .I2(n4_adj_4764), 
            .I3(n22339), .O(pwm_setpoint_22__N_3[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i24259_2_lut (.I0(displacement[8]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29861));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24259_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_8_i1_3_lut (.I0(encoder0_position[8]), .I1(encoder1_position[8]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4813));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_8_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11600_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n4772), .I3(GND_net), .O(n16175));   // verilog/coms.v(127[12] 300[6])
    defparam i11600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11601_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n4772), .I3(GND_net), .O(n16176));   // verilog/coms.v(127[12] 300[6])
    defparam i11601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11602_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n4772), .I3(GND_net), .O(n16177));   // verilog/coms.v(127[12] 300[6])
    defparam i11602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11603_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n4772), .I3(GND_net), .O(n16178));   // verilog/coms.v(127[12] 300[6])
    defparam i11603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14407_4_lut (.I0(n1_adj_4813), .I1(n28359), .I2(n29861), 
            .I3(control_mode[1]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14407_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i24260_2_lut (.I0(displacement[9]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29862));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24260_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_9_i1_3_lut (.I0(encoder0_position[9]), .I1(encoder1_position[9]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4814));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_9_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14408_4_lut (.I0(n1_adj_4814), .I1(n28359), .I2(n29862), 
            .I3(control_mode[1]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14408_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4790));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24267_2_lut (.I0(displacement[16]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29869));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24267_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_675_Mux_16_i1_3_lut (.I0(encoder0_position[16]), .I1(encoder1_position[16]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4821));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_16_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14415_4_lut (.I0(n1_adj_4821), .I1(n28359), .I2(n29869), 
            .I3(control_mode[1]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14415_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11180_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15755));   // verilog/coms.v(127[12] 300[6])
    defparam i11180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n26561), .I1(n2649), .I2(n14291), .I3(n4452), 
            .O(n26611));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_3_lut (.I0(n123), .I1(n26611), .I2(n63), .I3(GND_net), 
            .O(n7_adj_4829));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut.LUT_INIT = 16'h8c8c;
    SB_LUT4 i2_4_lut (.I0(n7_adj_4829), .I1(n123), .I2(n14253), .I3(n8595), 
            .O(n6));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'haeaf;
    SB_LUT4 i3_4_lut (.I0(n63_adj_4791), .I1(n6), .I2(n14288), .I3(\FRAME_MATCHER.state_31__N_2672 [1]), 
            .O(n31239));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hdfdd;
    SB_LUT4 i2_4_lut_adj_1635 (.I0(n122), .I1(\FRAME_MATCHER.state_31__N_2672 [2]), 
            .I2(n5_adj_4769), .I3(n14288), .O(n7));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1635.LUT_INIT = 16'ha0ec;
    SB_LUT4 i4_4_lut_adj_1636 (.I0(n7), .I1(n8_adj_4804), .I2(n63_adj_4791), 
            .I3(n7_adj_4803), .O(n31238));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1636.LUT_INIT = 16'hffef;
    SB_CARRY add_541_23 (.CI(n22339), .I0(n30633), .I1(n4_adj_4764), .CO(n22340));
    SB_LUT4 i11181_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15756));   // verilog/coms.v(127[12] 300[6])
    defparam i11181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24213_4_lut (.I0(state[0]), .I1(start), .I2(n19323), .I3(\neo_pixel_transmitter.done ), 
            .O(n29784));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24213_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 i18_4_lut (.I0(n4_adj_4802), .I1(n29784), .I2(state[1]), .I3(n66), 
            .O(n25291));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i11608_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n28904), 
            .I3(GND_net), .O(n16183));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11608_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11610_3_lut (.I0(quadA_debounced_adj_4792), .I1(reg_B_adj_4883[1]), 
            .I2(n28888), .I3(GND_net), .O(n16185));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11610_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut (.I0(n4677), .I1(DE_c), .I2(n14279), .I3(n4609), 
            .O(n25997));   // verilog/coms.v(127[12] 300[6])
    defparam i12_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i11132_3_lut (.I0(n15619), .I1(r_Bit_Index[0]), .I2(n15508), 
            .I3(GND_net), .O(n15707));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11132_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i11614_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n15460), .I3(GND_net), .O(n16189));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11615_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n15460), .I3(GND_net), .O(n16190));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11616_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n15460), .I3(GND_net), .O(n16191));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11617_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n15460), .I3(GND_net), .O(n16192));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11618_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n15460), .I3(GND_net), .O(n16193));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11619_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n15460), .I3(GND_net), .O(n16194));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11620_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n15460), .I3(GND_net), .O(n16195));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11621_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n1929), .I3(GND_net), .O(n16196));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11621_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_26[22]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_26[21]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_26[20]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_26[19]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_26[18]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_26[17]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_26[16]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_26[15]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_26[14]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_26[13]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_26[12]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_26[11]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_26[10]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_26[9]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_26[8]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_26[7]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_26[6]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_26[5]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_26[4]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_26[3]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_26[2]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_26[1]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[22]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[21]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[20]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[19]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[18]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[17]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[16]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[15]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[14]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[13]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[12]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[11]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[10]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[9]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[8]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[7]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[6]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[5]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[4]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[3]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[2]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[1]));   // verilog/TinyFPGA_B.v(98[10] 111[6])
    SB_LUT4 i11622_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n1929), .I3(GND_net), .O(n16197));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11623_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n1929), .I3(GND_net), .O(n16198));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11624_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n1929), .I3(GND_net), .O(n16199));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11625_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n1929), .I3(GND_net), .O(n16200));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4789));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11626_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n1929), .I3(GND_net), .O(n16201));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11627_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n1929), .I3(GND_net), .O(n16202));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11628_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n1929), .I3(GND_net), .O(n16203));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11629_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n1929), .I3(GND_net), .O(n16204));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11630_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n1929), .I3(GND_net), .O(n16205));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11631_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n1929), .I3(GND_net), .O(n16206));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11632_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n1929), .I3(GND_net), .O(n16207));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11633_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n1929), .I3(GND_net), .O(n16208));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11634_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n1929), .I3(GND_net), .O(n16209));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11635_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n1929), .I3(GND_net), .O(n16210));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11636_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n1929), .I3(GND_net), .O(n16211));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11637_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n1929), .I3(GND_net), .O(n16212));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11638_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n1929), .I3(GND_net), .O(n16213));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11639_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n1929), .I3(GND_net), .O(n16214));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11640_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n1929), .I3(GND_net), .O(n16215));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_22_lut (.I0(duty[20]), .I1(n30633), .I2(n5_adj_4765), 
            .I3(n22338), .O(pwm_setpoint_22__N_3[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_22 (.CI(n22338), .I0(n30633), .I1(n5_adj_4765), .CO(n22339));
    SB_LUT4 i11641_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n1929), .I3(GND_net), .O(n16216));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11642_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n1929), .I3(GND_net), .O(n16217));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11643_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n1929), .I3(GND_net), .O(n16218));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11644_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n1929), .I3(GND_net), .O(n16219));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11645_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n1929), .I3(GND_net), .O(n16220));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11646_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n1929), .I3(GND_net), .O(n16221));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_21_lut (.I0(duty[19]), .I1(n30633), .I2(n6_adj_4766), 
            .I3(n22337), .O(pwm_setpoint_22__N_3[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_541_21 (.CI(n22337), .I0(n30633), .I1(n6_adj_4766), .CO(n22338));
    SB_LUT4 i11647_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n1929), .I3(GND_net), .O(n16222));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11648_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n1929), .I3(GND_net), .O(n16223));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11648_3_lut.LUT_INIT = 16'hcaca;
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i11649_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n1929), .I3(GND_net), .O(n16224));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11650_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n1929), .I3(GND_net), .O(n16225));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11651_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n1929), .I3(GND_net), .O(n16226));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11652_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n18753), 
            .I3(n14264), .O(n16227));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11652_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11129_3_lut (.I0(n27476), .I1(r_Bit_Index_adj_4873[0]), .I2(n27464), 
            .I3(GND_net), .O(n15704));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11129_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 add_541_20_lut (.I0(duty[18]), .I1(n30633), .I2(n7_adj_4767), 
            .I3(n22336), .O(pwm_setpoint_22__N_3[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24261_2_lut (.I0(displacement[10]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29863));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24261_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_10_i1_3_lut (.I0(encoder0_position[10]), .I1(encoder1_position[10]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4815));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_10_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14409_4_lut (.I0(n1_adj_4815), .I1(n28359), .I2(n29863), 
            .I3(control_mode[1]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14409_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11136_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4768), 
            .I3(n14259), .O(n15711));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11136_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11140_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n4772), .I3(GND_net), .O(n15715));   // verilog/coms.v(127[12] 300[6])
    defparam i11140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11141_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n4772), .I3(GND_net), .O(n15716));   // verilog/coms.v(127[12] 300[6])
    defparam i11141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11142_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n4772), .I3(GND_net), .O(n15717));   // verilog/coms.v(127[12] 300[6])
    defparam i11142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11143_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n4772), .I3(GND_net), .O(n15718));   // verilog/coms.v(127[12] 300[6])
    defparam i11143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11144_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n4772), .I3(GND_net), .O(n15719));   // verilog/coms.v(127[12] 300[6])
    defparam i11144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11145_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n4772), .I3(GND_net), .O(n15720));   // verilog/coms.v(127[12] 300[6])
    defparam i11145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11146_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n4772), .I3(GND_net), .O(n15721));   // verilog/coms.v(127[12] 300[6])
    defparam i11146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11147_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n4772), .I3(GND_net), .O(n15722));   // verilog/coms.v(127[12] 300[6])
    defparam i11147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11148_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n4772), .I3(GND_net), .O(n15723));   // verilog/coms.v(127[12] 300[6])
    defparam i11148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11149_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n4772), .I3(GND_net), .O(n15724));   // verilog/coms.v(127[12] 300[6])
    defparam i11149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11150_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n4772), .I3(GND_net), .O(n15725));   // verilog/coms.v(127[12] 300[6])
    defparam i11150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24262_2_lut (.I0(displacement[11]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29864));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24262_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_11_i1_3_lut (.I0(encoder0_position[11]), .I1(encoder1_position[11]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4816));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_11_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14410_4_lut (.I0(n1_adj_4816), .I1(n28359), .I2(n29864), 
            .I3(control_mode[1]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14410_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11151_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n4772), .I3(GND_net), .O(n15726));   // verilog/coms.v(127[12] 300[6])
    defparam i11151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11152_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n4772), .I3(GND_net), .O(n15727));   // verilog/coms.v(127[12] 300[6])
    defparam i11152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11153_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n4772), .I3(GND_net), .O(n15728));   // verilog/coms.v(127[12] 300[6])
    defparam i11153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11154_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n4772), .I3(GND_net), .O(n15729));   // verilog/coms.v(127[12] 300[6])
    defparam i11154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11155_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n4772), .I3(GND_net), .O(n15730));   // verilog/coms.v(127[12] 300[6])
    defparam i11155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11156_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n4772), .I3(GND_net), .O(n15731));   // verilog/coms.v(127[12] 300[6])
    defparam i11156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11157_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n4772), .I3(GND_net), .O(n15732));   // verilog/coms.v(127[12] 300[6])
    defparam i11157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11158_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n4772), .I3(GND_net), .O(n15733));   // verilog/coms.v(127[12] 300[6])
    defparam i11158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24263_2_lut (.I0(displacement[12]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29865));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24263_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11159_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n4772), .I3(GND_net), .O(n15734));   // verilog/coms.v(127[12] 300[6])
    defparam i11159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11160_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n4772), .I3(GND_net), .O(n15735));   // verilog/coms.v(127[12] 300[6])
    defparam i11160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_675_Mux_12_i1_3_lut (.I0(encoder0_position[12]), .I1(encoder1_position[12]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4817));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11161_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n4772), .I3(GND_net), .O(n15736));   // verilog/coms.v(127[12] 300[6])
    defparam i11161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14411_4_lut (.I0(n1_adj_4817), .I1(n28359), .I2(n29865), 
            .I3(control_mode[1]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14411_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11162_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n4772), .I3(GND_net), .O(n15737));   // verilog/coms.v(127[12] 300[6])
    defparam i11162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11163_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15738));   // verilog/coms.v(127[12] 300[6])
    defparam i11163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24264_2_lut (.I0(displacement[13]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29866));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24264_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_13_i1_3_lut (.I0(encoder0_position[13]), .I1(encoder1_position[13]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4818));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_13_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14412_4_lut (.I0(n1_adj_4818), .I1(n28359), .I2(n29866), 
            .I3(control_mode[1]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14412_4_lut.LUT_INIT = 16'h3022;
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i24265_2_lut (.I0(displacement[14]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29867));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24265_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_14_i1_3_lut (.I0(encoder0_position[14]), .I1(encoder1_position[14]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4819));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14413_4_lut (.I0(n1_adj_4819), .I1(n28359), .I2(n29867), 
            .I3(control_mode[1]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14413_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11164_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15739));   // verilog/coms.v(127[12] 300[6])
    defparam i11164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24266_2_lut (.I0(displacement[15]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29868));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24266_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_15_i1_3_lut (.I0(encoder0_position[15]), .I1(encoder1_position[15]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4820));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14414_4_lut (.I0(n1_adj_4820), .I1(n28359), .I2(n29868), 
            .I3(control_mode[1]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14414_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11185_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15760));   // verilog/coms.v(127[12] 300[6])
    defparam i11185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4788));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11188_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15763));   // verilog/coms.v(127[12] 300[6])
    defparam i11188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4773));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11189_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15764));   // verilog/coms.v(127[12] 300[6])
    defparam i11189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11190_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15765));   // verilog/coms.v(127[12] 300[6])
    defparam i11190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11165_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15740));   // verilog/coms.v(127[12] 300[6])
    defparam i11165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11191_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15766));   // verilog/coms.v(127[12] 300[6])
    defparam i11191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11192_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15767));   // verilog/coms.v(127[12] 300[6])
    defparam i11192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11193_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15768));   // verilog/coms.v(127[12] 300[6])
    defparam i11193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11194_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n27965), 
            .I3(GND_net), .O(n15769));   // verilog/coms.v(127[12] 300[6])
    defparam i11194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11195_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n27965), 
            .I3(GND_net), .O(n15770));   // verilog/coms.v(127[12] 300[6])
    defparam i11195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11196_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n27965), 
            .I3(GND_net), .O(n15771));   // verilog/coms.v(127[12] 300[6])
    defparam i11196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11197_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n27965), 
            .I3(GND_net), .O(n15772));   // verilog/coms.v(127[12] 300[6])
    defparam i11197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4779));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24271_2_lut (.I0(displacement[20]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29873));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24271_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_20_i1_3_lut (.I0(encoder0_position[20]), .I1(encoder1_position[20]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4825));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_20_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14419_4_lut (.I0(n1_adj_4825), .I1(n28359), .I2(n29873), 
            .I3(control_mode[1]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14419_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11198_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n27965), 
            .I3(GND_net), .O(n15773));   // verilog/coms.v(127[12] 300[6])
    defparam i11198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11199_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n27965), 
            .I3(GND_net), .O(n15774));   // verilog/coms.v(127[12] 300[6])
    defparam i11199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11200_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n27965), 
            .I3(GND_net), .O(n15775));   // verilog/coms.v(127[12] 300[6])
    defparam i11200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11201_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n27965), 
            .I3(GND_net), .O(n15776));   // verilog/coms.v(127[12] 300[6])
    defparam i11201_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24272_2_lut (.I0(displacement[21]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29874));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24272_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_21_i1_3_lut (.I0(encoder0_position[21]), .I1(encoder1_position[21]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4826));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14420_4_lut (.I0(n1_adj_4826), .I1(n28359), .I2(n29874), 
            .I3(control_mode[1]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14420_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11202_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n27965), 
            .I3(GND_net), .O(n15777));   // verilog/coms.v(127[12] 300[6])
    defparam i11202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11186_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15761));   // verilog/coms.v(127[12] 300[6])
    defparam i11186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4778));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11203_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n27965), 
            .I3(GND_net), .O(n15778));   // verilog/coms.v(127[12] 300[6])
    defparam i11203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11204_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n27965), 
            .I3(GND_net), .O(n15779));   // verilog/coms.v(127[12] 300[6])
    defparam i11204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11205_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n27965), 
            .I3(GND_net), .O(n15780));   // verilog/coms.v(127[12] 300[6])
    defparam i11205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11206_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n27965), 
            .I3(GND_net), .O(n15781));   // verilog/coms.v(127[12] 300[6])
    defparam i11206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11207_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n27965), 
            .I3(GND_net), .O(n15782));   // verilog/coms.v(127[12] 300[6])
    defparam i11207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4777));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11208_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n27965), 
            .I3(GND_net), .O(n15783));   // verilog/coms.v(127[12] 300[6])
    defparam i11208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11209_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n27965), 
            .I3(GND_net), .O(n15784));   // verilog/coms.v(127[12] 300[6])
    defparam i11209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4772));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11210_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n27965), 
            .I3(GND_net), .O(n15785));   // verilog/coms.v(127[12] 300[6])
    defparam i11210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11211_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n27965), 
            .I3(GND_net), .O(n15786));   // verilog/coms.v(127[12] 300[6])
    defparam i11211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11212_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n27965), 
            .I3(GND_net), .O(n15787));   // verilog/coms.v(127[12] 300[6])
    defparam i11212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4776));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11213_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n27965), 
            .I3(GND_net), .O(n15788));   // verilog/coms.v(127[12] 300[6])
    defparam i11213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11214_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n27965), 
            .I3(GND_net), .O(n15789));   // verilog/coms.v(127[12] 300[6])
    defparam i11214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4775));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11215_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n27965), 
            .I3(GND_net), .O(n15790));   // verilog/coms.v(127[12] 300[6])
    defparam i11215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11216_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n27965), 
            .I3(GND_net), .O(n15791));   // verilog/coms.v(127[12] 300[6])
    defparam i11216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11217_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n27965), 
            .I3(GND_net), .O(n15792));   // verilog/coms.v(127[12] 300[6])
    defparam i11217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11218_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n27965), 
            .I3(GND_net), .O(n15793));   // verilog/coms.v(127[12] 300[6])
    defparam i11218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4771));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11219_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n27965), 
            .I3(GND_net), .O(n15794));   // verilog/coms.v(127[12] 300[6])
    defparam i11219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11220_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n27965), 
            .I3(GND_net), .O(n15795));   // verilog/coms.v(127[12] 300[6])
    defparam i11220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11221_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n27965), 
            .I3(GND_net), .O(n15796));   // verilog/coms.v(127[12] 300[6])
    defparam i11221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11222_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n27965), 
            .I3(GND_net), .O(n15797));   // verilog/coms.v(127[12] 300[6])
    defparam i11222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11223_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n27965), 
            .I3(GND_net), .O(n15798));   // verilog/coms.v(127[12] 300[6])
    defparam i11223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11224_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n11648), .I3(GND_net), .O(n15799));   // verilog/coms.v(127[12] 300[6])
    defparam i11224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11225_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n11648), .I3(GND_net), .O(n15800));   // verilog/coms.v(127[12] 300[6])
    defparam i11225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11226_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n11648), .I3(GND_net), .O(n15801));   // verilog/coms.v(127[12] 300[6])
    defparam i11226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11227_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n11648), .I3(GND_net), .O(n15802));   // verilog/coms.v(127[12] 300[6])
    defparam i11227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11228_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n11648), .I3(GND_net), .O(n15803));   // verilog/coms.v(127[12] 300[6])
    defparam i11228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11229_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n11648), .I3(GND_net), .O(n15804));   // verilog/coms.v(127[12] 300[6])
    defparam i11229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11230_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n11648), .I3(GND_net), .O(n15805));   // verilog/coms.v(127[12] 300[6])
    defparam i11230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24273_2_lut (.I0(displacement[22]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29875));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24273_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_675_Mux_22_i1_3_lut (.I0(encoder0_position[22]), .I1(encoder1_position[22]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4827));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14421_4_lut (.I0(n1_adj_4827), .I1(n28359), .I2(n29875), 
            .I3(control_mode[1]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14421_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i11231_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n11648), .I3(GND_net), .O(n15806));   // verilog/coms.v(127[12] 300[6])
    defparam i11231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11232_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n11648), .I3(GND_net), .O(n15807));   // verilog/coms.v(127[12] 300[6])
    defparam i11232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11233_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n11648), .I3(GND_net), .O(n15808));   // verilog/coms.v(127[12] 300[6])
    defparam i11233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4774));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11234_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n11648), .I3(GND_net), .O(n15809));   // verilog/coms.v(127[12] 300[6])
    defparam i11234_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_541_20 (.CI(n22336), .I0(n30633), .I1(n7_adj_4767), .CO(n22337));
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n2), .I3(n22558), .O(displacement_23__N_26[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_541_19_lut (.I0(duty[17]), .I1(n30633), .I2(n8), .I3(n22335), 
            .O(pwm_setpoint_22__N_3[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11235_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n11648), .I3(GND_net), .O(n15810));   // verilog/coms.v(127[12] 300[6])
    defparam i11235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4795), .I3(n22557), .O(displacement_23__N_26[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_541_19 (.CI(n22335), .I0(n30633), .I1(n8), .CO(n22336));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4794));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n22557), .I0(encoder1_position[22]), 
            .I1(n3_adj_4795), .CO(n22558));
    SB_LUT4 i11236_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n11648), .I3(GND_net), .O(n15811));   // verilog/coms.v(127[12] 300[6])
    defparam i11236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11237_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n11648), .I3(GND_net), .O(n15812));   // verilog/coms.v(127[12] 300[6])
    defparam i11237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11238_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n11648), .I3(GND_net), .O(n15813));   // verilog/coms.v(127[12] 300[6])
    defparam i11238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11239_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n11648), .I3(GND_net), .O(n15814));   // verilog/coms.v(127[12] 300[6])
    defparam i11239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11240_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n11648), .I3(GND_net), .O(n15815));   // verilog/coms.v(127[12] 300[6])
    defparam i11240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11241_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n11648), .I3(GND_net), .O(n15816));   // verilog/coms.v(127[12] 300[6])
    defparam i11241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24274_2_lut (.I0(displacement[23]), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n29876));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i24274_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n4_adj_4794), .I3(n22556), .O(displacement_23__N_26[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_675_Mux_23_i1_3_lut (.I0(encoder0_position[23]), .I1(encoder1_position[23]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n1_adj_4828));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam mux_675_Mux_23_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14422_4_lut (.I0(n1_adj_4828), .I1(n28359), .I2(n29876), 
            .I3(control_mode[1]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(166[5] 170[10])
    defparam i14422_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4795));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3426[2]), 
            .I3(r_SM_Main[0]), .O(n15446));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(203[21:58])
    defparam encoder1_position_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n15446), 
            .I3(rx_data_ready), .O(n26153));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i24759_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n26557));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i24759_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n22556), .I0(encoder1_position[21]), 
            .I1(n4_adj_4794), .CO(n22557));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5), .I3(n22555), .O(displacement_23__N_26[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(108[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n22555), .I0(encoder1_position[20]), 
            .I1(n5), .CO(n22556));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4771), .I3(n22554), .O(displacement_23__N_26[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n22554), .I0(encoder1_position[19]), 
            .I1(n6_adj_4771), .CO(n22555));
    SB_LUT4 add_541_18_lut (.I0(duty[16]), .I1(n30633), .I2(n9), .I3(n22334), 
            .O(pwm_setpoint_22__N_3[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11242_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n11648), .I3(GND_net), .O(n15817));   // verilog/coms.v(127[12] 300[6])
    defparam i11242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11243_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n11648), .I3(GND_net), .O(n15818));   // verilog/coms.v(127[12] 300[6])
    defparam i11243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4772), .I3(n22553), .O(displacement_23__N_26[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n22553), .I0(encoder1_position[18]), 
            .I1(n7_adj_4772), .CO(n22554));
    SB_LUT4 i11244_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n11648), .I3(GND_net), .O(n15819));   // verilog/coms.v(127[12] 300[6])
    defparam i11244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11245_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n11648), .I3(GND_net), .O(n15820));   // verilog/coms.v(127[12] 300[6])
    defparam i11245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11246_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n11648), .I3(GND_net), .O(n15821));   // verilog/coms.v(127[12] 300[6])
    defparam i11246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11247_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n11648), .I3(GND_net), .O(n15822));   // verilog/coms.v(127[12] 300[6])
    defparam i11247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11248_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n11648), .I3(GND_net), .O(n15823));   // verilog/coms.v(127[12] 300[6])
    defparam i11248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11249_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n11648), .I3(GND_net), .O(n15824));   // verilog/coms.v(127[12] 300[6])
    defparam i11249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11250_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n11648), .I3(GND_net), .O(n15825));   // verilog/coms.v(127[12] 300[6])
    defparam i11250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11251_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n11648), .I3(GND_net), .O(n15826));   // verilog/coms.v(127[12] 300[6])
    defparam i11251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11252_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n11648), .I3(GND_net), .O(n15827));   // verilog/coms.v(127[12] 300[6])
    defparam i11252_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_541_11 (.CI(n22327), .I0(n30633), .I1(n16), .CO(n22328));
    SB_LUT4 i11253_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n11648), .I3(GND_net), .O(n15828));   // verilog/coms.v(127[12] 300[6])
    defparam i11253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11254_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n11648), .I3(GND_net), .O(n15829));   // verilog/coms.v(127[12] 300[6])
    defparam i11254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11255_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n11648), .I3(GND_net), .O(n15830));   // verilog/coms.v(127[12] 300[6])
    defparam i11255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11256_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n11648), .I3(GND_net), .O(n15831));   // verilog/coms.v(127[12] 300[6])
    defparam i11256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4773), .I3(n22552), .O(displacement_23__N_26[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11257_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n11648), .I3(GND_net), .O(n15832));   // verilog/coms.v(127[12] 300[6])
    defparam i11257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11258_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n11648), .I3(GND_net), .O(n15833));   // verilog/coms.v(127[12] 300[6])
    defparam i11258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11259_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n11648), .I3(GND_net), .O(n15834));   // verilog/coms.v(127[12] 300[6])
    defparam i11259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11260_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n11648), .I3(GND_net), .O(n15835));   // verilog/coms.v(127[12] 300[6])
    defparam i11260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11261_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n11648), .I3(GND_net), .O(n15836));   // verilog/coms.v(127[12] 300[6])
    defparam i11261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11262_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n11648), .I3(GND_net), .O(n15837));   // verilog/coms.v(127[12] 300[6])
    defparam i11262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11263_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n11648), .I3(GND_net), .O(n15838));   // verilog/coms.v(127[12] 300[6])
    defparam i11263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11264_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n11648), .I3(GND_net), .O(n15839));   // verilog/coms.v(127[12] 300[6])
    defparam i11264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11265_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n11648), .I3(GND_net), .O(n15840));   // verilog/coms.v(127[12] 300[6])
    defparam i11265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11105_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n18753), 
            .I3(n14259), .O(n15680));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11105_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i11106_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n14264), 
            .O(n15681));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11106_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11107_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n4772), .I3(GND_net), .O(n15682));   // verilog/coms.v(127[12] 300[6])
    defparam i11107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11108_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n14259), 
            .O(n15683));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11108_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11109_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4763), 
            .I3(n14264), .O(n15684));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11109_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11110_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4763), 
            .I3(n14259), .O(n15685));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11110_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_541_18 (.CI(n22334), .I0(n30633), .I1(n9), .CO(n22335));
    SB_LUT4 i11111_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4768), 
            .I3(n14264), .O(n15686));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11111_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11266_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n11648), .I3(GND_net), .O(n15841));   // verilog/coms.v(127[12] 300[6])
    defparam i11266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11267_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n11648), .I3(GND_net), .O(n15842));   // verilog/coms.v(127[12] 300[6])
    defparam i11267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11268_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n11648), .I3(GND_net), .O(n15843));   // verilog/coms.v(127[12] 300[6])
    defparam i11268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11269_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n11648), .I3(GND_net), .O(n15844));   // verilog/coms.v(127[12] 300[6])
    defparam i11269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11270_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n11648), .I3(GND_net), .O(n15845));   // verilog/coms.v(127[12] 300[6])
    defparam i11270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11271_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n11648), .I3(GND_net), .O(n15846));   // verilog/coms.v(127[12] 300[6])
    defparam i11271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11272_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n11648), .I3(GND_net), .O(n15847));   // verilog/coms.v(127[12] 300[6])
    defparam i11272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11114_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15689));   // verilog/coms.v(127[12] 300[6])
    defparam i11114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11115_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n27965), 
            .I3(GND_net), .O(n15690));   // verilog/coms.v(127[12] 300[6])
    defparam i11115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11116_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n27965), 
            .I3(GND_net), .O(n15691));   // verilog/coms.v(127[12] 300[6])
    defparam i11116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11117_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n4774), .I3(GND_net), .O(n15692));   // verilog/coms.v(127[12] 300[6])
    defparam i11117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11119_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4772), .I3(GND_net), .O(n15694));   // verilog/coms.v(127[12] 300[6])
    defparam i11119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11273_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n11648), .I3(GND_net), .O(n15848));   // verilog/coms.v(127[12] 300[6])
    defparam i11273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11274_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n11648), .I3(GND_net), .O(n15849));   // verilog/coms.v(127[12] 300[6])
    defparam i11274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11275_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n11648), .I3(GND_net), .O(n15850));   // verilog/coms.v(127[12] 300[6])
    defparam i11275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11276_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n11648), .I3(GND_net), .O(n15851));   // verilog/coms.v(127[12] 300[6])
    defparam i11276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11277_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n11648), .I3(GND_net), .O(n15852));   // verilog/coms.v(127[12] 300[6])
    defparam i11277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n14254), .I3(n4609), .O(n63_adj_4791));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i11278_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n11648), .I3(GND_net), .O(n15853));   // verilog/coms.v(127[12] 300[6])
    defparam i11278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11279_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n11648), .I3(GND_net), .O(n15854));   // verilog/coms.v(127[12] 300[6])
    defparam i11279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11280_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n11648), .I3(GND_net), .O(n15855));   // verilog/coms.v(127[12] 300[6])
    defparam i11280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11281_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n11648), .I3(GND_net), .O(n15856));   // verilog/coms.v(127[12] 300[6])
    defparam i11281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11282_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n11648), .I3(GND_net), .O(n15857));   // verilog/coms.v(127[12] 300[6])
    defparam i11282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11283_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n11648), .I3(GND_net), .O(n15858));   // verilog/coms.v(127[12] 300[6])
    defparam i11283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11284_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n11648), .I3(GND_net), .O(n15859));   // verilog/coms.v(127[12] 300[6])
    defparam i11284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11285_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n11648), .I3(GND_net), .O(n15860));   // verilog/coms.v(127[12] 300[6])
    defparam i11285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11286_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n11648), .I3(GND_net), .O(n15861));   // verilog/coms.v(127[12] 300[6])
    defparam i11286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11287_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n11648), .I3(GND_net), .O(n15862));   // verilog/coms.v(127[12] 300[6])
    defparam i11287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11288_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n11648), .I3(GND_net), .O(n15863));   // verilog/coms.v(127[12] 300[6])
    defparam i11288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11289_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n11648), .I3(GND_net), .O(n15864));   // verilog/coms.v(127[12] 300[6])
    defparam i11289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_17_lut (.I0(duty[15]), .I1(n30633), .I2(n10), .I3(n22333), 
            .O(pwm_setpoint_22__N_3[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11290_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n11648), .I3(GND_net), .O(n15865));   // verilog/coms.v(127[12] 300[6])
    defparam i11290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11291_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n11648), .I3(GND_net), .O(n15866));   // verilog/coms.v(127[12] 300[6])
    defparam i11291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11292_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n11648), .I3(GND_net), .O(n15867));   // verilog/coms.v(127[12] 300[6])
    defparam i11292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11293_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n11648), .I3(GND_net), .O(n15868));   // verilog/coms.v(127[12] 300[6])
    defparam i11293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11294_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n11648), .I3(GND_net), .O(n15869));   // verilog/coms.v(127[12] 300[6])
    defparam i11294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11295_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n11648), .I3(GND_net), .O(n15870));   // verilog/coms.v(127[12] 300[6])
    defparam i11295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11296_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n11648), .I3(GND_net), .O(n15871));   // verilog/coms.v(127[12] 300[6])
    defparam i11296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11297_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n11648), .I3(GND_net), .O(n15872));   // verilog/coms.v(127[12] 300[6])
    defparam i11297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11298_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n11648), .I3(GND_net), .O(n15873));   // verilog/coms.v(127[12] 300[6])
    defparam i11298_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_541_17 (.CI(n22333), .I0(n30633), .I1(n10), .CO(n22334));
    SB_LUT4 i11299_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n11648), .I3(GND_net), .O(n15874));   // verilog/coms.v(127[12] 300[6])
    defparam i11299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11300_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n11648), .I3(GND_net), .O(n15875));   // verilog/coms.v(127[12] 300[6])
    defparam i11300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11301_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n11648), .I3(GND_net), .O(n15876));   // verilog/coms.v(127[12] 300[6])
    defparam i11301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11302_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n11648), .I3(GND_net), .O(n15877));   // verilog/coms.v(127[12] 300[6])
    defparam i11302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11303_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n11648), .I3(GND_net), .O(n15878));   // verilog/coms.v(127[12] 300[6])
    defparam i11303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11304_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n11648), 
            .I3(GND_net), .O(n15879));   // verilog/coms.v(127[12] 300[6])
    defparam i11304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11305_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n11648), 
            .I3(GND_net), .O(n15880));   // verilog/coms.v(127[12] 300[6])
    defparam i11305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_16_lut (.I0(duty[14]), .I1(n30633), .I2(n11), .I3(n22332), 
            .O(pwm_setpoint_22__N_3[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11120_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n4772), .I3(GND_net), .O(n15695));   // verilog/coms.v(127[12] 300[6])
    defparam i11120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1637 (.I0(n26611), .I1(n14253), .I2(n27374), 
            .I3(n771), .O(n28987));
    defparam i3_4_lut_adj_1637.LUT_INIT = 16'hafbf;
    SB_LUT4 i1_4_lut_adj_1638 (.I0(n63_adj_4791), .I1(n28987), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n9520), .O(n25861));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1638.LUT_INIT = 16'hd5dd;
    SB_LUT4 i11122_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n28904), 
            .I3(GND_net), .O(n15697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11187_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15762));   // verilog/coms.v(127[12] 300[6])
    defparam i11187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11123_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_4871[1]), .I2(n8439), 
            .I3(n4_adj_4805), .O(n15698));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11123_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_4871[1]), .I1(r_SM_Main_adj_4871[0]), 
            .I2(r_SM_Main_adj_4871[2]), .I3(r_SM_Main_2__N_3497[1]), .O(n31237));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1_4_lut_4_lut (.I0(n14253), .I1(n63), .I2(n771), .I3(n26561), 
            .O(n5_adj_4769));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hcc04;
    SB_LUT4 i11124_3_lut (.I0(quadB_debounced_adj_4793), .I1(reg_B_adj_4883[0]), 
            .I2(n28888), .I3(GND_net), .O(n15699));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11125_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n15460), .I3(GND_net), .O(n15700));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i11125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11126_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n1929), .I3(GND_net), .O(n15701));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11306_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n11648), 
            .I3(GND_net), .O(n15881));   // verilog/coms.v(127[12] 300[6])
    defparam i11306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11307_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n11648), 
            .I3(GND_net), .O(n15882));   // verilog/coms.v(127[12] 300[6])
    defparam i11307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11308_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n11648), 
            .I3(GND_net), .O(n15883));   // verilog/coms.v(127[12] 300[6])
    defparam i11308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11309_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n11648), 
            .I3(GND_net), .O(n15884));   // verilog/coms.v(127[12] 300[6])
    defparam i11309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11310_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n11648), 
            .I3(GND_net), .O(n15885));   // verilog/coms.v(127[12] 300[6])
    defparam i11310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11311_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n11648), 
            .I3(GND_net), .O(n15886));   // verilog/coms.v(127[12] 300[6])
    defparam i11311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11312_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n11648), 
            .I3(GND_net), .O(n15887));   // verilog/coms.v(127[12] 300[6])
    defparam i11312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11313_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n11648), 
            .I3(GND_net), .O(n15888));   // verilog/coms.v(127[12] 300[6])
    defparam i11313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11314_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n11648), 
            .I3(GND_net), .O(n15889));   // verilog/coms.v(127[12] 300[6])
    defparam i11314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11315_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n11648), 
            .I3(GND_net), .O(n15890));   // verilog/coms.v(127[12] 300[6])
    defparam i11315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11316_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n11648), 
            .I3(GND_net), .O(n15891));   // verilog/coms.v(127[12] 300[6])
    defparam i11316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11317_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n11648), 
            .I3(GND_net), .O(n15892));   // verilog/coms.v(127[12] 300[6])
    defparam i11317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11318_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n11648), 
            .I3(GND_net), .O(n15893));   // verilog/coms.v(127[12] 300[6])
    defparam i11318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11319_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n11648), 
            .I3(GND_net), .O(n15894));   // verilog/coms.v(127[12] 300[6])
    defparam i11319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11320_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n11648), 
            .I3(GND_net), .O(n15895));   // verilog/coms.v(127[12] 300[6])
    defparam i11320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11321_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n11648), 
            .I3(GND_net), .O(n15896));   // verilog/coms.v(127[12] 300[6])
    defparam i11321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11322_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n11648), 
            .I3(GND_net), .O(n15897));   // verilog/coms.v(127[12] 300[6])
    defparam i11322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11323_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n11648), 
            .I3(GND_net), .O(n15898));   // verilog/coms.v(127[12] 300[6])
    defparam i11323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11324_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n11648), 
            .I3(GND_net), .O(n15899));   // verilog/coms.v(127[12] 300[6])
    defparam i11324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11325_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n11648), 
            .I3(GND_net), .O(n15900));   // verilog/coms.v(127[12] 300[6])
    defparam i11325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11326_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n11648), 
            .I3(GND_net), .O(n15901));   // verilog/coms.v(127[12] 300[6])
    defparam i11326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11327_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n11648), 
            .I3(GND_net), .O(n15902));   // verilog/coms.v(127[12] 300[6])
    defparam i11327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11328_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n11648), .I3(GND_net), .O(n15903));   // verilog/coms.v(127[12] 300[6])
    defparam i11328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11329_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n11648), .I3(GND_net), .O(n15904));   // verilog/coms.v(127[12] 300[6])
    defparam i11329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11330_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n11648), .I3(GND_net), .O(n15905));   // verilog/coms.v(127[12] 300[6])
    defparam i11330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11331_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n11648), .I3(GND_net), .O(n15906));   // verilog/coms.v(127[12] 300[6])
    defparam i11331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11332_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n11648), .I3(GND_net), .O(n15907));   // verilog/coms.v(127[12] 300[6])
    defparam i11332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11333_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n11648), .I3(GND_net), .O(n15908));   // verilog/coms.v(127[12] 300[6])
    defparam i11333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11334_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n11648), .I3(GND_net), .O(n15909));   // verilog/coms.v(127[12] 300[6])
    defparam i11334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11335_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n11648), .I3(GND_net), .O(n15910));   // verilog/coms.v(127[12] 300[6])
    defparam i11335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11336_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n11648), .I3(GND_net), .O(n15911));   // verilog/coms.v(127[12] 300[6])
    defparam i11336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11337_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n11648), .I3(GND_net), .O(n15912));   // verilog/coms.v(127[12] 300[6])
    defparam i11337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11338_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n11648), .I3(GND_net), .O(n15913));   // verilog/coms.v(127[12] 300[6])
    defparam i11338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11339_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n11648), .I3(GND_net), .O(n15914));   // verilog/coms.v(127[12] 300[6])
    defparam i11339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11340_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n11648), .I3(GND_net), .O(n15915));   // verilog/coms.v(127[12] 300[6])
    defparam i11340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11341_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n11648), .I3(GND_net), .O(n15916));   // verilog/coms.v(127[12] 300[6])
    defparam i11341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11342_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n11648), .I3(GND_net), .O(n15917));   // verilog/coms.v(127[12] 300[6])
    defparam i11342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11343_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n11648), .I3(GND_net), .O(n15918));   // verilog/coms.v(127[12] 300[6])
    defparam i11343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11344_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n11648), .I3(GND_net), .O(n15919));   // verilog/coms.v(127[12] 300[6])
    defparam i11344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11345_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n11648), .I3(GND_net), .O(n15920));   // verilog/coms.v(127[12] 300[6])
    defparam i11345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11346_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n11648), .I3(GND_net), .O(n15921));   // verilog/coms.v(127[12] 300[6])
    defparam i11346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11347_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n11648), .I3(GND_net), .O(n15922));   // verilog/coms.v(127[12] 300[6])
    defparam i11347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11348_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n11648), .I3(GND_net), .O(n15923));   // verilog/coms.v(127[12] 300[6])
    defparam i11348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11349_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n11648), .I3(GND_net), .O(n15924));   // verilog/coms.v(127[12] 300[6])
    defparam i11349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11350_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n11648), .I3(GND_net), .O(n15925));   // verilog/coms.v(127[12] 300[6])
    defparam i11350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11351_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n11648), .I3(GND_net), .O(n15926));   // verilog/coms.v(127[12] 300[6])
    defparam i11351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11352_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n11648), .I3(GND_net), .O(n15927));   // verilog/coms.v(127[12] 300[6])
    defparam i11352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11353_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n11648), .I3(GND_net), .O(n15928));   // verilog/coms.v(127[12] 300[6])
    defparam i11353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11354_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n11648), .I3(GND_net), .O(n15929));   // verilog/coms.v(127[12] 300[6])
    defparam i11354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11355_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n11648), .I3(GND_net), .O(n15930));   // verilog/coms.v(127[12] 300[6])
    defparam i11355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11356_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n11648), .I3(GND_net), .O(n15931));   // verilog/coms.v(127[12] 300[6])
    defparam i11356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11357_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n11648), .I3(GND_net), .O(n15932));   // verilog/coms.v(127[12] 300[6])
    defparam i11357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11358_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n11648), .I3(GND_net), .O(n15933));   // verilog/coms.v(127[12] 300[6])
    defparam i11358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11359_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n11648), .I3(GND_net), .O(n15934));   // verilog/coms.v(127[12] 300[6])
    defparam i11359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11360_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n11648), .I3(GND_net), .O(n15935));   // verilog/coms.v(127[12] 300[6])
    defparam i11360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11361_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n11648), .I3(GND_net), .O(n15936));   // verilog/coms.v(127[12] 300[6])
    defparam i11361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11362_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n11648), .I3(GND_net), .O(n15937));   // verilog/coms.v(127[12] 300[6])
    defparam i11362_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_26[0]));   // verilog/TinyFPGA_B.v(202[10] 204[6])
    SB_LUT4 i11363_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n11648), .I3(GND_net), .O(n15938));   // verilog/coms.v(127[12] 300[6])
    defparam i11363_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i11364_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n11648), .I3(GND_net), .O(n15939));   // verilog/coms.v(127[12] 300[6])
    defparam i11364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11365_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n11648), .I3(GND_net), .O(n15940));   // verilog/coms.v(127[12] 300[6])
    defparam i11365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11366_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n11648), .I3(GND_net), .O(n15941));   // verilog/coms.v(127[12] 300[6])
    defparam i11366_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_541_16 (.CI(n22332), .I0(n30633), .I1(n11), .CO(n22333));
    SB_LUT4 i11367_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n11648), .I3(GND_net), .O(n15942));   // verilog/coms.v(127[12] 300[6])
    defparam i11367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11368_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n11648), .I3(GND_net), .O(n15943));   // verilog/coms.v(127[12] 300[6])
    defparam i11368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11369_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n11648), .I3(GND_net), .O(n15944));   // verilog/coms.v(127[12] 300[6])
    defparam i11369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11370_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n11648), .I3(GND_net), .O(n15945));   // verilog/coms.v(127[12] 300[6])
    defparam i11370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11371_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n11648), .I3(GND_net), .O(n15946));   // verilog/coms.v(127[12] 300[6])
    defparam i11371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11372_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n11648), .I3(GND_net), .O(n15947));   // verilog/coms.v(127[12] 300[6])
    defparam i11372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11373_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n11648), .I3(GND_net), .O(n15948));   // verilog/coms.v(127[12] 300[6])
    defparam i11373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11374_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n11648), .I3(GND_net), .O(n15949));   // verilog/coms.v(127[12] 300[6])
    defparam i11374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_15_lut (.I0(duty[13]), .I1(n30633), .I2(n12), .I3(n22331), 
            .O(pwm_setpoint_22__N_3[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11375_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n11648), .I3(GND_net), .O(n15950));   // verilog/coms.v(127[12] 300[6])
    defparam i11375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11376_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n4774), .I3(GND_net), .O(n15951));   // verilog/coms.v(127[12] 300[6])
    defparam i11376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11377_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n4774), .I3(GND_net), .O(n15952));   // verilog/coms.v(127[12] 300[6])
    defparam i11377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11378_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n4774), .I3(GND_net), .O(n15953));   // verilog/coms.v(127[12] 300[6])
    defparam i11378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11379_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n4774), .I3(GND_net), .O(n15954));   // verilog/coms.v(127[12] 300[6])
    defparam i11379_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_541_15 (.CI(n22331), .I0(n30633), .I1(n12), .CO(n22332));
    SB_LUT4 i11380_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n4774), .I3(GND_net), .O(n15955));   // verilog/coms.v(127[12] 300[6])
    defparam i11380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11381_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n4774), .I3(GND_net), .O(n15956));   // verilog/coms.v(127[12] 300[6])
    defparam i11381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11382_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n4774), .I3(GND_net), .O(n15957));   // verilog/coms.v(127[12] 300[6])
    defparam i11382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11383_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n4774), .I3(GND_net), .O(n15958));   // verilog/coms.v(127[12] 300[6])
    defparam i11383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_541_14_lut (.I0(duty[12]), .I1(n30633), .I2(n13), .I3(n22330), 
            .O(pwm_setpoint_22__N_3[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_541_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11384_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n4774), .I3(GND_net), .O(n15959));   // verilog/coms.v(127[12] 300[6])
    defparam i11384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11385_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n4774), .I3(GND_net), .O(n15960));   // verilog/coms.v(127[12] 300[6])
    defparam i11385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11386_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n4774), .I3(GND_net), .O(n15961));   // verilog/coms.v(127[12] 300[6])
    defparam i11386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11387_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n4774), .I3(GND_net), .O(n15962));   // verilog/coms.v(127[12] 300[6])
    defparam i11387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11388_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n4774), .I3(GND_net), .O(n15963));   // verilog/coms.v(127[12] 300[6])
    defparam i11388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11389_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n4774), .I3(GND_net), .O(n15964));   // verilog/coms.v(127[12] 300[6])
    defparam i11389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11390_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n4774), .I3(GND_net), .O(n15965));   // verilog/coms.v(127[12] 300[6])
    defparam i11390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11391_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n4774), .I3(GND_net), .O(n15966));   // verilog/coms.v(127[12] 300[6])
    defparam i11391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11392_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n4774), .I3(GND_net), .O(n15967));   // verilog/coms.v(127[12] 300[6])
    defparam i11392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11393_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n4774), .I3(GND_net), .O(n15968));   // verilog/coms.v(127[12] 300[6])
    defparam i11393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11394_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n4774), .I3(GND_net), .O(n15969));   // verilog/coms.v(127[12] 300[6])
    defparam i11394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11395_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n4774), .I3(GND_net), .O(n15970));   // verilog/coms.v(127[12] 300[6])
    defparam i11395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11396_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n4774), .I3(GND_net), .O(n15971));   // verilog/coms.v(127[12] 300[6])
    defparam i11396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11397_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n4774), .I3(GND_net), .O(n15972));   // verilog/coms.v(127[12] 300[6])
    defparam i11397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11398_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n4774), .I3(GND_net), .O(n15973));   // verilog/coms.v(127[12] 300[6])
    defparam i11398_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n22552), .I0(encoder1_position[17]), 
            .I1(n8_adj_4773), .CO(n22553));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4774), .I3(n22551), .O(displacement_23__N_26[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    motorControl control (.\Kp[6] (Kp[6]), .GND_net(GND_net), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .motor_state({motor_state}), .IntegralLimit({IntegralLimit}), 
            .duty({duty}), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), 
            .PWMLimit({PWMLimit}), .\Kp[3] (Kp[3]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
            .\Ki[11] (Ki[11]), .\Ki[8] (Ki[8]), .\Kp[9] (Kp[9]), .\Ki[1] (Ki[1]), 
            .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), 
            .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Kp[4] (Kp[4]), 
            .\Kp[5] (Kp[5]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), 
            .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .setpoint({setpoint}), 
            .\Ki[12] (Ki[12]), .\Ki[15] (Ki[15]), .\Ki[14] (Ki[14]), .\Ki[13] (Ki[13]), 
            .clk32MHz(clk32MHz), .VCC_net(VCC_net), .n25(n25), .n30633(n30633)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(172[16] 184[4])
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n22551), .I0(encoder1_position[16]), 
            .I1(n9_adj_4774), .CO(n22552));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4775), .I3(n22550), .O(displacement_23__N_26[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n22550), .I0(encoder1_position[15]), 
            .I1(n10_adj_4775), .CO(n22551));
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.data_o({quadA_debounced_adj_4792, 
            quadB_debounced_adj_4793}), .GND_net(GND_net), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n28888(n28888), .reg_B({reg_B_adj_4883}), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .VCC_net(VCC_net), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n16185(n16185), .n15699(n15699)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(195[15] 200[4])
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4776), .I3(n22549), .O(displacement_23__N_26[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n22549), .I0(encoder1_position[14]), 
            .I1(n11_adj_4776), .CO(n22550));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4777), .I3(n22548), .O(displacement_23__N_26[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n22548), .I0(encoder1_position[13]), 
            .I1(n12_adj_4777), .CO(n22549));
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4778), .I3(n22547), .O(displacement_23__N_26[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n22547), .I0(encoder1_position[12]), 
            .I1(n13_adj_4778), .CO(n22548));
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4779), .I3(n22546), .O(displacement_23__N_26[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_541_14 (.CI(n22330), .I0(n30633), .I1(n13), .CO(n22331));
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n22546), .I0(encoder1_position[11]), 
            .I1(n14_adj_4779), .CO(n22547));
    \pwm(32000000,20000,8000000,23,1)  PWM (.INHA_c_0(INHA_c_0), .clk32MHz(clk32MHz), 
            .\half_duty_new[0] (half_duty_new[0]), .n15460(n15460), .\half_duty[0][0] (\half_duty[0] [0]), 
            .GND_net(GND_net), .\half_duty[0][1] (\half_duty[0] [1]), .\half_duty[0][2] (\half_duty[0] [2]), 
            .\half_duty[0][3] (\half_duty[0] [3]), .\half_duty[0][4] (\half_duty[0] [4]), 
            .\half_duty[0][5] (\half_duty[0] [5]), .\half_duty[0][6] (\half_duty[0] [6]), 
            .\half_duty[0][7] (\half_duty[0] [7]), .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint}), 
            .\half_duty_new[1] (half_duty_new[1]), .\half_duty_new[2] (half_duty_new[2]), 
            .\half_duty_new[3] (half_duty_new[3]), .\half_duty_new[4] (half_duty_new[4]), 
            .\half_duty_new[5] (half_duty_new[5]), .\half_duty_new[6] (half_duty_new[6]), 
            .\half_duty_new[7] (half_duty_new[7]), .n16195(n16195), .n16194(n16194), 
            .n16193(n16193), .n16192(n16192), .n16191(n16191), .n16190(n16190), 
            .n16189(n16189), .n15700(n15700));   // verilog/TinyFPGA_B.v(90[42] 96[3])
    coms neopxl_color_23__I_0 (.\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .GND_net(GND_net), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .n15762(n15762), 
         .\data_in[3] ({\data_in[3] }), .clk32MHz(clk32MHz), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n15761(n15761), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n15760(n15760), .\data_in[2] ({\data_in[2] }), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .setpoint({setpoint}), .n15759(n15759), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .n15758(n15758), .n15757(n15757), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .n15756(n15756), .n15755(n15755), 
         .rx_data({rx_data}), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n15754(n15754), .n15753(n15753), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .n15752(n15752), .\data_in[1] ({\data_in[1] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .n15751(n15751), .rx_data_ready(rx_data_ready), 
         .n15750(n15750), .n15749(n15749), .n15748(n15748), .n15747(n15747), 
         .n14288(n14288), .n771(n771), .n9520(n9520), .n4609(n4609), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n14253(n14253), 
         .n123(n123), .n63(n63), .n26561(n26561), .n14291(n14291), .n4677(n4677), 
         .n14254(n14254), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .n15746(n15746), .\FRAME_MATCHER.state_31__N_2672[1] (\FRAME_MATCHER.state_31__N_2672 [1]), 
         .n8595(n8595), .n122(n122), .\FRAME_MATCHER.state_31__N_2672[2] (\FRAME_MATCHER.state_31__N_2672 [2]), 
         .n4452(n4452), .n7(n7_adj_4803), .n2649(n2649), .n8(n8_adj_4804), 
         .n14279(n14279), .n15745(n15745), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .tx_active(tx_active), .n15744(n15744), .\data_in[0] ({\data_in[0] }), 
         .n15743(n15743), .n15742(n15742), .n27362(n27362), .n4772(n4772), 
         .n15741(n15741), .LED_c(LED_c), .n27374(n27374), .n15740(n15740), 
         .n15739(n15739), .n15738(n15738), .n15737(n15737), .IntegralLimit({IntegralLimit}), 
         .n15736(n15736), .n15735(n15735), .n15734(n15734), .n15733(n15733), 
         .n15732(n15732), .n15731(n15731), .n15730(n15730), .n15729(n15729), 
         .n15728(n15728), .n15727(n15727), .n15726(n15726), .n15725(n15725), 
         .n15724(n15724), .n15723(n15723), .n15722(n15722), .n15721(n15721), 
         .n15720(n15720), .n15719(n15719), .n15718(n15718), .n15717(n15717), 
         .n15716(n15716), .n15715(n15715), .n63_adj_3(n63_adj_4791), .n27965(n27965), 
         .n25997(n25997), .DE_c(DE_c), .n31238(n31238), .n31239(n31239), 
         .n16178(n16178), .PWMLimit({PWMLimit}), .n16177(n16177), .n16176(n16176), 
         .n16175(n16175), .n16174(n16174), .n16173(n16173), .n16172(n16172), 
         .n16171(n16171), .n16170(n16170), .n16169(n16169), .n16168(n16168), 
         .n16167(n16167), .n16166(n16166), .n16165(n16165), .n16164(n16164), 
         .n16163(n16163), .n16162(n16162), .n16161(n16161), .n16160(n16160), 
         .n16159(n16159), .n16158(n16158), .n16157(n16157), .n16156(n16156), 
         .n16155(n16155), .control_mode({control_mode}), .n16154(n16154), 
         .n16153(n16153), .n16152(n16152), .n16151(n16151), .n16150(n16150), 
         .n16149(n16149), .n15973(n15973), .neopxl_color({neopxl_color}), 
         .n15972(n15972), .n15971(n15971), .n15970(n15970), .n15969(n15969), 
         .n15968(n15968), .n15967(n15967), .n15966(n15966), .n15965(n15965), 
         .n15964(n15964), .n15963(n15963), .n15962(n15962), .n15961(n15961), 
         .n15960(n15960), .n15959(n15959), .n15958(n15958), .n15957(n15957), 
         .n15956(n15956), .n15955(n15955), .n15954(n15954), .n15953(n15953), 
         .n15952(n15952), .n15951(n15951), .n15950(n15950), .n15949(n15949), 
         .n15948(n15948), .n15947(n15947), .n15946(n15946), .n15945(n15945), 
         .n15944(n15944), .n15943(n15943), .n15942(n15942), .n15941(n15941), 
         .n15940(n15940), .n15939(n15939), .n15938(n15938), .n15937(n15937), 
         .n15936(n15936), .n15935(n15935), .n15934(n15934), .n15933(n15933), 
         .n15932(n15932), .n15931(n15931), .n15930(n15930), .n15929(n15929), 
         .n15928(n15928), .n15927(n15927), .n15926(n15926), .n15925(n15925), 
         .n15924(n15924), .n15923(n15923), .n15922(n15922), .n15921(n15921), 
         .n15920(n15920), .n15919(n15919), .n15918(n15918), .n15917(n15917), 
         .n15916(n15916), .n15915(n15915), .n15914(n15914), .n15913(n15913), 
         .n15912(n15912), .n15911(n15911), .n15910(n15910), .n15909(n15909), 
         .n15908(n15908), .n15907(n15907), .n15906(n15906), .n15905(n15905), 
         .n15904(n15904), .n15903(n15903), .n15902(n15902), .n15901(n15901), 
         .n15900(n15900), .n15899(n15899), .n15898(n15898), .n15897(n15897), 
         .n15896(n15896), .n15895(n15895), .n15894(n15894), .n15893(n15893), 
         .n15892(n15892), .n15891(n15891), .n15890(n15890), .n15889(n15889), 
         .n15888(n15888), .n15887(n15887), .n15886(n15886), .n15885(n15885), 
         .n15884(n15884), .n15883(n15883), .n15882(n15882), .n15881(n15881), 
         .n25861(n25861), .n15695(n15695), .n15880(n15880), .n15879(n15879), 
         .n15878(n15878), .n15877(n15877), .n15876(n15876), .n15875(n15875), 
         .n15874(n15874), .n15873(n15873), .n15872(n15872), .n15871(n15871), 
         .n15870(n15870), .n15869(n15869), .n15868(n15868), .n15867(n15867), 
         .n15866(n15866), .n15865(n15865), .n15864(n15864), .n15863(n15863), 
         .n15862(n15862), .n15861(n15861), .n15860(n15860), .n15859(n15859), 
         .n15858(n15858), .n15857(n15857), .n15856(n15856), .n15855(n15855), 
         .n15854(n15854), .n15853(n15853), .n15852(n15852), .n15851(n15851), 
         .n15850(n15850), .n15849(n15849), .n15848(n15848), .n15694(n15694), 
         .n15692(n15692), .n15691(n15691), .\Ki[0] (Ki[0]), .n15690(n15690), 
         .\Kp[0] (Kp[0]), .n15689(n15689), .n15847(n15847), .n15846(n15846), 
         .n15845(n15845), .n15844(n15844), .n15843(n15843), .n15842(n15842), 
         .n15841(n15841), .n15682(n15682), .n15840(n15840), .n15839(n15839), 
         .n15838(n15838), .n15837(n15837), .n15836(n15836), .n15835(n15835), 
         .n15834(n15834), .n15833(n15833), .n15832(n15832), .n15831(n15831), 
         .n15830(n15830), .n15829(n15829), .n15828(n15828), .n15827(n15827), 
         .n15826(n15826), .n15825(n15825), .n15824(n15824), .n15823(n15823), 
         .n15822(n15822), .n15821(n15821), .n15820(n15820), .n15819(n15819), 
         .n15818(n15818), .n15817(n15817), .n11648(n11648), .n4774(n4774), 
         .n15816(n15816), .n15815(n15815), .n15814(n15814), .n15813(n15813), 
         .n15812(n15812), .n15811(n15811), .n15810(n15810), .n15809(n15809), 
         .n15808(n15808), .n15807(n15807), .n15806(n15806), .n15805(n15805), 
         .n15804(n15804), .n15803(n15803), .n15802(n15802), .n15801(n15801), 
         .n15800(n15800), .n15799(n15799), .n15798(n15798), .\Ki[15] (Ki[15]), 
         .n15797(n15797), .\Ki[14] (Ki[14]), .n15796(n15796), .\Ki[13] (Ki[13]), 
         .n15795(n15795), .\Ki[12] (Ki[12]), .n15794(n15794), .\Ki[11] (Ki[11]), 
         .n15793(n15793), .\Ki[10] (Ki[10]), .n15792(n15792), .\Ki[9] (Ki[9]), 
         .n15791(n15791), .\Ki[8] (Ki[8]), .n15790(n15790), .\Ki[7] (Ki[7]), 
         .n15789(n15789), .\Ki[6] (Ki[6]), .n15788(n15788), .\Ki[5] (Ki[5]), 
         .n15787(n15787), .\Ki[4] (Ki[4]), .n15786(n15786), .\Ki[3] (Ki[3]), 
         .n15785(n15785), .\Ki[2] (Ki[2]), .n15784(n15784), .\Ki[1] (Ki[1]), 
         .n15783(n15783), .\Kp[15] (Kp[15]), .n15782(n15782), .\Kp[14] (Kp[14]), 
         .n15781(n15781), .\Kp[13] (Kp[13]), .n15780(n15780), .\Kp[12] (Kp[12]), 
         .n15779(n15779), .\Kp[11] (Kp[11]), .n15778(n15778), .\Kp[10] (Kp[10]), 
         .n15777(n15777), .\Kp[9] (Kp[9]), .n15776(n15776), .\Kp[8] (Kp[8]), 
         .n15775(n15775), .\Kp[7] (Kp[7]), .n15774(n15774), .\Kp[6] (Kp[6]), 
         .n15773(n15773), .\Kp[5] (Kp[5]), .n15772(n15772), .\Kp[4] (Kp[4]), 
         .n15771(n15771), .\Kp[3] (Kp[3]), .n15770(n15770), .\Kp[2] (Kp[2]), 
         .n15769(n15769), .\Kp[1] (Kp[1]), .n15768(n15768), .n15767(n15767), 
         .n15766(n15766), .n15765(n15765), .n15764(n15764), .n15763(n15763), 
         .\r_Bit_Index[0] (r_Bit_Index_adj_4873[0]), .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_4871}), 
         .\r_SM_Main_2__N_3497[1] (r_SM_Main_2__N_3497[1]), .n27464(n27464), 
         .n27476(n27476), .n4(n4_adj_4805), .VCC_net(VCC_net), .n15704(n15704), 
         .n8439(n8439), .n31237(n31237), .n15698(n15698), .tx_enable(tx_enable), 
         .\r_SM_Main_2__N_3426[2] (r_SM_Main_2__N_3426[2]), .r_SM_Main_adj_11({r_SM_Main}), 
         .n26557(n26557), .\r_Bit_Index[0]_adj_7 (r_Bit_Index[0]), .r_Rx_Data(r_Rx_Data), 
         .RX_N_2(RX_N_2), .n14264(n14264), .n18753(n18753), .n14259(n14259), 
         .n4_adj_8(n4_adj_4768), .n15508(n15508), .n15619(n15619), .n4_adj_9(n4), 
         .n4_adj_10(n4_adj_4763), .n15711(n15711), .n16227(n16227), .n15707(n15707), 
         .n26153(n26153), .n15686(n15686), .n15685(n15685), .n15684(n15684), 
         .n15683(n15683), .n15681(n15681), .n15680(n15680)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(138[8] 161[4])
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4780), .I3(n22545), .O(displacement_23__N_26[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, clk32MHz, 
            data_o, n28904, reg_B, VCC_net, ENCODER0_B_c_0, n16183, 
            n15697, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output n28904;
    output [1:0]reg_B;
    input VCC_net;
    input ENCODER0_B_c_0;
    input n16183;
    input n15697;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2856;
    
    wire n2852, n22391, n22392, n22390, n22389, n22388, n22387, 
        count_enable, B_delayed, A_delayed, n22386, n22385, count_direction, 
        n22384, n22407, n22406, n22405, n22404, n22403, n22402, 
        n22401, n22400, n22399, n22398, n22397, n22396, n22395, 
        n22394, n22393;
    
    SB_LUT4 add_610_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2852), 
            .I3(n22391), .O(n2856[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_9 (.CI(n22391), .I0(encoder0_position[7]), .I1(n2852), 
            .CO(n22392));
    SB_LUT4 add_610_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2852), 
            .I3(n22390), .O(n2856[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_8 (.CI(n22390), .I0(encoder0_position[6]), .I1(n2852), 
            .CO(n22391));
    SB_LUT4 add_610_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2852), 
            .I3(n22389), .O(n2856[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_7 (.CI(n22389), .I0(encoder0_position[5]), .I1(n2852), 
            .CO(n22390));
    SB_LUT4 add_610_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2852), 
            .I3(n22388), .O(n2856[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_6 (.CI(n22388), .I0(encoder0_position[4]), .I1(n2852), 
            .CO(n22389));
    SB_LUT4 add_610_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2852), 
            .I3(n22387), .O(n2856[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_5 (.CI(n22387), .I0(encoder0_position[3]), .I1(n2852), 
            .CO(n22388));
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_610_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2852), 
            .I3(n22386), .O(n2856[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_4 (.CI(n22386), .I0(encoder0_position[2]), .I1(n2852), 
            .CO(n22387));
    SB_LUT4 add_610_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2852), 
            .I3(n22385), .O(n2856[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_3 (.CI(n22385), .I0(encoder0_position[1]), .I1(n2852), 
            .CO(n22386));
    SB_LUT4 add_610_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n22384), .O(n2856[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_2 (.CI(n22384), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n22385));
    SB_CARRY add_610_1 (.CI(GND_net), .I0(n2852), .I1(n2852), .CO(n22384));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_610_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2852), 
            .I3(n22407), .O(n2856[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_610_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2852), 
            .I3(n22406), .O(n2856[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_24 (.CI(n22406), .I0(encoder0_position[22]), .I1(n2852), 
            .CO(n22407));
    SB_LUT4 add_610_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2852), 
            .I3(n22405), .O(n2856[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_610_23 (.CI(n22405), .I0(encoder0_position[21]), .I1(n2852), 
            .CO(n22406));
    SB_LUT4 add_610_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2852), 
            .I3(n22404), .O(n2856[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_22 (.CI(n22404), .I0(encoder0_position[20]), .I1(n2852), 
            .CO(n22405));
    SB_LUT4 add_610_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2852), 
            .I3(n22403), .O(n2856[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_21 (.CI(n22403), .I0(encoder0_position[19]), .I1(n2852), 
            .CO(n22404));
    SB_LUT4 add_610_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2852), 
            .I3(n22402), .O(n2856[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_20 (.CI(n22402), .I0(encoder0_position[18]), .I1(n2852), 
            .CO(n22403));
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[23]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_610_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2852), 
            .I3(n22401), .O(n2856[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_19 (.CI(n22401), .I0(encoder0_position[17]), .I1(n2852), 
            .CO(n22402));
    SB_LUT4 add_610_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2852), 
            .I3(n22400), .O(n2856[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_18 (.CI(n22400), .I0(encoder0_position[16]), .I1(n2852), 
            .CO(n22401));
    SB_LUT4 add_610_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2852), 
            .I3(n22399), .O(n2856[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_17 (.CI(n22399), .I0(encoder0_position[15]), .I1(n2852), 
            .CO(n22400));
    SB_LUT4 add_610_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2852), 
            .I3(n22398), .O(n2856[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_16 (.CI(n22398), .I0(encoder0_position[14]), .I1(n2852), 
            .CO(n22399));
    SB_LUT4 add_610_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2852), 
            .I3(n22397), .O(n2856[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_15 (.CI(n22397), .I0(encoder0_position[13]), .I1(n2852), 
            .CO(n22398));
    SB_LUT4 add_610_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2852), 
            .I3(n22396), .O(n2856[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_14 (.CI(n22396), .I0(encoder0_position[12]), .I1(n2852), 
            .CO(n22397));
    SB_LUT4 i903_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2852));   // quad.v(37[5] 40[8])
    defparam i903_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_610_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2852), 
            .I3(n22395), .O(n2856[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_13 (.CI(n22395), .I0(encoder0_position[11]), .I1(n2852), 
            .CO(n22396));
    SB_LUT4 add_610_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2852), 
            .I3(n22394), .O(n2856[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_12 (.CI(n22394), .I0(encoder0_position[10]), .I1(n2852), 
            .CO(n22395));
    SB_LUT4 add_610_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2852), 
            .I3(n22393), .O(n2856[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_11 (.CI(n22393), .I0(encoder0_position[9]), .I1(n2852), 
            .CO(n22394));
    SB_LUT4 add_610_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2852), 
            .I3(n22392), .O(n2856[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_610_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_610_10 (.CI(n22392), .I0(encoder0_position[8]), .I1(n2852), 
            .CO(n22393));
    \grp_debouncer(2,100)_U0  debounce (.n28904(n28904), .reg_B({reg_B}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n16183(n16183), .data_o({data_o}), 
            .n15697(n15697), .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (n28904, reg_B, GND_net, clk32MHz, 
            VCC_net, ENCODER0_B_c_0, n16183, data_o, n15697, ENCODER0_A_c_1);
    output n28904;
    output [1:0]reg_B;
    input GND_net;
    input clk32MHz;
    input VCC_net;
    input ENCODER0_B_c_0;
    input n16183;
    output [1:0]data_o;
    input n15697;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3740;
    wire [6:0]n33;
    
    wire n22867, n22866, n22865, n22864, n22863, n22862;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n28904));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n28904), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1214__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 cnt_reg_1214_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n22867), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1214_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n22866), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1214_add_4_7 (.CI(n22866), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n22867));
    SB_LUT4 cnt_reg_1214_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n22865), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1214_add_4_6 (.CI(n22865), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n22866));
    SB_LUT4 cnt_reg_1214_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n22864), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1214_add_4_5 (.CI(n22864), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n22865));
    SB_LUT4 cnt_reg_1214_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n22863), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1214_add_4_4 (.CI(n22863), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n22864));
    SB_LUT4 cnt_reg_1214_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n22862), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1214_add_4_3 (.CI(n22862), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n22863));
    SB_LUT4 cnt_reg_1214_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1214_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1214_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n22862));
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n16183));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n15697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1214__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1214__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1214__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1214__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1214__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1214__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (timer, \neo_pixel_transmitter.done , clk32MHz, GND_net, 
            VCC_net, \neo_pixel_transmitter.t0 , start, n4, \state[0] , 
            n66, LED_c, \state[1] , n1929, n19323, neopxl_color, 
            n16226, n16225, n16224, n16223, n16222, n16221, n16220, 
            n16219, n16218, n16217, n16216, n16215, n16214, n16213, 
            n16212, n16211, n16210, n16209, n16208, n16207, n16206, 
            n16205, n16204, n16203, n16202, n16201, n16200, n16199, 
            n16198, n16197, n16196, n25291, NEOPXL_c, n15701) /* synthesis syn_module_defined=1 */ ;
    output [31:0]timer;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output start;
    output n4;
    output \state[0] ;
    output n66;
    input LED_c;
    output \state[1] ;
    output n1929;
    output n19323;
    input [23:0]neopxl_color;
    input n16226;
    input n16225;
    input n16224;
    input n16223;
    input n16222;
    input n16221;
    input n16220;
    input n16219;
    input n16218;
    input n16217;
    input n16216;
    input n16215;
    input n16214;
    input n16213;
    input n16212;
    input n16211;
    input n16210;
    input n16209;
    input n16208;
    input n16207;
    input n16206;
    input n16205;
    input n16204;
    input n16203;
    input n16202;
    input n16201;
    input n16200;
    input n16199;
    input n16198;
    input n16197;
    input n16196;
    input n25291;
    output NEOPXL_c;
    input n15701;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n2291, n2192, n2225, n22622, n22435;
    wire [31:0]n1;
    
    wire n22436, n22721, n1802, n1829, n22722, n23555, n2308, 
        n2324, n23556, n2292, n2193, n22621, n2405, n2306, n23557, 
        \neo_pixel_transmitter.done_N_580 , n28956, n2396, n2297, n23566, 
        n2293, n2194, n22620, n2406, n2307;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n3209, n19329, n35, n11, n29, n51, n48, n37, n23, 
        n53, n39, n46, n27, n57, n63, n43, n47, n25, n33, 
        n47_adj_4608, n61, n45, n59, n17, n15, n55, n44, n31, 
        n41, n49, n43_adj_4609, n54, n45_adj_4610, n13, n19, n21, 
        n49_adj_4611, n23810, n24143, n23567, n30631, n4_c;
    wire [31:0]one_wire_N_523;
    
    wire n2294, n2195, n22619, n2295, n2196, n22618, n1902, n1803, 
        n22720, n2296, n2197, n22617, n1903, n1804, n22719, n2198, 
        n22616, n1904, n1805, n22718, n2298, n2199, n22615, n1905, 
        n1806, n22717, n2299, n2200, n22614, n1906, n1807, n22716, 
        n1907, n1808, n22715, n2300, n2201, n22613, n1908, n1809, 
        n22714, n2301, n2202, n22612, n1909, n1994, n1895, n1928, 
        n22713, n1995, n1896, n22712, n1996, n1897, n22711, n1997, 
        n1898, n22710, n1998, n1899, n22709, n1999, n1900, n22708, 
        n2103, n2097, n18, n2109, n19377, n2093, n2108, n2100, 
        n30, n2000, n1901, n22707, n2302, n2203, n22611, n2098, 
        n2094, n2099, n28, n2001, n22706, n2105, n2096, n2095, 
        n2102, n29_adj_4613, n2303, n2204, n22610, n2002, n22705, 
        n2304, n2205, n22609, n2003, n22704, n2101, n2107, n2104, 
        n2106, n27_adj_4614, n2126, n2305, n2206, n22608, n2207, 
        n22607, n2004, n22703, n2005, n22702, n2208, n22606, n2006, 
        n22701, n2209, n30634, n22605, n2007, n22700, n2008, n30635, 
        n22699, n2309, n2009, n2027, n22698, n22697, n2693, n2704, 
        n28_adj_4616, n2699, n2706, n2694, n2691, n38, n2709, 
        n19339, n2701, n2696, n2697, n36, n2700, n2705, n42, 
        n22696, n2702, n2690, n2689, n2708, n40, n2687, n2703, 
        n2695, n41_adj_4617, n2688, n2698, n2692, n2707, n39_adj_4618, 
        n2720;
    wire [31:0]n255;
    
    wire n15464, n15593, n2819, n30641, n22695, n2404, n23558, 
        n2403, n23559, n2397, n23565, n2407, n23560, n2398, n23564, 
        n2489, n2390, n2423, n22427, n2798, n2804, n2791, n2795, 
        n40_adj_4621, n2796, n2793, n2788, n2808, n38_adj_4622, 
        n2789, n2800, n2803, n2805, n39_adj_4623, n2792, n2787, 
        n2801, n2799, n37_adj_4624, n2786, n2797, n34, n2794, 
        n2806, n2807, n2790, n42_adj_4625, n46_adj_4626, n22694, 
        n2802, n2809, n33_adj_4627, n2918, n30640, n22693, n22692, 
        n2894, n2909, n33_adj_4629, n2885, n2900, n2891, n2889, 
        n41_adj_4630, n2895, n2887, n2906, n38_adj_4631, n2896, 
        n2893, n2890, n2899, n43_adj_4632, n2892, n2901, n2902, 
        n2908, n40_adj_4633, n2903, n2886, n46_adj_4634, n2907, 
        n2897, n2898, n2904, n39_adj_4635, n2888, n2905, n47_adj_4636, 
        n22691, n3017, n30639, n3004, n2989, n2990, n3007, n40_adj_4639, 
        n3006, n2984, n2988, n2986, n44_adj_4640, n3008, n3003, 
        n2994, n3002, n42_adj_4641, n2999, n3000, n2992, n2997, 
        n43_adj_4642, n2996, n2985, n2995, n2987, n41_adj_4643, 
        n3001, n2993, n38_adj_4644, n2998, n2991, n46_adj_4645, 
        n50, n3005, n3009, n37_adj_4646, n3116, n30638, n30637, 
        n3103, n3109, n36_adj_4647, n3104, n3094, n3095, n3097, 
        n46_adj_4648, n3084, n3089, n3083, n3105, n42_adj_4649, 
        n3086, n3091, n32_adj_4650, n3092, n3098, n3100, n3107, 
        n44_adj_4651, n3085, n3093, n50_adj_4652, n3087, n3096, 
        n3099, n48_adj_4653, n3102, n3101, n49_adj_4654, n3106, 
        n3090, n3108, n3088, n47_adj_4655, n22690, n2591, n2608, 
        n2601, n2605, n36_adj_4656, n2606, n2609, n25_adj_4657, 
        n2593, n2596, n2600, n2590, n34_adj_4658, n2490, n2391, 
        n22426, n2594, n2589, n40_adj_4659, n2602, n2588, n2604, 
        n2607, n38_adj_4660, n2598, n2603, n39_adj_4661, n2592, 
        n2597, n2595, n2599, n37_adj_4662, n2621, n30642, n30636, 
        n22689, n2408, n30632, n23554, n22688, n2491, n2392, n22425, 
        n2409, n2492, n2393, n22424, n2493, n2394, n22423, n22687, 
        n22298, n2494, n2395, n22422, n22290, n22299, n2495, n22421, 
        n22297, n2496, n22420, n22318, n22317, n22316, n2497, 
        n22419, n22291, n2498, n2399, n22418, n22296, n22315, 
        n22289, n22314, n2499, n2400, n22417, n22313, n22686, 
        n2500, n2401, n22416, n22312, n22311, n2501, n2402, n22415, 
        n22, n22465, n2502, n22414, n22685, n22295, n22310, n23563, 
        n23562, n23_adj_4664, n22464, n22684, n28_adj_4665, n22463, 
        n2503, n22413, n22683, n23561, n2504, n22412, n26, n22462, 
        n2505, n22411, n21_adj_4666, n22461, n22294, n2506, n22410, 
        n22309, n23572, n22308, n23067, n23066, n23065, n23064, 
        n2507, n22409, n23063, n22460, n22288, n23062, n23061, 
        n2508, n22408, n23060, n23059, n23058, n23057, n23056, 
        n23055, n2509, n23054, n23053, n23052, n23051, n23050, 
        n22459, n23049, n22307, n23048, n23047, n22306, n22305, 
        n23046, n23571, n22293, n23045, n23044, n23043, n23042, 
        n22458, n23041, n23040, n23039, n23038, n23037, n23036, 
        n23035, n30_adj_4667, n22457, n23034, n23033, n23032, n23031, 
        n23030, n23029, n23028, n23027, n23026, n23025, n23024, 
        n23023, n24, n22456, n27_adj_4668, n33_adj_4669, n32_adj_4670, 
        n31_adj_4671, n35_adj_4672, n37_adj_4673, n23022, n23021, 
        n23020, n23019, n25_adj_4674, n22455, n23018, n23017;
    wire [31:0]n133;
    
    wire n14_adj_4675, n23016, n13_adj_4676, n23015, n22_adj_4677, 
        n32_adj_4678, n29_adj_4679, n22454, n23014, n23013, n22453, 
        n23012, n23011, n23010, n23009, n23008, n36_adj_4680, n23007, 
        n23006, n23005, n23004, n34_adj_4681, n23003, n35_adj_4682, 
        n33_adj_4683, n23002, n24963, n23001, n19291, n27307, n23000, 
        n22999, n22998, n22997, n22996, n22995, n22994, n22993, 
        n22992, n14151, n19313, n22991, n22990, n10_adj_4685, n14275, 
        n14_adj_4686, n22452, n76, n4659, n22989, n22988, n22987, 
        n27_adj_4687, n22451, n22986, n29835, n22985, n28213, n22984, 
        n22983, n22982, n22981, n22980, n22979, n22978, n1304, 
        n1305, n10_adj_4688, n22977, n22976, n1303, n1309, n12_adj_4689, 
        n22975, n22974, n1306, n1308, n1302, n16_adj_4690, n22973, 
        n1307, n1301, n1334, n22972, n22450, n22449, n22971, n22970, 
        n22969, n22968, n22967, n22966, n22965, n22964, n22963, 
        n22448, n83, n22639, n22962, n22961, n22960, n22447, n22638, 
        n22959, n22958, n22637, n22957, n22956, n22955, n22636, 
        n22954, n18_adj_4692, n28_adj_4693, n22635, n26_adj_4694, 
        n27_adj_4695, n25_adj_4696, n22634, n22953, n22952, n22951, 
        n22950, n27317, n12884, n807, n838, n18_adj_4699, n26_adj_4700, 
        n11_adj_4701, n24_adj_4702, n19309, n25_adj_4703, n27428, 
        n29787, n20768, n19471, n27462, n29821, n15468, n23_adj_4704, 
        n19317;
    wire [4:0]color_bit_N_566;
    
    wire n30880, n30808, n29829, n30784;
    wire [3:0]state_3__N_372;
    
    wire n30949, n29081, n78, n30877, n22949, n27356, n27855, 
        n1235, n30648, n36_adj_4705, n37_adj_4706, n30823, n29210, 
        n30817, n29213, n30805, n30787, n30389, n30781, n14_adj_4707, 
        n22948, n22947, n22946, n22945, n22944, n22943, n15_adj_4708, 
        n22942, n22941, n27482, n22940, n22633, n22939, n26579, 
        n103, n22938, n22937, n22936, n1205, n1206, n1204, n1207, 
        n14_adj_4709, n1203, n1209, n9_adj_4710, n1202, n1208, n1136, 
        n30647, n30643, n22935, n22934, n22933, n22932, n22931, 
        n22930, n1106, n1104, n8_adj_4713, n1105, n1103, n1107, 
        n1108, n12_adj_4714, n1109, n1730, n30653, n1037, n30646, 
        n2_adj_4716;
    wire [31:0]n971;
    
    wire n1007, n1006, n906, n1005, n15523, n905, n8_adj_4717, 
        n12882, n1009, n1008, n29077, n6_adj_4718, n4_adj_4719, 
        n60, n608, n708, n27340, n29790, n22929, n22928, n22927, 
        n22926, n22925, n22924, n22923, n22304, n2522, n30645, 
        n22446, n22922, n30644, n22921, n22920, n22919, n22918, 
        n22632, n24_adj_4724, n34_adj_4725, n22_adj_4726, n38_adj_4727, 
        n36_adj_4728, n37_adj_4729, n22917, n35_adj_4730, n22916, 
        n22915, n22914, n22913, n22631, n22912, n1699, n1709, 
        n17_adj_4731, n22911, n22910, n22303, n22909, n1698, n1707, 
        n1703, n1705, n21_adj_4732, n1704, n1701, n1708, n20_adj_4733, 
        n1702, n1697, n24_adj_4734, n22908, n22_adj_4735, n1700, 
        n1706, n22907, n22906, n1631, n30652, n22905, n22904, 
        n22903, n22902, n22630, n22901, n22900, n30_adj_4736, n27488, 
        n4_adj_4737, n34_adj_4738, n22899, n22898, n22897, n22896, 
        n22629, n22895, n22445, n22444, n22628, n22627, n22894, 
        n22893, n22892, n22891, n22890, n22292, n22889, n22888, 
        n22887, n22886, n22885, n22884, n22626, n22883, n22443, 
        n22882, n22442, n22881, n22880, n22879, n22878, n22877, 
        n28974, n22876, n22875, n22874, n32_adj_4739, n33_adj_4740, 
        n31_adj_4741, n1608, n1606, n1604, n1603, n20_adj_4742, 
        n1602, n1609, n13_adj_4743, n1598, n1600, n18_adj_4744, 
        n22441, n1605, n1599, n22_adj_4745, n22440, n1601, n1607, 
        n22302, n12_adj_4746, n22439, n20_adj_4747, n1801, n1800, 
        n23_adj_4748, n1798, n1799, n22_adj_4749, n1797, n26_adj_4750, 
        n1796, n28_adj_4751, n32_adj_4752, n30_adj_4753, n22813, n31_adj_4754, 
        n22812, n29_adj_4755, n22811, n22810, n22809, n22808, n22807, 
        n22806, n22805, n22804, n22803, n22802, n22801, n22800, 
        n22799, n22798, n22797, n22796, n22795, n22794, n22793, 
        n23570, n22792, n22791, n22790, n22789, n22788, n22787, 
        n22786, n22785, n22784, n22783, n1400, n22782, n1401, 
        n22781, n1532, n30651, n1500, n1506, n1499, n1501, n18_adj_4756, 
        n1508, n1504, n1502, n20_adj_4757, n1505, n1509, n15_adj_4758, 
        n1402, n22780, n1503, n1507, n1433, n30650, n1407, n1406, 
        n1403, n1404, n16_adj_4760, n22779, n22778, n1408, n18_adj_4761, 
        n1409, n13_adj_4762, n1405, n30649, n27450, n22777, n22776, 
        n91, n26470, n15422, \neo_pixel_transmitter.done_N_586 , n22775, 
        n22774, n22773, n22772, n22771, n22770, n22769, n22768, 
        n22438, n22767, n22766, n22765, n22764, n22763, n22301, 
        n22762, n22761, n22760, n22759, n22758, n22757, n22756, 
        n22755, n22754, n22753, n23569, n22752, n22751, n22750, 
        n22749, n22300, n22748, n22747, n22746, n22745, n22744, 
        n22743, n22742, n22741, n22740, n22739, n22738, n22737, 
        n22736, n22735, n22437, n22734, n22625, n22733, n22732, 
        n22731, n22730, n22624, n22729, n22728, n22727, n22726, 
        n22725, n22724, n22623, n23568, n22723;
    
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n22622), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_3 (.CI(n22435), .I0(timer[1]), .I1(n1[1]), .CO(n22436));
    SB_CARRY mod_5_add_1272_10 (.CI(n22721), .I0(n1802), .I1(n1829), .CO(n22722));
    SB_CARRY mod_5_add_1607_4 (.CI(n23555), .I0(n2308), .I1(n2324), .CO(n23556));
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n22621), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n23557), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n28956), .D(\neo_pixel_transmitter.done_N_580 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n23566), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n22621), .I0(n2193), .I1(n2225), .CO(n22622));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n22620), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n23556), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n23556), .I0(n2307), .I1(n2324), .CO(n23557));
    SB_LUT4 i14762_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n19329));
    defparam i14762_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n11), .I2(n29), .I3(n51), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n37), .I1(n23), .I2(n53), .I3(n39), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n27), .I1(n57), .I2(n63), .I3(n43), .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n25), .I1(n33), .I2(n47_adj_4608), .I3(n61), 
            .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n59), .I1(n17), .I2(n15), .I3(n55), .O(n44));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n31), .I1(n41), .I2(n49), .I3(n19329), .O(n43_adj_4609));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n45_adj_4610), .I1(n13), .I2(n19), .I3(n21), 
            .O(n49_adj_4611));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4611), .I1(n54), .I2(n43_adj_4609), 
            .I3(n44), .O(n23810));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[3]), .I1(n23810), .I2(GND_net), .I3(GND_net), 
            .O(n24143));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mod_5_add_1607_15 (.CI(n23566), .I0(n2297), .I1(n2324), .CO(n23567));
    SB_LUT4 i24780_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30631));
    defparam i24780_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_523[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_c)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1540_18 (.CI(n22620), .I0(n2194), .I1(n2225), .CO(n22621));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n22619), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n22619), .I0(n2195), .I1(n2225), .CO(n22620));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n22618), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n22720), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n22720), .I0(n1803), .I1(n1829), .CO(n22721));
    SB_CARRY mod_5_add_1540_16 (.CI(n22618), .I0(n2196), .I1(n2225), .CO(n22619));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n22617), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n22719), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n22617), .I0(n2197), .I1(n2225), .CO(n22618));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n22616), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n22719), .I0(n1804), .I1(n1829), .CO(n22720));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n22718), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n22718), .I0(n1805), .I1(n1829), .CO(n22719));
    SB_CARRY mod_5_add_1540_14 (.CI(n22616), .I0(n2198), .I1(n2225), .CO(n22617));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n22615), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n22717), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n22717), .I0(n1806), .I1(n1829), .CO(n22718));
    SB_CARRY mod_5_add_1540_13 (.CI(n22615), .I0(n2199), .I1(n2225), .CO(n22616));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n22614), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n22716), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n22716), .I0(n1807), .I1(n1829), .CO(n22717));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n22715), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n22715), .I0(n1808), .I1(n1829), .CO(n22716));
    SB_CARRY mod_5_add_1540_12 (.CI(n22614), .I0(n2200), .I1(n2225), .CO(n22615));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n22613), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n30631), 
            .I3(n22714), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_11 (.CI(n22613), .I0(n2201), .I1(n2225), .CO(n22614));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n22612), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_3 (.CI(n22714), .I0(n1809), .I1(n30631), .CO(n22715));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n30631), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n30631), 
            .CO(n22714));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n22713), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n22712), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n22712), .I0(n1896), .I1(n1928), .CO(n22713));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n22711), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n22711), .I0(n1897), .I1(n1928), .CO(n22712));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n22710), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n22710), .I0(n1898), .I1(n1928), .CO(n22711));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n22709), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n22709), .I0(n1899), .I1(n1928), .CO(n22710));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n22708), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1499 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i1_2_lut_adj_1499.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1540_10 (.CI(n22612), .I0(n2202), .I1(n2225), .CO(n22613));
    SB_CARRY mod_5_add_1339_12 (.CI(n22708), .I0(n1900), .I1(n1928), .CO(n22709));
    SB_LUT4 i14810_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n19377));
    defparam i14810_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n22435));
    SB_LUT4 i13_4_lut (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18), 
            .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n22707), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n22611), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n22611), .I0(n2203), .I1(n2225), .CO(n22612));
    SB_CARRY mod_5_add_1339_11 (.CI(n22707), .I0(n1901), .I1(n1928), .CO(n22708));
    SB_LUT4 i11_4_lut (.I0(n2098), .I1(n19377), .I2(n2094), .I3(n2099), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n22706), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4613));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n22610), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n22706), .I0(n1902), .I1(n1928), .CO(n22707));
    SB_CARRY mod_5_add_1540_8 (.CI(n22610), .I0(n2204), .I1(n2225), .CO(n22611));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n22705), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n22609), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n22705), .I0(n1903), .I1(n1928), .CO(n22706));
    SB_CARRY mod_5_add_1540_7 (.CI(n22609), .I0(n2205), .I1(n2225), .CO(n22610));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n22704), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4614));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1500 (.I0(n27_adj_4614), .I1(n29_adj_4613), .I2(n28), 
            .I3(n30), .O(n2126));
    defparam i16_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n22608), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_6 (.CI(n22608), .I0(n2206), .I1(n2225), .CO(n22609));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n22607), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n22704), .I0(n1904), .I1(n1928), .CO(n22705));
    SB_CARRY mod_5_add_1540_5 (.CI(n22607), .I0(n2207), .I1(n2225), .CO(n22608));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n22703), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n22703), .I0(n1905), .I1(n1928), .CO(n22704));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n22702), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n22702), .I0(n1906), .I1(n1928), .CO(n22703));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n22606), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n22701), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n22701), .I0(n1907), .I1(n1928), .CO(n22702));
    SB_CARRY mod_5_add_1540_4 (.CI(n22606), .I0(n2208), .I1(n2225), .CO(n22607));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n30634), 
            .I3(n22605), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n22700), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_3 (.CI(n22605), .I0(n2209), .I1(n30634), .CO(n22606));
    SB_CARRY mod_5_add_1339_4 (.CI(n22700), .I0(n1908), .I1(n1928), .CO(n22701));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n30635), 
            .I3(n22699), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n30634), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n30634), 
            .CO(n22605));
    SB_CARRY mod_5_add_1339_3 (.CI(n22699), .I0(n1909), .I1(n30635), .CO(n22700));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n30635), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n30635), 
            .CO(n22699));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n22698), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n22697), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4616));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1501 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38));
    defparam i15_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i14772_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n19339));
    defparam i14772_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1502 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n19339), 
            .O(n36));
    defparam i13_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_17 (.CI(n22697), .I0(n1995), .I1(n2027), .CO(n22698));
    SB_LUT4 i19_4_lut_adj_1503 (.I0(n2700), .I1(n38), .I2(n28_adj_4616), 
            .I3(n2705), .O(n42));
    defparam i19_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n22696), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_4_lut_adj_1504 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40));
    defparam i17_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1505 (.I0(n2687), .I1(n36), .I2(n2703), .I3(n2695), 
            .O(n41_adj_4617));
    defparam i18_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1506 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4618));
    defparam i16_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4618), .I1(n41_adj_4617), .I2(n40), 
            .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr__i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n15464), 
            .D(n255[31]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n15464), 
            .D(n255[30]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1406_16 (.CI(n22696), .I0(n1996), .I1(n2027), .CO(n22697));
    SB_DFFESR bit_ctr__i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n15464), 
            .D(n255[29]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i24790_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30641));
    defparam i24790_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n22695), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n23558), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n23559), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n23565), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n23555), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n23558), .I0(n2305), .I1(n2324), .CO(n23559));
    SB_CARRY mod_5_add_1607_8 (.CI(n23559), .I0(n2304), .I1(n2324), .CO(n23560));
    SB_CARRY mod_5_add_1607_14 (.CI(n23565), .I0(n2298), .I1(n2324), .CO(n23566));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n23564), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n22695), .I0(n1997), .I1(n2027), .CO(n22696));
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n22427), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1507 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4621));
    defparam i16_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4622));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1508 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4623));
    defparam i15_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1509 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4624));
    defparam i13_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1510 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4625));
    defparam i18_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1511 (.I0(n37_adj_4624), .I1(n39_adj_4623), .I2(n38_adj_4622), 
            .I3(n40_adj_4621), .O(n46_adj_4626));
    defparam i22_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n22694), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n22694), .I0(n1998), .I1(n2027), .CO(n22695));
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4627));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4627), .I1(n46_adj_4626), .I2(n42_adj_4625), 
            .I3(n34), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24789_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30640));
    defparam i24789_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n22693), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_13 (.CI(n22693), .I0(n1999), .I1(n2027), .CO(n22694));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n22692), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2894), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4629));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1406_12 (.CI(n22692), .I0(n2000), .I1(n2027), .CO(n22693));
    SB_LUT4 i16_4_lut_adj_1512 (.I0(n2885), .I1(n2900), .I2(n2891), .I3(n2889), 
            .O(n41_adj_4630));
    defparam i16_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2895), .I1(n2887), .I2(n2906), .I3(GND_net), 
            .O(n38_adj_4631));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1513 (.I0(n2896), .I1(n2893), .I2(n2890), .I3(n2899), 
            .O(n43_adj_4632));
    defparam i18_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1514 (.I0(n2892), .I1(n2901), .I2(n2902), .I3(n2908), 
            .O(n40_adj_4633));
    defparam i15_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1515 (.I0(n41_adj_4630), .I1(n33_adj_4629), .I2(n2903), 
            .I3(n2886), .O(n46_adj_4634));
    defparam i21_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1516 (.I0(n2907), .I1(n2897), .I2(n2898), .I3(n2904), 
            .O(n39_adj_4635));
    defparam i14_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1517 (.I0(n43_adj_4632), .I1(n2888), .I2(n38_adj_4631), 
            .I3(n2905), .O(n47_adj_4636));
    defparam i22_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_4636), .I1(n39_adj_4635), .I2(n46_adj_4634), 
            .I3(n40_adj_4633), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n22691), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n22691), .I0(n2001), .I1(n2027), .CO(n22692));
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr__i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n15464), 
            .D(n255[28]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i24788_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30639));
    defparam i24788_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1518 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4639));
    defparam i14_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1519 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4640));
    defparam i18_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1520 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4641));
    defparam i16_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1521 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4642));
    defparam i17_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1522 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4643));
    defparam i15_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_4644));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4639), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4645));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut_adj_1523 (.I0(n41_adj_4643), .I1(n43_adj_4642), .I2(n42_adj_4641), 
            .I3(n44_adj_4640), .O(n50));
    defparam i24_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4646));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_4646), .I1(n50), .I2(n46_adj_4645), 
            .I3(n38_adj_4644), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24787_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30638));
    defparam i24787_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24786_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30637));
    defparam i24786_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_3_lut_adj_1524 (.I0(bit_ctr[4]), .I1(n3103), .I2(n3109), 
            .I3(GND_net), .O(n36_adj_4647));
    defparam i9_3_lut_adj_1524.LUT_INIT = 16'hecec;
    SB_LUT4 i19_4_lut_adj_1525 (.I0(n3104), .I1(n3094), .I2(n3095), .I3(n3097), 
            .O(n46_adj_4648));
    defparam i19_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1526 (.I0(n3084), .I1(n3089), .I2(n3083), .I3(n3105), 
            .O(n42_adj_4649));
    defparam i15_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut_adj_1527 (.I0(n3086), .I1(n3091), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_4650));
    defparam i5_2_lut_adj_1527.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1528 (.I0(n3092), .I1(n3098), .I2(n3100), .I3(n3107), 
            .O(n44_adj_4651));
    defparam i17_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1529 (.I0(n3085), .I1(n46_adj_4648), .I2(n36_adj_4647), 
            .I3(n3093), .O(n50_adj_4652));
    defparam i23_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1530 (.I0(n3087), .I1(n42_adj_4649), .I2(n3096), 
            .I3(n3099), .O(n48_adj_4653));
    defparam i21_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1531 (.I0(n3102), .I1(n44_adj_4651), .I2(n32_adj_4650), 
            .I3(n3101), .O(n49_adj_4654));
    defparam i22_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1532 (.I0(n3106), .I1(n3090), .I2(n3108), .I3(n3088), 
            .O(n47_adj_4655));
    defparam i20_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1533 (.I0(n47_adj_4655), .I1(n49_adj_4654), .I2(n48_adj_4653), 
            .I3(n50_adj_4652), .O(n3116));
    defparam i26_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr__i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n15464), 
            .D(n255[27]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n22690), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1534 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4656));
    defparam i14_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n25_adj_4657));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1535 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4658));
    defparam i12_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr__i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n15464), 
            .D(n255[26]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n15464), 
            .D(n255[25]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n22426), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1536 (.I0(n25_adj_4657), .I1(n36_adj_4656), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4659));
    defparam i18_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1537 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4660));
    defparam i16_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4658), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4661));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1538 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4662));
    defparam i15_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1539 (.I0(n37_adj_4662), .I1(n39_adj_4661), .I2(n38_adj_4660), 
            .I3(n40_adj_4659), .O(n2621));
    defparam i21_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i24791_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30642));
    defparam i24791_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24785_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30636));
    defparam i24785_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_10 (.CI(n22690), .I0(n2002), .I1(n2027), .CO(n22691));
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n22689), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n30632), 
            .I3(n23554), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n23554), .I0(n2309), .I1(n30632), .CO(n23555));
    SB_CARRY mod_5_add_1406_9 (.CI(n22689), .I0(n2003), .I1(n2027), .CO(n22690));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n22688), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n22426), .I0(n2391), .I1(n2423), .CO(n22427));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n22425), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr__i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n15464), .D(n255[4]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n30632), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_20 (.CI(n22425), .I0(n2392), .I1(n2423), .CO(n22426));
    SB_DFFESR bit_ctr__i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n15464), .D(n255[3]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n22424), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n22424), .I0(n2393), .I1(n2423), .CO(n22425));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n22423), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n22688), .I0(n2004), .I1(n2027), .CO(n22689));
    SB_CARRY mod_5_add_1674_18 (.CI(n22423), .I0(n2394), .I1(n2423), .CO(n22424));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n22687), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n22298), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n22422), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n22290), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_13 (.CI(n22298), .I0(bit_ctr[11]), .I1(GND_net), .CO(n22299));
    SB_CARRY mod_5_add_1674_17 (.CI(n22422), .I0(n2395), .I1(n2423), .CO(n22423));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n22421), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n22297), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n22421), .I0(n2396), .I1(n2423), .CO(n22422));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n22420), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n22420), .I0(n2397), .I1(n2423), .CO(n22421));
    SB_CARRY add_21_12 (.CI(n22297), .I0(bit_ctr[10]), .I1(GND_net), .CO(n22298));
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n30632), 
            .CO(n23554));
    SB_CARRY mod_5_add_1607_6 (.CI(n23557), .I0(n2306), .I1(n2324), .CO(n23558));
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n22318), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n22317), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_32 (.CI(n22317), .I0(bit_ctr[30]), .I1(GND_net), .CO(n22318));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n22316), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_31 (.CI(n22316), .I0(bit_ctr[29]), .I1(GND_net), .CO(n22317));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n22419), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr__i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n15464), 
            .D(n255[24]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_5 (.CI(n22290), .I0(bit_ctr[3]), .I1(GND_net), .CO(n22291));
    SB_CARRY mod_5_add_1674_14 (.CI(n22419), .I0(n2398), .I1(n2423), .CO(n22420));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n22418), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n22296), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n22315), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr__i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n15464), 
            .D(n255[23]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n22289), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_13 (.CI(n22418), .I0(n2399), .I1(n2423), .CO(n22419));
    SB_CARRY add_21_11 (.CI(n22296), .I0(bit_ctr[9]), .I1(GND_net), .CO(n22297));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_30 (.CI(n22315), .I0(bit_ctr[28]), .I1(GND_net), .CO(n22316));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n22314), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n22314), .I0(bit_ctr[27]), .I1(GND_net), .CO(n22315));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n22417), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n22313), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_7 (.CI(n22687), .I0(n2005), .I1(n2027), .CO(n22688));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n22686), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n22417), .I0(n2400), .I1(n2423), .CO(n22418));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n22416), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_28 (.CI(n22313), .I0(bit_ctr[26]), .I1(GND_net), .CO(n22314));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n22312), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_11 (.CI(n22416), .I0(n2401), .I1(n2423), .CO(n22417));
    SB_DFFESR bit_ctr__i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n15464), 
            .D(n255[22]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_27 (.CI(n22312), .I0(bit_ctr[25]), .I1(GND_net), .CO(n22313));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n22311), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_26 (.CI(n22311), .I0(bit_ctr[24]), .I1(GND_net), .CO(n22312));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n22415), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n22686), .I0(n2006), .I1(n2027), .CO(n22687));
    SB_CARRY mod_5_add_1674_10 (.CI(n22415), .I0(n2402), .I1(n2423), .CO(n22416));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_523[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n22465), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n22414), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n22685), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n23564), .I0(n2299), .I1(n2324), .CO(n23565));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n22295), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n22310), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n22414), .I0(n2403), .I1(n2423), .CO(n22415));
    SB_CARRY add_21_4 (.CI(n22289), .I0(bit_ctr[2]), .I1(GND_net), .CO(n22290));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n23563), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n23563), .I0(n2300), .I1(n2324), .CO(n23564));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n23562), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_523[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n22464), .O(n23_adj_4664)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n22464), .I0(timer[30]), .I1(n1[30]), 
            .CO(n22465));
    SB_CARRY mod_5_add_1406_5 (.CI(n22685), .I0(n2007), .I1(n2027), .CO(n22686));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n22684), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n22684), .I0(n2008), .I1(n2027), .CO(n22685));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_523[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n22463), .O(n28_adj_4665)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n22413), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n30636), 
            .I3(n22683), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_11 (.CI(n23562), .I0(n2301), .I1(n2324), .CO(n23563));
    SB_CARRY mod_5_add_1406_3 (.CI(n22683), .I0(n2009), .I1(n30636), .CO(n22684));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n23561), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n30636), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_8 (.CI(n22413), .I0(n2404), .I1(n2423), .CO(n22414));
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n30636), 
            .CO(n22683));
    SB_CARRY sub_14_add_2_31 (.CI(n22463), .I0(timer[29]), .I1(n1[29]), 
            .CO(n22464));
    SB_CARRY mod_5_add_1607_10 (.CI(n23561), .I0(n2302), .I1(n2324), .CO(n23562));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n22412), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_523[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n22462), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1674_7 (.CI(n22412), .I0(n2405), .I1(n2423), .CO(n22413));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n22411), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_30 (.CI(n22462), .I0(timer[28]), .I1(n1[28]), 
            .CO(n22463));
    SB_CARRY mod_5_add_1674_6 (.CI(n22411), .I0(n2406), .I1(n2423), .CO(n22412));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_523[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n22461), .O(n21_adj_4666)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_10 (.CI(n22295), .I0(bit_ctr[8]), .I1(GND_net), .CO(n22296));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n22294), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n22410), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n22310), .I0(bit_ctr[23]), .I1(GND_net), .CO(n22311));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n22309), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_24 (.CI(n22309), .I0(bit_ctr[22]), .I1(GND_net), .CO(n22310));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n23572), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n22410), .I0(n2407), .I1(n2423), .CO(n22411));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n22308), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24781_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30632));
    defparam i24781_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n23067), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n23066), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n23066), .I0(n3084), .I1(n3116), .CO(n23067));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n23065), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n23065), .I0(n3085), .I1(n3116), .CO(n23066));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n23064), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n22409), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n22409), .I0(n2408), .I1(n2423), .CO(n22410));
    SB_CARRY mod_5_add_2143_26 (.CI(n23064), .I0(n3086), .I1(n3116), .CO(n23065));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n23063), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_29 (.CI(n22461), .I0(timer[27]), .I1(n1[27]), 
            .CO(n22462));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n22460), .O(one_wire_N_523[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n22288), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_25 (.CI(n23063), .I0(n3087), .I1(n3116), .CO(n23064));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n23062), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n23062), .I0(n3088), .I1(n3116), .CO(n23063));
    SB_CARRY sub_14_add_2_28 (.CI(n22460), .I0(timer[26]), .I1(n1[26]), 
            .CO(n22461));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n23061), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n30637), 
            .I3(n22408), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n22408), .I0(n2409), .I1(n30637), .CO(n22409));
    SB_CARRY mod_5_add_2143_23 (.CI(n23061), .I0(n3089), .I1(n3116), .CO(n23062));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n23060), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n23060), .I0(n3090), .I1(n3116), .CO(n23061));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n23059), .O(n47_adj_4608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n23059), .I0(n3091), .I1(n3116), .CO(n23060));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n23058), .O(n45_adj_4610)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n23058), .I0(n3092), .I1(n3116), .CO(n23059));
    SB_CARRY add_21_23 (.CI(n22308), .I0(bit_ctr[21]), .I1(GND_net), .CO(n22309));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n23057), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n23057), .I0(n3093), .I1(n3116), .CO(n23058));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n23056), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n23056), .I0(n3094), .I1(n3116), .CO(n23057));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n23055), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr__i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n15464), .D(n255[0]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n30637), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_17 (.CI(n23055), .I0(n3095), .I1(n3116), .CO(n23056));
    SB_CARRY add_21_9 (.CI(n22294), .I0(bit_ctr[7]), .I1(GND_net), .CO(n22295));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n23054), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n23054), .I0(n3096), .I1(n3116), .CO(n23055));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n23053), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n23053), .I0(n3097), .I1(n3116), .CO(n23054));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n23052), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n23052), .I0(n3098), .I1(n3116), .CO(n23053));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n23051), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n23051), .I0(n3099), .I1(n3116), .CO(n23052));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n23050), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n22459), .O(one_wire_N_523[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n30637), 
            .CO(n22408));
    SB_CARRY mod_5_add_2143_12 (.CI(n23050), .I0(n3100), .I1(n3116), .CO(n23051));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n23049), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n22307), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_22 (.CI(n22307), .I0(bit_ctr[20]), .I1(GND_net), .CO(n22308));
    SB_CARRY mod_5_add_2143_11 (.CI(n23049), .I0(n3101), .I1(n3116), .CO(n23050));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n23048), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n23048), .I0(n3102), .I1(n3116), .CO(n23049));
    SB_DFFESR bit_ctr__i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n15464), 
            .D(n255[21]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n23047), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n22306), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_21 (.CI(n22306), .I0(bit_ctr[19]), .I1(GND_net), .CO(n22307));
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n22305), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_9 (.CI(n23047), .I0(n3103), .I1(n3116), .CO(n23048));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n23046), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n23571), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n23560), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n22293), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_27 (.CI(n22459), .I0(timer[25]), .I1(n1[25]), 
            .CO(n22460));
    SB_CARRY mod_5_add_2143_8 (.CI(n23046), .I0(n3104), .I1(n3116), .CO(n23047));
    SB_CARRY mod_5_add_1607_9 (.CI(n23560), .I0(n2303), .I1(n2324), .CO(n23561));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n23045), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n23045), .I0(n3105), .I1(n3116), .CO(n23046));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n23044), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n23044), .I0(n3106), .I1(n3116), .CO(n23045));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n23043), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n23043), .I0(n3107), .I1(n3116), .CO(n23044));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n23042), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n22458), .O(one_wire_N_523[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_4 (.CI(n23042), .I0(n3108), .I1(n3116), .CO(n23043));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n30638), 
            .I3(n23041), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n23041), .I0(n3109), .I1(n30638), .CO(n23042));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n30638), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n30638), 
            .CO(n23041));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n23040), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n23039), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n23039), .I0(n2985), .I1(n3017), .CO(n23040));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n23038), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n23038), .I0(n2986), .I1(n3017), .CO(n23039));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n23037), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n23037), .I0(n2987), .I1(n3017), .CO(n23038));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n23036), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n23036), .I0(n2988), .I1(n3017), .CO(n23037));
    SB_CARRY sub_14_add_2_26 (.CI(n22458), .I0(timer[24]), .I1(n1[24]), 
            .CO(n22459));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n23035), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_523[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n22457), .O(n30_adj_4667)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_23 (.CI(n23035), .I0(n2989), .I1(n3017), .CO(n23036));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n23034), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n23034), .I0(n2990), .I1(n3017), .CO(n23035));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n23033), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n23033), .I0(n2991), .I1(n3017), .CO(n23034));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n23032), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n23032), .I0(n2992), .I1(n3017), .CO(n23033));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n23031), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n23031), .I0(n2993), .I1(n3017), .CO(n23032));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n23030), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n23030), .I0(n2994), .I1(n3017), .CO(n23031));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n23029), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n23029), .I0(n2995), .I1(n3017), .CO(n23030));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n23028), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n23028), .I0(n2996), .I1(n3017), .CO(n23029));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n23027), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n23027), .I0(n2997), .I1(n3017), .CO(n23028));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n23026), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n23026), .I0(n2998), .I1(n3017), .CO(n23027));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n23025), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n23025), .I0(n2999), .I1(n3017), .CO(n23026));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n23024), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n23024), .I0(n3000), .I1(n3017), .CO(n23025));
    SB_CARRY sub_14_add_2_25 (.CI(n22457), .I0(timer[23]), .I1(n1[23]), 
            .CO(n22458));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n23023), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_523[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n22456), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_11 (.CI(n23023), .I0(n3001), .I1(n3017), .CO(n23024));
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), .I3(GND_net), 
            .O(n27_adj_4668));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1540 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4669));
    defparam i13_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1541 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4670));
    defparam i12_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1542 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4671));
    defparam i11_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1543 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4672));
    defparam i15_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1544 (.I0(n33_adj_4669), .I1(n27_adj_4668), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4673));
    defparam i17_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1545 (.I0(n37_adj_4673), .I1(n35_adj_4672), .I2(n31_adj_4671), 
            .I3(n32_adj_4670), .O(n2423));
    defparam i19_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr__i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n15464), 
            .D(n255[20]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n23022), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n23022), .I0(n3002), .I1(n3017), .CO(n23023));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n23021), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n23021), .I0(n3003), .I1(n3017), .CO(n23022));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n23020), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_24 (.CI(n22456), .I0(timer[22]), .I1(n1[22]), 
            .CO(n22457));
    SB_CARRY mod_5_add_2076_8 (.CI(n23020), .I0(n3004), .I1(n3017), .CO(n23021));
    SB_CARRY mod_5_add_1607_20 (.CI(n23571), .I0(n2292), .I1(n2324), .CO(n23572));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n23019), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_523[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n22455), .O(n25_adj_4674)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_20 (.CI(n22305), .I0(bit_ctr[18]), .I1(GND_net), .CO(n22306));
    SB_CARRY mod_5_add_2076_7 (.CI(n23019), .I0(n3005), .I1(n3017), .CO(n23020));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n23018), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n23018), .I0(n3006), .I1(n3017), .CO(n23019));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n23017), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n23017), .I0(n3007), .I1(n3017), .CO(n23018));
    SB_DFF timer_1207__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i6_4_lut (.I0(bit_ctr[15]), .I1(bit_ctr[12]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[8]), .O(n14_adj_4675));   // verilog/neopixel.v(18[12:19])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n23016), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n23016), .I0(n3008), .I1(n3017), .CO(n23017));
    SB_LUT4 i5_4_lut (.I0(bit_ctr[23]), .I1(bit_ctr[28]), .I2(bit_ctr[13]), 
            .I3(bit_ctr[29]), .O(n13_adj_4676));   // verilog/neopixel.v(18[12:19])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_23 (.CI(n22455), .I0(timer[21]), .I1(n1[21]), 
            .CO(n22456));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n30639), 
            .I3(n23015), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i2_3_lut (.I0(n13_adj_4676), .I1(bit_ctr[30]), .I2(n14_adj_4675), 
            .I3(GND_net), .O(n22_adj_4677));   // verilog/neopixel.v(18[12:19])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1546 (.I0(bit_ctr[20]), .I1(bit_ctr[5]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[16]), .O(n32_adj_4678));   // verilog/neopixel.v(18[12:19])
    defparam i12_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_523[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n22454), .O(n29_adj_4679)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2076_3 (.CI(n23015), .I0(n3009), .I1(n30639), .CO(n23016));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n30639), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_22 (.CI(n22454), .I0(timer[20]), .I1(n1[20]), 
            .CO(n22455));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n30639), 
            .CO(n23015));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n23014), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n23013), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n22453), .O(one_wire_N_523[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_26 (.CI(n23013), .I0(n2886), .I1(n2918), .CO(n23014));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n23012), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n23012), .I0(n2887), .I1(n2918), .CO(n23013));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n23011), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n23011), .I0(n2888), .I1(n2918), .CO(n23012));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n23010), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n23010), .I0(n2889), .I1(n2918), .CO(n23011));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n23009), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n23009), .I0(n2890), .I1(n2918), .CO(n23010));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n23008), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1547 (.I0(bit_ctr[31]), .I1(n32_adj_4678), .I2(n22_adj_4677), 
            .I3(bit_ctr[10]), .O(n36_adj_4680));   // verilog/neopixel.v(18[12:19])
    defparam i16_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_21 (.CI(n23008), .I0(n2891), .I1(n2918), .CO(n23009));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n23007), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n23007), .I0(n2892), .I1(n2918), .CO(n23008));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n23006), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n23006), .I0(n2893), .I1(n2918), .CO(n23007));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n23005), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n23005), .I0(n2894), .I1(n2918), .CO(n23006));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n23004), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n23004), .I0(n2895), .I1(n2918), .CO(n23005));
    SB_LUT4 i14_4_lut_adj_1548 (.I0(bit_ctr[26]), .I1(bit_ctr[7]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[24]), .O(n34_adj_4681));   // verilog/neopixel.v(18[12:19])
    defparam i14_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n23003), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1549 (.I0(bit_ctr[25]), .I1(bit_ctr[11]), .I2(bit_ctr[22]), 
            .I3(bit_ctr[19]), .O(n35_adj_4682));   // verilog/neopixel.v(18[12:19])
    defparam i15_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_16 (.CI(n23003), .I0(n2896), .I1(n2918), .CO(n23004));
    SB_LUT4 i13_4_lut_adj_1550 (.I0(bit_ctr[17]), .I1(bit_ctr[27]), .I2(bit_ctr[14]), 
            .I3(bit_ctr[6]), .O(n33_adj_4683));   // verilog/neopixel.v(18[12:19])
    defparam i13_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n23002), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n23002), .I0(n2897), .I1(n2918), .CO(n23003));
    SB_LUT4 i19_4_lut_adj_1551 (.I0(n33_adj_4683), .I1(n35_adj_4682), .I2(n34_adj_4681), 
            .I3(n36_adj_4680), .O(n24963));   // verilog/neopixel.v(18[12:19])
    defparam i19_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n23001), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n23001), .I0(n2898), .I1(n2918), .CO(n23002));
    SB_LUT4 i21463_2_lut (.I0(n19291), .I1(one_wire_N_523[4]), .I2(GND_net), 
            .I3(GND_net), .O(n27307));
    defparam i21463_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n23000), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n23000), .I0(n2899), .I1(n2918), .CO(n23001));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n22999), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n22999), .I0(n2900), .I1(n2918), .CO(n23000));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n22998), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n22998), .I0(n2901), .I1(n2918), .CO(n22999));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n22997), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n22997), .I0(n2902), .I1(n2918), .CO(n22998));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n22996), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n22996), .I0(n2903), .I1(n2918), .CO(n22997));
    SB_LUT4 i1_2_lut_adj_1552 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n22995), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n22995), .I0(n2904), .I1(n2918), .CO(n22996));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n22994), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n22994), .I0(n2905), .I1(n2918), .CO(n22995));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n22993), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n22993), .I0(n2906), .I1(n2918), .CO(n22994));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n22992), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut (.I0(n14151), .I1(n19313), .I2(n27307), .I3(\state[0] ), 
            .O(n66));   // verilog/neopixel.v(16[20:25])
    defparam i1_4_lut.LUT_INIT = 16'hfaee;
    SB_CARRY mod_5_add_2009_5 (.CI(n22992), .I0(n2907), .I1(n2918), .CO(n22993));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n22991), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n22991), .I0(n2908), .I1(n2918), .CO(n22992));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n30640), 
            .I3(n22990), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n22990), .I0(n2909), .I1(n30640), .CO(n22991));
    SB_LUT4 i2_3_lut_adj_1553 (.I0(one_wire_N_523[3]), .I1(one_wire_N_523[4]), 
            .I2(one_wire_N_523[2]), .I3(GND_net), .O(n19313));
    defparam i2_3_lut_adj_1553.LUT_INIT = 16'h8080;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n30640), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_523[10]), .I1(one_wire_N_523[8]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4685));   // verilog/neopixel.v(104[14:39])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY sub_14_add_2_21 (.CI(n22453), .I0(timer[19]), .I1(n1[19]), 
            .CO(n22454));
    SB_LUT4 i6_4_lut_adj_1554 (.I0(one_wire_N_523[5]), .I1(one_wire_N_523[11]), 
            .I2(one_wire_N_523[7]), .I3(n14275), .O(n14_adj_4686));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(one_wire_N_523[9]), .I1(n14_adj_4686), .I2(n10_adj_4685), 
            .I3(one_wire_N_523[6]), .O(n14151));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n22452), .O(one_wire_N_523[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n30640), 
            .CO(n22990));
    SB_LUT4 i3_4_lut (.I0(n76), .I1(LED_c), .I2(\state[0] ), .I3(\state[1] ), 
            .O(n4659));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n22989), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n22988), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n22988), .I0(n2787), .I1(n2819), .CO(n22989));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n22987), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n22987), .I0(n2788), .I1(n2819), .CO(n22988));
    SB_CARRY sub_14_add_2_20 (.CI(n22452), .I0(timer[18]), .I1(n1[18]), 
            .CO(n22453));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_523[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n22451), .O(n27_adj_4687)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i11018_2_lut (.I0(n15464), .I1(n4659), .I2(GND_net), .I3(GND_net), 
            .O(n15593));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11018_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n22986), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_19 (.CI(n22451), .I0(timer[17]), .I1(n1[17]), 
            .CO(n22452));
    SB_LUT4 i24210_3_lut (.I0(n14151), .I1(\state[0] ), .I2(n19313), .I3(GND_net), 
            .O(n29835));   // verilog/neopixel.v(16[20:25])
    defparam i24210_3_lut.LUT_INIT = 16'h3232;
    SB_CARRY mod_5_add_1942_23 (.CI(n22986), .I0(n2789), .I1(n2819), .CO(n22987));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n22985), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_4_lut (.I0(n66), .I1(n4), .I2(n29835), .I3(\state[1] ), 
            .O(n28213));   // verilog/neopixel.v(16[20:25])
    defparam i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY mod_5_add_1942_22 (.CI(n22985), .I0(n2790), .I1(n2819), .CO(n22986));
    SB_LUT4 i1_4_lut_adj_1555 (.I0(n28213), .I1(\state[1] ), .I2(n4659), 
            .I3(\state[0] ), .O(n15464));
    defparam i1_4_lut_adj_1555.LUT_INIT = 16'hfa32;
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n22984), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n22984), .I0(n2791), .I1(n2819), .CO(n22985));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n22983), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n22983), .I0(n2792), .I1(n2819), .CO(n22984));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n22982), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n22982), .I0(n2793), .I1(n2819), .CO(n22983));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n22981), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n22981), .I0(n2794), .I1(n2819), .CO(n22982));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n22980), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n22980), .I0(n2795), .I1(n2819), .CO(n22981));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n22979), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n22979), .I0(n2796), .I1(n2819), .CO(n22980));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n22978), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4688));
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1942_15 (.CI(n22978), .I0(n2797), .I1(n2819), .CO(n22979));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n22977), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n22977), .I0(n2798), .I1(n2819), .CO(n22978));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n22976), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n22976), .I0(n2799), .I1(n2819), .CO(n22977));
    SB_LUT4 i3_3_lut_adj_1557 (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), 
            .I3(GND_net), .O(n12_adj_4689));
    defparam i3_3_lut_adj_1557.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n22975), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n22975), .I0(n2800), .I1(n2819), .CO(n22976));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n22974), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1558 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4688), 
            .O(n16_adj_4690));
    defparam i7_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_11 (.CI(n22974), .I0(n2801), .I1(n2819), .CO(n22975));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n22973), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16_adj_4690), .I2(n12_adj_4689), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_10 (.CI(n22973), .I0(n2802), .I1(n2819), .CO(n22974));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n22972), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n22450), .O(one_wire_N_523[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n22450), .I0(timer[16]), .I1(n1[16]), 
            .CO(n22451));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n22449), .O(one_wire_N_523[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_9 (.CI(n22972), .I0(n2803), .I1(n2819), .CO(n22973));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n22971), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n22971), .I0(n2804), .I1(n2819), .CO(n22972));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n22970), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n22970), .I0(n2805), .I1(n2819), .CO(n22971));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n22969), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n22969), .I0(n2806), .I1(n2819), .CO(n22970));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n22968), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n22968), .I0(n2807), .I1(n2819), .CO(n22969));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n22967), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n22967), .I0(n2808), .I1(n2819), .CO(n22968));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n30641), 
            .I3(n22966), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n22966), .I0(n2809), .I1(n30641), .CO(n22967));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n30641), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n30641), 
            .CO(n22966));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n22965), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n22964), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n22964), .I0(n2688), .I1(n2720), .CO(n22965));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n22963), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n22963), .I0(n2689), .I1(n2720), .CO(n22964));
    SB_CARRY sub_14_add_2_17 (.CI(n22449), .I0(timer[15]), .I1(n1[15]), 
            .CO(n22450));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n22448), .O(one_wire_N_523[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i95_4_lut (.I0(n27307), .I1(n19313), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n83));
    defparam i95_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i1_4_lut_adj_1559 (.I0(start), .I1(\state[1] ), .I2(n14151), 
            .I3(n83), .O(n1929));
    defparam i1_4_lut_adj_1559.LUT_INIT = 16'h3332;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n22639), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n22962), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n22962), .I0(n2690), .I1(n2720), .CO(n22963));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n22961), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_16 (.CI(n22448), .I0(timer[14]), .I1(n1[14]), 
            .CO(n22449));
    SB_CARRY mod_5_add_1875_21 (.CI(n22961), .I0(n2691), .I1(n2720), .CO(n22962));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n22960), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n22447), .O(one_wire_N_523[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_20 (.CI(n22960), .I0(n2692), .I1(n2720), .CO(n22961));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n22638), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n22638), .I0(n2094), .I1(n2126), .CO(n22639));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n22959), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1875_19 (.CI(n22959), .I0(n2693), .I1(n2720), .CO(n22960));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n22958), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n22958), .I0(n2694), .I1(n2720), .CO(n22959));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n22637), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n22957), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n22957), .I0(n2695), .I1(n2720), .CO(n22958));
    SB_CARRY mod_5_add_1473_17 (.CI(n22637), .I0(n2095), .I1(n2126), .CO(n22638));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n22956), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n22956), .I0(n2696), .I1(n2720), .CO(n22957));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n22955), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n22955), .I0(n2697), .I1(n2720), .CO(n22956));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n22636), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n22954), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_2_lut_adj_1560 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4692));
    defparam i2_2_lut_adj_1560.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1473_16 (.CI(n22636), .I0(n2096), .I1(n2126), .CO(n22637));
    SB_LUT4 i12_4_lut_adj_1561 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4693));
    defparam i12_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n22635), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n22635), .I0(n2097), .I1(n2126), .CO(n22636));
    SB_CARRY mod_5_add_1875_14 (.CI(n22954), .I0(n2698), .I1(n2720), .CO(n22955));
    SB_LUT4 i10_4_lut_adj_1562 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4694));
    defparam i10_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1563 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4695));
    defparam i11_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(bit_ctr[15]), .I1(n18_adj_4692), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4696));
    defparam i9_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1564 (.I0(n25_adj_4696), .I1(n27_adj_4695), .I2(n26_adj_4694), 
            .I3(n28_adj_4693), .O(n2027));
    defparam i15_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n22634), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_15 (.CI(n22447), .I0(timer[13]), .I1(n1[13]), 
            .CO(n22448));
    SB_DFFESR bit_ctr__i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n15464), 
            .D(n255[19]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n22953), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n22953), .I0(n2699), .I1(n2720), .CO(n22954));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n22952), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n22952), .I0(n2700), .I1(n2720), .CO(n22953));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n22951), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n22634), .I0(n2098), .I1(n2126), .CO(n22635));
    SB_CARRY mod_5_add_1875_11 (.CI(n22951), .I0(n2701), .I1(n2720), .CO(n22952));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n22950), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24784_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30635));
    defparam i24784_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24783_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30634));
    defparam i24783_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut (.I0(n27317), .I1(n12884), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i3_2_lut (.I0(n1908), .I1(n1907), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4699));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1875_10 (.CI(n22950), .I0(n2702), .I1(n2720), .CO(n22951));
    SB_LUT4 i11_4_lut_adj_1565 (.I0(n1895), .I1(n1903), .I2(n1901), .I3(n1896), 
            .O(n26_adj_4700));
    defparam i11_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1566 (.I0(start), .I1(n66), .I2(GND_net), .I3(GND_net), 
            .O(n11_adj_4701));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_adj_1566.LUT_INIT = 16'h4444;
    SB_LUT4 i9_4_lut_adj_1567 (.I0(bit_ctr[16]), .I1(n18_adj_4699), .I2(n1906), 
            .I3(n1909), .O(n24_adj_4702));
    defparam i9_4_lut_adj_1567.LUT_INIT = 16'hfefc;
    SB_LUT4 i14742_3_lut (.I0(one_wire_N_523[9]), .I1(one_wire_N_523[11]), 
            .I2(one_wire_N_523[10]), .I3(GND_net), .O(n19309));
    defparam i14742_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i10_4_lut_adj_1568 (.I0(n1900), .I1(n1905), .I2(n1904), .I3(n1899), 
            .O(n25_adj_4703));
    defparam i10_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i24705_3_lut_4_lut (.I0(n12884), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n27317), .O(n27428));   // verilog/neopixel.v(22[26:36])
    defparam i24705_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i14_4_lut_adj_1569 (.I0(n29787), .I1(n11_adj_4701), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n20768));   // verilog/neopixel.v(16[20:25])
    defparam i14_4_lut_adj_1569.LUT_INIT = 16'h0aca;
    SB_LUT4 i24195_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n19471), .I2(n27462), 
            .I3(bit_ctr[28]), .O(n27317));
    defparam i24195_3_lut_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 i24047_3_lut (.I0(n19323), .I1(\state[0] ), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n29821));
    defparam i24047_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i20_4_lut_adj_1570 (.I0(n11_adj_4701), .I1(n29821), .I2(\state[1] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n15468));
    defparam i20_4_lut_adj_1570.LUT_INIT = 16'hcac0;
    SB_LUT4 i8_3_lut_adj_1571 (.I0(n1902), .I1(n1897), .I2(n1898), .I3(GND_net), 
            .O(n23_adj_4704));
    defparam i8_3_lut_adj_1571.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut_adj_1572 (.I0(n23_adj_4704), .I1(n25_adj_4703), .I2(n24_adj_4702), 
            .I3(n26_adj_4700), .O(n1928));
    defparam i14_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i14750_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n19317));   // verilog/neopixel.v(22[26:36])
    defparam i14750_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i24371_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n23810), .I3(GND_net), 
            .O(color_bit_N_566[4]));
    defparam i24371_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i24366_4_lut (.I0(n30880), .I1(n24143), .I2(n30808), .I3(bit_ctr[2]), 
            .O(n29829));
    defparam i24366_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i24765_4_lut (.I0(n30784), .I1(n76), .I2(n29829), .I3(color_bit_N_566[4]), 
            .O(state_3__N_372[0]));   // verilog/neopixel.v(18[12:19])
    defparam i24765_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n30949));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30949_bdd_4_lut (.I0(n30949), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n29081));
    defparam n30949_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1573 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n78));
    defparam i1_2_lut_adj_1573.LUT_INIT = 16'h2222;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25045 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n30877));
    defparam bit_ctr_0__bdd_4_lut_25045.LUT_INIT = 16'he4aa;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n22949), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i21510_2_lut (.I0(one_wire_N_523[2]), .I1(one_wire_N_523[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27356));
    defparam i21510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14724_2_lut (.I0(n27855), .I1(one_wire_N_523[3]), .I2(GND_net), 
            .I3(GND_net), .O(n19291));
    defparam i14724_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24797_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30648));
    defparam i24797_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1574 (.I0(n21_adj_4666), .I1(n23_adj_4664), .I2(n22), 
            .I3(n24), .O(n36_adj_4705));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1575 (.I0(n25_adj_4674), .I1(n27_adj_4687), .I2(n26), 
            .I3(n28_adj_4665), .O(n37_adj_4706));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 n30877_bdd_4_lut (.I0(n30877), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n30880));
    defparam n30877_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19_4_lut_adj_1576 (.I0(n37_adj_4706), .I1(n29_adj_4679), .I2(n36_adj_4705), 
            .I3(n30_adj_4667), .O(n14275));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_24986 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n30823));
    defparam bit_ctr_0__bdd_4_lut_24986.LUT_INIT = 16'he4aa;
    SB_LUT4 n30823_bdd_4_lut (.I0(n30823), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n29210));
    defparam n30823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_24941 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n30817));
    defparam bit_ctr_0__bdd_4_lut_24941.LUT_INIT = 16'he4aa;
    SB_LUT4 n30817_bdd_4_lut (.I0(n30817), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n29213));
    defparam n30817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_24936 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n30805));
    defparam bit_ctr_0__bdd_4_lut_24936.LUT_INIT = 16'he4aa;
    SB_LUT4 n30805_bdd_4_lut (.I0(n30805), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n30808));
    defparam n30805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_24926 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n30787));
    defparam bit_ctr_0__bdd_4_lut_24926.LUT_INIT = 16'he4aa;
    SB_LUT4 n30787_bdd_4_lut (.I0(n30787), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n30389));
    defparam n30787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n29210), .I2(n29213), 
            .I3(n24143), .O(n30781));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30781_bdd_4_lut (.I0(n30781), .I1(n30389), .I2(n29081), .I3(n24143), 
            .O(n30784));
    defparam n30781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut (.I0(one_wire_N_523[10]), .I1(one_wire_N_523[5]), .I2(start), 
            .I3(GND_net), .O(n14_adj_4707));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1875_9 (.CI(n22949), .I0(n2703), .I1(n2720), .CO(n22950));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n22948), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n22948), .I0(n2704), .I1(n2720), .CO(n22949));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n22947), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n22947), .I0(n2705), .I1(n2720), .CO(n22948));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n22946), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n22946), .I0(n2706), .I1(n2720), .CO(n22947));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n22945), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n22945), .I0(n2707), .I1(n2720), .CO(n22946));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n22944), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n22944), .I0(n2708), .I1(n2720), .CO(n22945));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n30642), 
            .I3(n22943), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n22943), .I0(n2709), .I1(n30642), .CO(n22944));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n30642), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n30642), 
            .CO(n22943));
    SB_LUT4 i6_4_lut_adj_1577 (.I0(one_wire_N_523[11]), .I1(one_wire_N_523[7]), 
            .I2(one_wire_N_523[9]), .I3(one_wire_N_523[8]), .O(n15_adj_4708));
    defparam i6_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n22942), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n22941), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n22941), .I0(n2589), .I1(n2621), .CO(n22942));
    SB_LUT4 i8_4_lut_adj_1578 (.I0(n15_adj_4708), .I1(\state[1] ), .I2(n14_adj_4707), 
            .I3(one_wire_N_523[6]), .O(n27482));
    defparam i8_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n22940), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n22633), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n22940), .I0(n2590), .I1(n2621), .CO(n22941));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n22939), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(one_wire_N_523[4]), .I1(n26579), .I2(n19291), 
            .I3(n27356), .O(n103));
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'h45cd;
    SB_CARRY mod_5_add_1808_21 (.CI(n22939), .I0(n2591), .I1(n2621), .CO(n22940));
    SB_LUT4 i24710_3_lut (.I0(n27482), .I1(n103), .I2(n14275), .I3(GND_net), 
            .O(n28956));
    defparam i24710_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n22938), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mux_642_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_580 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_642_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY mod_5_add_1808_20 (.CI(n22938), .I0(n2592), .I1(n2621), .CO(n22939));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n22937), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n22937), .I0(n2593), .I1(n2621), .CO(n22938));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n22936), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n22936), .I0(n2594), .I1(n2621), .CO(n22937));
    SB_LUT4 i24028_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n19323), 
            .I3(GND_net), .O(n29787));   // verilog/neopixel.v(16[20:25])
    defparam i24028_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i6_4_lut_adj_1580 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4709));
    defparam i6_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr__i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n15464), .D(n255[2]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n15464), .D(n255[1]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n15464), 
            .D(n255[18]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n15464), 
            .D(n255[17]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_3_lut (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), .I3(GND_net), 
            .O(n9_adj_4710));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1581 (.I0(n9_adj_4710), .I1(n14_adj_4709), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24796_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30647));
    defparam i24796_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24792_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30643));
    defparam i24792_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n22935), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n22935), .I0(n2595), .I1(n2621), .CO(n22936));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n22934), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n22934), .I0(n2596), .I1(n2621), .CO(n22935));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n22933), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n22933), .I0(n2597), .I1(n2621), .CO(n22934));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n22932), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n22932), .I0(n2598), .I1(n2621), .CO(n22933));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n22931), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n22931), .I0(n2599), .I1(n2621), .CO(n22932));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n22930), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(n1106), .I1(n1104), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4713));
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1583 (.I0(n1105), .I1(n1103), .I2(n1107), .I3(n1108), 
            .O(n12_adj_4714));
    defparam i5_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1584 (.I0(bit_ctr[24]), .I1(n12_adj_4714), .I2(n8_adj_4713), 
            .I3(n1109), .O(n1136));
    defparam i6_4_lut_adj_1584.LUT_INIT = 16'hfefc;
    SB_LUT4 i24802_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30653));
    defparam i24802_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24795_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30646));
    defparam i24795_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24753_2_lut (.I0(n2_adj_4716), .I1(n971[28]), .I2(GND_net), 
            .I3(GND_net), .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i24753_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24751_2_lut (.I0(n2_adj_4716), .I1(n971[29]), .I2(GND_net), 
            .I3(GND_net), .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i24751_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2_adj_4716), 
            .I3(GND_net), .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_3_lut_adj_1585 (.I0(n15523), .I1(n905), .I2(n27428), .I3(GND_net), 
            .O(n8_adj_4717));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut_adj_1585.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n8_adj_4717), .I2(n906), .I3(n12882), 
            .O(n2_adj_4716));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h040c;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2_adj_4716), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n12882), .I1(n971[27]), .I2(n2_adj_4716), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23225_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n29077));
    defparam i23225_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1586 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4718));
    defparam i2_3_lut_adj_1586.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut_adj_1587 (.I0(n2_adj_4716), .I1(n6_adj_4718), .I2(n1005), 
            .I3(n29077), .O(n1037));
    defparam i3_4_lut_adj_1587.LUT_INIT = 16'hfdfc;
    SB_LUT4 i24770_2_lut (.I0(n2_adj_4716), .I1(n971[31]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4719));   // verilog/neopixel.v(22[26:36])
    defparam i24770_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1588 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n12882));
    defparam i1_2_lut_adj_1588.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n24963), 
            .I3(GND_net), .O(n76));   // verilog/neopixel.v(18[12:19])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i14719_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i14719_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1589 (.I0(n708), .I1(n19317), .I2(n27340), .I3(n608), 
            .O(n27462));
    defparam i2_4_lut_adj_1589.LUT_INIT = 16'hfefa;
    SB_LUT4 i24278_3_lut_4_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n24963), 
            .I3(\state[0] ), .O(n29790));   // verilog/neopixel.v(18[12:19])
    defparam i24278_3_lut_4_lut.LUT_INIT = 16'h0700;
    SB_LUT4 i1_2_lut_adj_1590 (.I0(bit_ctr[28]), .I1(n27462), .I2(GND_net), 
            .I3(GND_net), .O(n12884));
    defparam i1_2_lut_adj_1590.LUT_INIT = 16'h9999;
    SB_LUT4 i23152_3_lut (.I0(n27462), .I1(n708), .I2(n27340), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i23152_3_lut.LUT_INIT = 16'h8282;
    SB_CARRY mod_5_add_1808_12 (.CI(n22930), .I0(n2600), .I1(n2621), .CO(n22931));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n22929), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n22929), .I0(n2601), .I1(n2621), .CO(n22930));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n22928), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n22928), .I0(n2602), .I1(n2621), .CO(n22929));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n22927), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n22927), .I0(n2603), .I1(n2621), .CO(n22928));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n22926), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n22926), .I0(n2604), .I1(n2621), .CO(n22927));
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n22925), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n22925), .I0(n2605), .I1(n2621), .CO(n22926));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n22924), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n22924), .I0(n2606), .I1(n2621), .CO(n22925));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n22923), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n22923), .I0(n2607), .I1(n2621), .CO(n22924));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n22304), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24794_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30645));
    defparam i24794_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n22446), .O(one_wire_N_523[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n22922), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n22922), .I0(n2608), .I1(n2621), .CO(n22923));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n30644), 
            .I3(n22921), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n22921), .I0(n2609), .I1(n30644), .CO(n22922));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n30644), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n30644), 
            .CO(n22921));
    SB_CARRY mod_5_add_1473_13 (.CI(n22633), .I0(n2099), .I1(n2126), .CO(n22634));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n22920), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n22919), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n22919), .I0(n2490), .I1(n2522), .CO(n22920));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n22918), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n22632), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n22632), .I0(n2100), .I1(n2126), .CO(n22633));
    SB_CARRY mod_5_add_1741_21 (.CI(n22918), .I0(n2491), .I1(n2522), .CO(n22919));
    SB_LUT4 i3_2_lut_adj_1591 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4724));
    defparam i3_2_lut_adj_1591.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1592 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4725));
    defparam i13_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1593 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4726));
    defparam i1_3_lut_adj_1593.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1594 (.I0(n2490), .I1(n34_adj_4725), .I2(n24_adj_4724), 
            .I3(n2494), .O(n38_adj_4727));
    defparam i17_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1595 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4728));
    defparam i15_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1596 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4726), 
            .O(n37_adj_4729));
    defparam i16_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n22917), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1597 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4730));
    defparam i14_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1598 (.I0(n35_adj_4730), .I1(n37_adj_4729), .I2(n36_adj_4728), 
            .I3(n38_adj_4727), .O(n2522));
    defparam i20_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_20 (.CI(n22917), .I0(n2492), .I1(n2522), .CO(n22918));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n22916), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n22916), .I0(n2493), .I1(n2522), .CO(n22917));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n22915), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n22915), .I0(n2494), .I1(n2522), .CO(n22916));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n22914), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n22914), .I0(n2495), .I1(n2522), .CO(n22915));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n22913), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n22631), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n22913), .I0(n2496), .I1(n2522), .CO(n22914));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n22912), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n22912), .I0(n2497), .I1(n2522), .CO(n22913));
    SB_LUT4 i4_3_lut (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), .I3(GND_net), 
            .O(n17_adj_4731));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n22911), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n22631), .I0(n2101), .I1(n2126), .CO(n22632));
    SB_CARRY add_21_19 (.CI(n22304), .I0(bit_ctr[17]), .I1(GND_net), .CO(n22305));
    SB_CARRY mod_5_add_1741_14 (.CI(n22911), .I0(n2498), .I1(n2522), .CO(n22912));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n22910), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n22910), .I0(n2499), .I1(n2522), .CO(n22911));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n22303), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n22909), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24793_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30644));
    defparam i24793_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1599 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4732));
    defparam i8_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut_adj_1600 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4733));
    defparam i7_3_lut_adj_1600.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1601 (.I0(n21_adj_4732), .I1(n17_adj_4731), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4734));
    defparam i11_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_12 (.CI(n22909), .I0(n2500), .I1(n2522), .CO(n22910));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n22908), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut_adj_1602 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4735));
    defparam i3_2_lut_adj_1602.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1603 (.I0(n1700), .I1(n24_adj_4734), .I2(n20_adj_4733), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_11 (.CI(n22908), .I0(n2501), .I1(n2522), .CO(n22909));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n22907), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n22907), .I0(n2502), .I1(n2522), .CO(n22908));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n22906), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24801_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30652));
    defparam i24801_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_9 (.CI(n22906), .I0(n2503), .I1(n2522), .CO(n22907));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n22905), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n22905), .I0(n2504), .I1(n2522), .CO(n22906));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n22904), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n22904), .I0(n2505), .I1(n2522), .CO(n22905));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n22903), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n22903), .I0(n2506), .I1(n2522), .CO(n22904));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n22902), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr__i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n15464), 
            .D(n255[16]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n22630), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n22902), .I0(n2507), .I1(n2522), .CO(n22903));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n22901), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n22630), .I0(n2102), .I1(n2126), .CO(n22631));
    SB_CARRY mod_5_add_1741_4 (.CI(n22901), .I0(n2508), .I1(n2522), .CO(n22902));
    SB_CARRY add_21_8 (.CI(n22293), .I0(bit_ctr[6]), .I1(GND_net), .CO(n22294));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n30645), 
            .I3(n22900), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i11_4_lut_adj_1604 (.I0(bit_ctr[12]), .I1(n22_adj_4735), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4736));
    defparam i11_4_lut_adj_1604.LUT_INIT = 16'hfefc;
    SB_LUT4 i21639_2_lut_3_lut (.I0(n27482), .I1(one_wire_N_523[4]), .I2(n27356), 
            .I3(GND_net), .O(n27488));
    defparam i21639_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[1] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(GND_net), .O(n4_adj_4737));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h3b3b;
    SB_LUT4 i15_4_lut_adj_1605 (.I0(n2294), .I1(n30_adj_4736), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4738));
    defparam i15_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_3 (.CI(n22900), .I0(n2509), .I1(n30645), .CO(n22901));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n30645), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n30645), 
            .CO(n22900));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n22899), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n22898), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n22898), .I0(n906), .I1(VCC_net), .CO(n22899));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n27428), .I2(VCC_net), 
            .I3(n22897), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n22897), .I0(n27428), .I1(VCC_net), 
            .CO(n22898));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n15523), .I2(VCC_net), 
            .I3(n22896), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n22896), .I0(n15523), .I1(VCC_net), 
            .CO(n22897));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n22629), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n12882), .I2(GND_net), 
            .I3(n22895), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n22446), .I0(timer[12]), .I1(n1[12]), 
            .CO(n22447));
    SB_CARRY mod_5_add_669_3 (.CI(n22895), .I0(n12882), .I1(GND_net), 
            .CO(n22896));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n22445), .O(one_wire_N_523[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n22445), .I0(timer[11]), .I1(n1[11]), 
            .CO(n22446));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n22444), .O(one_wire_N_523[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_9 (.CI(n22629), .I0(n2103), .I1(n2126), .CO(n22630));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n22628), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n22628), .I0(n2104), .I1(n2126), .CO(n22629));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n22627), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_12 (.CI(n22444), .I0(timer[10]), .I1(n1[10]), 
            .CO(n22445));
    SB_CARRY mod_5_add_1473_7 (.CI(n22627), .I0(n2105), .I1(n2126), .CO(n22628));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n22895));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4719), .I1(n4_adj_4719), .I2(n1037), 
            .I3(n22894), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n22893), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n22893), .I0(n1005), .I1(n1037), .CO(n22894));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n22892), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n22892), .I0(n1006), .I1(n1037), .CO(n22893));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n22891), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n22891), .I0(n1007), .I1(n1037), .CO(n22892));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n22890), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n22292), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_736_4 (.CI(n22890), .I0(n1008), .I1(n1037), .CO(n22891));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n30646), 
            .I3(n22889), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n22889), .I0(n1009), .I1(n30646), .CO(n22890));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n30646), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n30646), 
            .CO(n22889));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n22888), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n22887), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n22887), .I0(n1104), .I1(n1136), .CO(n22888));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n22886), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n22886), .I0(n1105), .I1(n1136), .CO(n22887));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n22885), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n22885), .I0(n1106), .I1(n1136), .CO(n22886));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n22884), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n22884), .I0(n1107), .I1(n1136), .CO(n22885));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n22626), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n22883), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n22443), .O(one_wire_N_523[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_4 (.CI(n22883), .I0(n1108), .I1(n1136), .CO(n22884));
    SB_CARRY sub_14_add_2_11 (.CI(n22443), .I0(timer[9]), .I1(n1[9]), 
            .CO(n22444));
    SB_LUT4 i14902_2_lut_3_lut (.I0(n19317), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n19471));   // verilog/neopixel.v(22[26:36])
    defparam i14902_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n30647), 
            .I3(n22882), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n22442), .O(one_wire_N_523[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_3 (.CI(n22882), .I0(n1109), .I1(n30647), .CO(n22883));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n30647), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n30647), 
            .CO(n22882));
    SB_LUT4 i24281_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n27462), .I2(bit_ctr[27]), 
            .I3(n838), .O(n15523));
    defparam i24281_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n22881), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n22880), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n22880), .I0(n1203), .I1(n1235), .CO(n22881));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n22879), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n22879), .I0(n1204), .I1(n1235), .CO(n22880));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n22878), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n22878), .I0(n1205), .I1(n1235), .CO(n22879));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n22877), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n19323), 
            .I3(\neo_pixel_transmitter.done ), .O(n28974));   // verilog/neopixel.v(16[20:25])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY mod_5_add_870_6 (.CI(n22877), .I0(n1206), .I1(n1235), .CO(n22878));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n22876), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n22876), .I0(n1207), .I1(n1235), .CO(n22877));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n22875), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_10 (.CI(n22442), .I0(timer[8]), .I1(n1[8]), 
            .CO(n22443));
    SB_CARRY mod_5_add_870_4 (.CI(n22875), .I0(n1208), .I1(n1235), .CO(n22876));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n30648), 
            .I3(n22874), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n22874), .I0(n1209), .I1(n30648), .CO(n22875));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n30648), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n30648), 
            .CO(n22874));
    SB_LUT4 i13_4_lut_adj_1606 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4739));
    defparam i13_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr__i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n15464), 
            .D(n255[15]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n15464), 
            .D(n255[14]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i14_4_lut_adj_1607 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4740));
    defparam i14_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1608 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4741));
    defparam i12_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr__i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n15464), 
            .D(n255[13]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n15468), .D(state_3__N_372[0]), 
            .S(n20768));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n26579));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1609 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4742));
    defparam i8_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1610 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4743));
    defparam i1_3_lut_adj_1610.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4744));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_21_18 (.CI(n22303), .I0(bit_ctr[16]), .I1(GND_net), .CO(n22304));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n22441), .O(one_wire_N_523[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1611 (.I0(n13_adj_4743), .I1(n20_adj_4742), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4745));
    defparam i10_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_9 (.CI(n22441), .I0(timer[7]), .I1(n1[7]), .CO(n22442));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n22440), .O(one_wire_N_523[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21495_2_lut_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n19317), .I2(n608), 
            .I3(bit_ctr[28]), .O(n27340));
    defparam i21495_2_lut_3_lut_4_lut.LUT_INIT = 16'h5600;
    SB_LUT4 i14756_2_lut_4_lut (.I0(one_wire_N_523[9]), .I1(one_wire_N_523[11]), 
            .I2(one_wire_N_523[10]), .I3(n14275), .O(n19323));
    defparam i14756_2_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i11_4_lut_adj_1612 (.I0(n1601), .I1(n22_adj_4745), .I2(n18_adj_4744), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n22302), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2259_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n27462), .I2(bit_ctr[27]), 
            .I3(n27317), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i2259_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_CARRY add_21_3 (.CI(n22288), .I0(bit_ctr[1]), .I1(GND_net), .CO(n22289));
    SB_CARRY add_21_17 (.CI(n22302), .I0(bit_ctr[15]), .I1(GND_net), .CO(n22303));
    SB_CARRY sub_14_add_2_8 (.CI(n22440), .I0(timer[6]), .I1(n1[6]), .CO(n22441));
    SB_LUT4 i26_4_lut_adj_1613 (.I0(n11_adj_4701), .I1(n29790), .I2(\state[1] ), 
            .I3(n4_adj_4737), .O(n12_adj_4746));   // verilog/neopixel.v(16[20:25])
    defparam i26_4_lut_adj_1613.LUT_INIT = 16'h303a;
    SB_LUT4 i18_4_lut_adj_1614 (.I0(n31_adj_4741), .I1(n33_adj_4740), .I2(n32_adj_4739), 
            .I3(n34_adj_4738), .O(n2324));
    defparam i18_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n22439), .O(one_wire_N_523[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr__i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n15464), 
            .D(n255[12]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_7 (.CI(n22439), .I0(timer[5]), .I1(n1[5]), .CO(n22440));
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(n19317), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hd622;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[17]), .I1(n1807), .I2(n1809), .I3(GND_net), 
            .O(n20_adj_4747));
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i9_4_lut_adj_1615 (.I0(n1801), .I1(n1800), .I2(n1803), .I3(n1804), 
            .O(n23_adj_4748));
    defparam i9_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1616 (.I0(n1808), .I1(n1798), .I2(n1799), .I3(n1805), 
            .O(n22_adj_4749));
    defparam i8_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1617 (.I0(n23_adj_4748), .I1(n1806), .I2(n20_adj_4747), 
            .I3(n1797), .O(n26_adj_4750));
    defparam i12_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1618 (.I0(n1796), .I1(n26_adj_4750), .I2(n22_adj_4749), 
            .I3(n1802), .O(n1829));
    defparam i13_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1619 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4751));
    defparam i10_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1620 (.I0(n2203), .I1(n28_adj_4751), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4752));
    defparam i14_4_lut_adj_1620.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1621 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4753));
    defparam i12_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1207_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n22813), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1622 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4754));
    defparam i13_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1207_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n22812), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_32 (.CI(n22812), .I0(GND_net), .I1(timer[30]), 
            .CO(n22813));
    SB_LUT4 i11_4_lut_adj_1623 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4755));
    defparam i11_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1207_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n22811), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut_adj_1624 (.I0(n29_adj_4755), .I1(n31_adj_4754), .I2(n30_adj_4753), 
            .I3(n32_adj_4752), .O(n2225));
    defparam i17_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1207_add_4_31 (.CI(n22811), .I0(GND_net), .I1(timer[29]), 
            .CO(n22812));
    SB_LUT4 timer_1207_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n22810), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_30 (.CI(n22810), .I0(GND_net), .I1(timer[28]), 
            .CO(n22811));
    SB_LUT4 timer_1207_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n22809), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_29 (.CI(n22809), .I0(GND_net), .I1(timer[27]), 
            .CO(n22810));
    SB_LUT4 timer_1207_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n22808), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_28 (.CI(n22808), .I0(GND_net), .I1(timer[26]), 
            .CO(n22809));
    SB_LUT4 timer_1207_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n22807), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_27 (.CI(n22807), .I0(GND_net), .I1(timer[25]), 
            .CO(n22808));
    SB_LUT4 timer_1207_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n22806), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_26 (.CI(n22806), .I0(GND_net), .I1(timer[24]), 
            .CO(n22807));
    SB_LUT4 timer_1207_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n22805), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_25 (.CI(n22805), .I0(GND_net), .I1(timer[23]), 
            .CO(n22806));
    SB_LUT4 timer_1207_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n22804), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_24 (.CI(n22804), .I0(GND_net), .I1(timer[22]), 
            .CO(n22805));
    SB_LUT4 timer_1207_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n22803), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_23 (.CI(n22803), .I0(GND_net), .I1(timer[21]), 
            .CO(n22804));
    SB_LUT4 timer_1207_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n22802), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_22 (.CI(n22802), .I0(GND_net), .I1(timer[20]), 
            .CO(n22803));
    SB_LUT4 timer_1207_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n22801), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_21 (.CI(n22801), .I0(GND_net), .I1(timer[19]), 
            .CO(n22802));
    SB_LUT4 timer_1207_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n22800), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_20 (.CI(n22800), .I0(GND_net), .I1(timer[18]), 
            .CO(n22801));
    SB_LUT4 timer_1207_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n22799), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_19 (.CI(n22799), .I0(GND_net), .I1(timer[17]), 
            .CO(n22800));
    SB_LUT4 timer_1207_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n22798), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_18 (.CI(n22798), .I0(GND_net), .I1(timer[16]), 
            .CO(n22799));
    SB_LUT4 timer_1207_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n22797), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_17 (.CI(n22797), .I0(GND_net), .I1(timer[15]), 
            .CO(n22798));
    SB_LUT4 timer_1207_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n22796), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_16 (.CI(n22796), .I0(GND_net), .I1(timer[14]), 
            .CO(n22797));
    SB_LUT4 timer_1207_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n22795), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_15 (.CI(n22795), .I0(GND_net), .I1(timer[13]), 
            .CO(n22796));
    SB_LUT4 timer_1207_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n22794), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_14 (.CI(n22794), .I0(GND_net), .I1(timer[12]), 
            .CO(n22795));
    SB_LUT4 timer_1207_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n22793), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_13 (.CI(n22793), .I0(GND_net), .I1(timer[11]), 
            .CO(n22794));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n23570), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1207_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n22792), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_12 (.CI(n22792), .I0(GND_net), .I1(timer[10]), 
            .CO(n22793));
    SB_LUT4 timer_1207_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n22791), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_11 (.CI(n22791), .I0(GND_net), .I1(timer[9]), 
            .CO(n22792));
    SB_LUT4 timer_1207_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n22790), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_10 (.CI(n22790), .I0(GND_net), .I1(timer[8]), 
            .CO(n22791));
    SB_LUT4 timer_1207_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n22789), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_9 (.CI(n22789), .I0(GND_net), .I1(timer[7]), 
            .CO(n22790));
    SB_LUT4 timer_1207_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n22788), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_8 (.CI(n22788), .I0(GND_net), .I1(timer[6]), 
            .CO(n22789));
    SB_LUT4 timer_1207_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n22787), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_7 (.CI(n22787), .I0(GND_net), .I1(timer[5]), 
            .CO(n22788));
    SB_LUT4 timer_1207_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n22786), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_6 (.CI(n22786), .I0(GND_net), .I1(timer[4]), 
            .CO(n22787));
    SB_LUT4 timer_1207_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n22785), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_5 (.CI(n22785), .I0(GND_net), .I1(timer[3]), 
            .CO(n22786));
    SB_LUT4 timer_1207_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n22784), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_4 (.CI(n22784), .I0(GND_net), .I1(timer[2]), 
            .CO(n22785));
    SB_LUT4 timer_1207_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n22783), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_3 (.CI(n22783), .I0(GND_net), .I1(timer[1]), 
            .CO(n22784));
    SB_LUT4 timer_1207_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1207_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1207_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n22783));
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n16226));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n16225));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n16224));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n16223));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n16222));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n16221));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n22782), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n16220));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n22781), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n16219));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n16218));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n16217));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n16216));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n16215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n16214));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i24800_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30651));
    defparam i24800_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1625 (.I0(n1500), .I1(n1506), .I2(n1499), .I3(n1501), 
            .O(n18_adj_4756));
    defparam i7_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1626 (.I0(n1508), .I1(n18_adj_4756), .I2(n1504), 
            .I3(n1502), .O(n20_adj_4757));
    defparam i9_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1627 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4758));
    defparam i4_3_lut_adj_1627.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_937_10 (.CI(n22781), .I0(n1302), .I1(n1334), .CO(n22782));
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n16213));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n22780), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n16212));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n16211));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n16210));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n16209));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n16208));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i10_4_lut_adj_1628 (.I0(n15_adj_4758), .I1(n20_adj_4757), .I2(n1503), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n16207));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n16206));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i24799_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30650));
    defparam i24799_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n16205));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n16204));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n16203));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n16202));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n16201));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n16200));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n16199));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n16198));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n16197));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n16196));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_937_9 (.CI(n22780), .I0(n1303), .I1(n1334), .CO(n22781));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1629 (.I0(n1407), .I1(n1406), .I2(n1403), .I3(n1404), 
            .O(n16_adj_4760));
    defparam i6_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n25291));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n22779), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n22779), .I0(n1304), .I1(n1334), .CO(n22780));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n22778), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_3_lut_adj_1630 (.I0(n1408), .I1(n16_adj_4760), .I2(n1401), 
            .I3(GND_net), .O(n18_adj_4761));
    defparam i8_3_lut_adj_1630.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut_adj_1631 (.I0(n1402), .I1(bit_ctr[21]), .I2(n1409), 
            .I3(GND_net), .O(n13_adj_4762));
    defparam i3_3_lut_adj_1631.LUT_INIT = 16'heaea;
    SB_LUT4 i9_4_lut_adj_1632 (.I0(n13_adj_4762), .I1(n18_adj_4761), .I2(n1405), 
            .I3(n1400), .O(n1433));
    defparam i9_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i24798_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30649));
    defparam i24798_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21601_2_lut (.I0(one_wire_N_523[4]), .I1(n27356), .I2(GND_net), 
            .I3(GND_net), .O(n27450));
    defparam i21601_2_lut.LUT_INIT = 16'h8888;
    SB_DFF timer_1207__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_937_7 (.CI(n22778), .I0(n1305), .I1(n1334), .CO(n22779));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n22777), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n22777), .I0(n1306), .I1(n1334), .CO(n22778));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n22776), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n22776), .I0(n1307), .I1(n1334), .CO(n22777));
    SB_LUT4 i116_4_lut (.I0(n19309), .I1(n27488), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n91));
    defparam i116_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1633 (.I0(n27482), .I1(n27307), .I2(n27450), 
            .I3(n78), .O(n26470));
    defparam i1_4_lut_adj_1633.LUT_INIT = 16'h1511;
    SB_DFFESR bit_ctr__i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n15464), 
            .D(n255[11]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n15464), 
            .D(n255[10]), .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_4_lut_adj_1634 (.I0(n14275), .I1(\state[0] ), .I2(n26470), 
            .I3(n91), .O(n15422));
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'h5150;
    SB_DFFESR bit_ctr__i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n15464), .D(n255[9]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr__i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n15464), .D(n255[8]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i2_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_586 ));
    defparam i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n15422), .D(\neo_pixel_transmitter.done_N_586 ), 
            .R(n28974));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n22775), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n22775), .I0(n1308), .I1(n1334), .CO(n22776));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n30649), 
            .I3(n22774), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n22774), .I0(n1309), .I1(n30649), .CO(n22775));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n30649), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n30649), 
            .CO(n22774));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n22773), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n22772), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n22772), .I0(n1401), .I1(n1433), .CO(n22773));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n22771), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n22771), .I0(n1402), .I1(n1433), .CO(n22772));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n22770), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n22770), .I0(n1403), .I1(n1433), .CO(n22771));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n22769), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n22769), .I0(n1404), .I1(n1433), .CO(n22770));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n22768), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n22438), .O(one_wire_N_523[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_7 (.CI(n22768), .I0(n1405), .I1(n1433), .CO(n22769));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n22767), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n22767), .I0(n1406), .I1(n1433), .CO(n22768));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n22766), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n22766), .I0(n1407), .I1(n1433), .CO(n22767));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n22765), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n22765), .I0(n1408), .I1(n1433), .CO(n22766));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n30650), 
            .I3(n22764), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n22764), .I0(n1409), .I1(n30650), .CO(n22765));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n30650), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_7 (.CI(n22292), .I0(bit_ctr[5]), .I1(GND_net), .CO(n22293));
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n30650), 
            .CO(n22764));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n22763), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n22291), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n22301), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n22762), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n22762), .I0(n1500), .I1(n1532), .CO(n22763));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n22761), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n22761), .I0(n1501), .I1(n1532), .CO(n22762));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n22760), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n22760), .I0(n1502), .I1(n1532), .CO(n22761));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n22759), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_9 (.CI(n22759), .I0(n1503), .I1(n1532), .CO(n22760));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n22758), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n22758), .I0(n1504), .I1(n1532), .CO(n22759));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n22757), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n22757), .I0(n1505), .I1(n1532), .CO(n22758));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n22756), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n22756), .I0(n1506), .I1(n1532), .CO(n22757));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n22755), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n22755), .I0(n1507), .I1(n1532), .CO(n22756));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n22754), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n22754), .I0(n1508), .I1(n1532), .CO(n22755));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n30651), 
            .I3(n22753), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_19 (.CI(n23570), .I0(n2293), .I1(n2324), .CO(n23571));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n23569), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr__i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n15464), .D(n255[7]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_3 (.CI(n22753), .I0(n1509), .I1(n30651), .CO(n22754));
    SB_DFF timer_1207__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n30651), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n30651), 
            .CO(n22753));
    SB_DFF timer_1207__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1207__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n15701));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n12_adj_4746));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n22752), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n22751), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_16 (.CI(n22301), .I0(bit_ctr[14]), .I1(GND_net), .CO(n22302));
    SB_CARRY mod_5_add_1138_13 (.CI(n22751), .I0(n1599), .I1(n1631), .CO(n22752));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n22750), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n22750), .I0(n1600), .I1(n1631), .CO(n22751));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n22749), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n22300), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n22288));
    SB_CARRY mod_5_add_1138_11 (.CI(n22749), .I0(n1601), .I1(n1631), .CO(n22750));
    SB_CARRY add_21_15 (.CI(n22300), .I0(bit_ctr[13]), .I1(GND_net), .CO(n22301));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n22748), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n22748), .I0(n1602), .I1(n1631), .CO(n22749));
    SB_CARRY sub_14_add_2_6 (.CI(n22438), .I0(timer[4]), .I1(n1[4]), .CO(n22439));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n22747), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n22747), .I0(n1603), .I1(n1631), .CO(n22748));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n22746), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n22746), .I0(n1604), .I1(n1631), .CO(n22747));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n22745), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n22745), .I0(n1605), .I1(n1631), .CO(n22746));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n22299), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n22744), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_14 (.CI(n22299), .I0(bit_ctr[12]), .I1(GND_net), .CO(n22300));
    SB_CARRY add_21_6 (.CI(n22291), .I0(bit_ctr[4]), .I1(GND_net), .CO(n22292));
    SB_CARRY mod_5_add_1138_6 (.CI(n22744), .I0(n1606), .I1(n1631), .CO(n22745));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n22743), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n22743), .I0(n1607), .I1(n1631), .CO(n22744));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n22742), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n22742), .I0(n1608), .I1(n1631), .CO(n22743));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n30652), 
            .I3(n22741), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n22741), .I0(n1609), .I1(n30652), .CO(n22742));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n30652), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n30652), 
            .CO(n22741));
    SB_CARRY mod_5_add_1473_6 (.CI(n22626), .I0(n2106), .I1(n2126), .CO(n22627));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n22740), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n22739), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n22739), .I0(n1698), .I1(n1730), .CO(n22740));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n22738), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n22738), .I0(n1699), .I1(n1730), .CO(n22739));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n22737), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n22737), .I0(n1700), .I1(n1730), .CO(n22738));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n22736), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n22736), .I0(n1701), .I1(n1730), .CO(n22737));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n22735), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n22437), .O(one_wire_N_523[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_10 (.CI(n22735), .I0(n1702), .I1(n1730), .CO(n22736));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n22734), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n22734), .I0(n1703), .I1(n1730), .CO(n22735));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n22625), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n22733), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n22625), .I0(n2107), .I1(n2126), .CO(n22626));
    SB_CARRY sub_14_add_2_5 (.CI(n22437), .I0(timer[3]), .I1(n1[3]), .CO(n22438));
    SB_CARRY mod_5_add_1205_8 (.CI(n22733), .I0(n1704), .I1(n1730), .CO(n22734));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n22732), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n22732), .I0(n1705), .I1(n1730), .CO(n22733));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n22731), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n22731), .I0(n1706), .I1(n1730), .CO(n22732));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n22730), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n22730), .I0(n1707), .I1(n1730), .CO(n22731));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n22624), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n22729), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n22729), .I0(n1708), .I1(n1730), .CO(n22730));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n22436), .O(one_wire_N_523[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n30653), 
            .I3(n22728), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n22728), .I0(n1709), .I1(n30653), .CO(n22729));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n30653), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n30653), 
            .CO(n22728));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n22727), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n22624), .I0(n2108), .I1(n2126), .CO(n22625));
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n22726), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr__i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n15464), .D(n255[6]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1272_15 (.CI(n22726), .I0(n1797), .I1(n1829), .CO(n22727));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n22725), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n22725), .I0(n1798), .I1(n1829), .CO(n22726));
    SB_CARRY mod_5_add_1607_18 (.CI(n23569), .I0(n2294), .I1(n2324), .CO(n23570));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n22724), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n30643), 
            .I3(n22623), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n22623), .I0(n2109), .I1(n30643), .CO(n22624));
    SB_CARRY mod_5_add_1272_13 (.CI(n22724), .I0(n1799), .I1(n1829), .CO(n22725));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n30643), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_4 (.CI(n22436), .I0(timer[2]), .I1(n1[2]), .CO(n22437));
    SB_DFFESR bit_ctr__i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n15464), .D(n255[5]), 
            .R(n15593));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n23568), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n22723), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n23568), .I0(n2295), .I1(n2324), .CO(n23569));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n23567), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n23567), .I0(n2296), .I1(n2324), .CO(n23568));
    SB_CARRY mod_5_add_1272_12 (.CI(n22723), .I0(n1800), .I1(n1829), .CO(n22724));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n22722), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n22722), .I0(n1801), .I1(n1829), .CO(n22723));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n22721), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n30643), 
            .CO(n22623));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_c), .I1(timer[1]), .I2(n1[1]), 
            .I3(n22435), .O(n27855)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[6] , GND_net, \Kp[7] , \Kp[8] , motor_state, 
            IntegralLimit, duty, \Kp[1] , \Kp[0] , \Kp[2] , PWMLimit, 
            \Kp[3] , \Ki[9] , \Ki[10] , \Ki[11] , \Ki[8] , \Kp[9] , 
            \Ki[1] , \Ki[0] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , 
            \Ki[6] , \Ki[7] , \Kp[4] , \Kp[5] , \Kp[10] , \Kp[11] , 
            \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] , setpoint, \Ki[12] , 
            \Ki[15] , \Ki[14] , \Ki[13] , clk32MHz, VCC_net, n25, 
            n30633) /* synthesis syn_module_defined=1 */ ;
    input \Kp[6] ;
    input GND_net;
    input \Kp[7] ;
    input \Kp[8] ;
    input [23:0]motor_state;
    input [23:0]IntegralLimit;
    output [23:0]duty;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input [23:0]PWMLimit;
    input \Kp[3] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[8] ;
    input \Kp[9] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input [23:0]setpoint;
    input \Ki[12] ;
    input \Ki[15] ;
    input \Ki[14] ;
    input \Ki[13] ;
    input clk32MHz;
    input VCC_net;
    input n25;
    output n30633;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(21[23:26])
    
    wire n478, n23338;
    wire [21:0]n7725;
    
    wire n585, n23339;
    wire [47:0]n155;
    
    wire n512, n23337, n53, n122, n23300, n439, n23336;
    wire [7:0]n7673;
    wire [6:0]n7683;
    
    wire n630, n23299, n557, n23298, n366, n23335, n293, n23334, 
        n220, n23333, n147, n23332, n484, n23297;
    wire [19:0]n7772;
    wire [18:0]n7794;
    
    wire n23389, n5, n74, n23390, n1105, n23387, n411, n23296, 
        n23388, n1032, n23386;
    wire [20:0]n7749;
    
    wire n23331, n23330, n959, n23385, n338, n23295, n265, n23294, 
        n192, n23293, n23329, n886, n23384, n23328, n50, n119, 
        n551, n813, n23383, n624, n23327, n23326, n23325, n1099, 
        n23324, n1026, n23323, n953, n23322, n880, n23321, n807, 
        n23320, n734, n23319, n661, n23318, n588, n23317, n515, 
        n23316, n442, n23315, n369, n23314, n296, n23313, n223, 
        n23312, n150, n23311, n8, n77;
    wire [5:0]n7692;
    
    wire n28160, n490, n23310;
    wire [4:0]n7700;
    
    wire n417, n23309, n344, n23308, n271, n23307, n198_adj_4178, 
        n23306, n56, n125;
    wire [8:0]n7662;
    
    wire n700, n23292, n627, n23291, n554, n23290, n481, n23289, 
        n22484;
    wire [23:0]n1;
    
    wire n22485;
    wire [23:0]\PID_CONTROLLER.err_23__N_3556 ;
    
    wire n22483, n408, n23288, n335, n23287, n262, n23286, n22482, 
        n195, n23301, n268, n23302, n341, n23303, n189, n23285, 
        n47, n116;
    wire [9:0]n7650;
    
    wire n770, n23284, n697, n23283, n23282, n23281, n23280, n405, 
        n23279, n332, n23278, n259, n23277, n186, n23276, n44, 
        n113;
    wire [10:0]n7637;
    
    wire n840, n23275, n767, n23274, n694, n23273, n621, n23272, 
        n548, n23271, n475, n23270, n402, n23269, n329, n23268, 
        n256, n23267, n183, n23266, n41, n110;
    wire [11:0]n7623;
    
    wire n910, n23265, n837, n23264, n764, n23263, n691, n23262, 
        n618, n23261, n545, n23260, n472, n23259, n399, n23258, 
        n326, n23257, n253, n23256, n487, n23304, n414, n180, 
        n23255, n38, n107;
    wire [12:0]n7608;
    
    wire n980, n23254;
    wire [23:0]n1_adj_4606;
    
    wire n907, n23253, n834, n23252, n761, n23251, n23305, n560, 
        n688, n23250, n615, n23249, n542, n23248, n469, n23247, 
        n396, n23246, n323, n23245, n250, n23244, n177, n23243, 
        n35, n104;
    wire [13:0]n7592;
    
    wire n1050, n23242, n977, n23241, n904, n23240, n831, n23239, 
        n758, n23238, n685, n23237, n612, n23236, n539, n23235, 
        n466, n23234, n22481;
    wire [23:0]duty_23__N_3655;
    wire [23:0]n2908;
    wire [23:0]n2933;
    
    wire n22535, n22534, n393, n23233, n320, n23232, n247, n23231, 
        n174, n23230, n32, n101;
    wire [14:0]n7575;
    
    wire n1120, n23229, n1047, n23228, n974, n23227, n901, n23226, 
        n828, n23225, n755, n23224, n22533, n22480, n22479, n22532, 
        n22531, n22478, n22530, n22477, n22529, n22476, n22528, 
        n22475, n47_adj_4180;
    wire [23:0]n1_adj_4607;
    
    wire n22604, n682, n23223, n609, n23222, n536, n23221, n463, 
        n23220, n390, n23219, n317, n23218, n244, n23217, n171, 
        n23216, n29, n98;
    wire [15:0]n7557;
    
    wire n23215, n1117, n23214;
    wire [23:0]n257;
    
    wire n22603, n1044, n23213;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n17, n22602, n9_adj_4182, n22601, n11_adj_4184, n22527, 
        n971, n23212, n30048, n30045, n898, n23211, n31459, n30387, 
        n30291, n31441, n30289, n825, n23210, n30287, n31435, 
        n27, n15_adj_4185, n13_adj_4186, n11_adj_4187, n29996, n21_adj_4188, 
        n19, n17_adj_4189, n9_adj_4190, n30002, n43, n16, n29977, 
        n8_adj_4191, n45, n24_adj_4192, n7_adj_4193, n5_adj_4194, 
        n30012, n30263, n752, n23209, n679, n23208, n30259, n25_c, 
        n23_adj_4195, n30490, n31, n29_adj_4196, n30365, n37, n35_adj_4197, 
        n33, n30514, n30293, n31428, n30281, n31423, n12_adj_4198, 
        n30025, n31446, n10_adj_4199, n30, n30437, n30033, n31426, 
        n30381, n31452, n30494, n256_adj_4200, n31417, n30536, n31414, 
        n16_adj_4201, n30014, n24_adj_4202, n6_adj_4203, n30407, n30408, 
        n30016, n8_adj_4204, n31412, n30343, n30200;
    wire [10:0]n7934;
    wire [9:0]n7947;
    
    wire n402_adj_4205, n23512;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3631 ;
    
    wire n3_adj_4206, n4_adj_4207, n30397, n30398, n12_adj_4208, n29990, 
        n10_adj_4209, n30_adj_4210, n606, n23207, n29992, n30504, 
        n30212, n30544, n30545, n39, n30525, n6_adj_4211, n30399, 
        n30400, n29979, n30345, n30210, n41_adj_4212, n29982, n30470, 
        n30218, n30512, n4_adj_4213, n30405, n30406, n30027, n30502, 
        n30202, n30542, n30543, n30527, n30018, n30468, n30208, 
        \PID_CONTROLLER.integral_23__N_3630 , n30510, \PID_CONTROLLER.integral_23__N_3628 , 
        n533, n23206, n460, n23205, n387, n23204, n22526, n694_adj_4214, 
        n314, n23203, n767_adj_4216, n840_adj_4217, n241, n23202, 
        n700_adj_4218, n168, n23201, n26, n95;
    wire [16:0]n7538;
    
    wire n23200, n23199, n1114, n23198, n1041, n23197, n968, n23196, 
        n895, n23195, n822, n23194, n749, n23193, n621_adj_4219, 
        n22474, n22473, n676, n23192, n603, n23191, n530, n23190, 
        n457, n23189, n384, n23188, n311, n23187, n22525, n238, 
        n23186, n165, n23185, n113_adj_4226, n44_adj_4227, n186_adj_4228, 
        n259_adj_4229, n332_adj_4231, n405_adj_4233, n478_adj_4234, 
        n551_adj_4235, n624_adj_4237, n697_adj_4238, n770_adj_4239, 
        n116_adj_4240, n47_adj_4241, n189_adj_4242, n262_adj_4243, n335_adj_4244, 
        n23_adj_4245, n92, n408_adj_4246, n481_adj_4247;
    wire [17:0]n7518;
    
    wire n23184, n554_adj_4252, n627_adj_4253, n119_adj_4254, n50_adj_4255, 
        n77_adj_4263, n8_adj_4264, n150_adj_4265, n223_adj_4266, n296_adj_4267, 
        n369_adj_4268, n442_adj_4269, n515_adj_4270, n588_adj_4271, 
        n661_adj_4272, n734_adj_4273, n807_adj_4274, n880_adj_4275, 
        n953_adj_4276, n1026_adj_4277, n1099_adj_4278, n23183, n74_adj_4281, 
        n5_adj_4282, n147_adj_4283, n220_adj_4284, n293_adj_4285, n366_adj_4286, 
        n439_adj_4287, n512_adj_4288, n585_adj_4289, n658, n23182, 
        n731, n804, n877, n950, n1023, n1111, n23181, n521, 
        n156, n1096, n737, n664, n591, n18939, n265_adj_4297, 
        n80, n11_adj_4298, n153, n226, n299, n372, n445, n518, 
        n591_adj_4299, n664_adj_4300, n737_adj_4301, n810, n883, n956, 
        n1029, n560_adj_4303, n630_adj_4304, n195_adj_4305, n487_adj_4306, 
        n1102, n341_adj_4307, n268_adj_4308, n414_adj_4309, n411_adj_4310, 
        n557_adj_4311, n338_adj_4312, n484_adj_4313, n198_adj_4315, 
        n125_adj_4316, n56_adj_4317, n271_adj_4318, n344_adj_4319, n83, 
        n14_adj_4320, n156_adj_4321, n229, n302, n375, n448, n521_adj_4323, 
        n594, n667, n740, n813_adj_4325, n229_adj_4326, n886_adj_4327, 
        n959_adj_4328, n1032_adj_4329, n1105_adj_4330, n31_adj_4331, 
        n877_adj_4332, n1096_adj_4333, n417_adj_4334, n6_adj_4335;
    wire [3:0]n8004;
    wire [4:0]n7997;
    
    wire n518_adj_4336, n445_adj_4337, n372_adj_4339, n86, n17_adj_4340, 
        n1023_adj_4341, n153_adj_4342, n80_adj_4343, n35_adj_4344, n11_adj_4345, 
        n302_adj_4346, n299_adj_4347, n226_adj_4348, n594_adj_4349, 
        n159, n950_adj_4350, n804_adj_4351, n33_adj_4353, n232, n192_adj_4354, 
        n122_adj_4355, n53_adj_4356, n305, n378, n11_adj_4359, n204;
    wire [1:0]n8015;
    
    wire n131, n62, n13_adj_4360, n1038, n23180, n965, n23179, 
        n4_adj_4361;
    wire [2:0]n8010;
    
    wire n490_adj_4362, n892, n23178, n12_adj_4363, n8_adj_4364, n11_adj_4365, 
        n6_adj_4366, n22260, n18_adj_4367, n13_adj_4368, n4_adj_4369, 
        n28011, n15_adj_4370, n819, n23177, n810_adj_4371, n883_adj_4372, 
        n23382, n740_adj_4373, n956_adj_4374, n451, n731_adj_4375, 
        n746, n23176, n475_adj_4376, n22600, n22524, n673, n23175, 
        n658_adj_4379, n600, n23174, n524, n27_adj_4381, n667_adj_4385, 
        n23381, n527, n23173, n454, n23172, n22472, n381, n23171, 
        n23391, n448_adj_4387, n23378, n308, n23170;
    wire [23:0]duty_23__N_3532;
    
    wire n235, n23169, n162, n23168, n597, n20_adj_4389, n89, 
        n14_adj_4390, n83_adj_4391, n23369, n23370, n22599, n23368, 
        n23374, n670;
    wire [18:0]n7497;
    
    wire n23167, n23166, n23165, n1029_adj_4395, n23366, n23367, 
        n22523, n23373, n23164, n1108, n23163, n743, n375_adj_4397, 
        n1035, n23162, n23379, n22471, n962, n23161, n889, n23160, 
        n816, n23159, n23372, n1102_adj_4399, n23377, n9_adj_4400, 
        n17_adj_4401, n22598, n23158, n19_adj_4402, n22522, n22470, 
        n22597, n23157, n21_adj_4404, n22521, n22469, n23156, n22468, 
        n29928, n22520, n22596, n23155, n23340, n23513, n23514, 
        n23341, n29922, n12_adj_4405, n10_adj_4406, n30_adj_4407, 
        n23154, n23365, n23364, n23363;
    wire [5:0]n7989;
    
    wire n23553, n22595, n22467, n23153, n23371, n23152;
    wire [6:0]n7980;
    wire [7:0]n7970;
    
    wire n23536, n23151, n29938, n30171, n30167, n25_adj_4408, n23_adj_4409, 
        n30458, n22519, n29_adj_4410, n30325, n23342, n23343, n23150, 
        n23380, n23348, n23355, n37_adj_4411, n30506, n23356, n23357, 
        n23376, n23354, n23349, n23350, n23344, n23345, n23351, 
        n43_adj_4412, n16_adj_4413, n23358, n22466, n6_adj_4415, n30446, 
        n23359, n23360, n23352, n30447, n23552;
    wire [19:0]n7475;
    
    wire n23149, n23148, n23147, n23146, n8_adj_4417, n23346, n23145, 
        n23353, n45_adj_4419, n24_adj_4420, n23347, n29838, n23144, 
        n23143, n23142, n29908, n23141, n23375, n23140, n22594, 
        n23139, n23138, n23137, n23136, n23135, n23134, n22518, 
        n23133, n39_adj_4422, n23132, n23131, n41_adj_4423, n45_adj_4424, 
        n37_adj_4425, n43_adj_4426, n29906, n30349, n23_adj_4427, 
        n23551, n25_adj_4428, n23550;
    wire [20:0]n7452;
    
    wire n23130, n23129, n23128, n29_adj_4429, n23127, n23549, n23126, 
        n31_adj_4430, n35_adj_4431, n22593, n23125, n33_adj_4432, 
        n23540, n23541, n23538, n23539, n22517, n23546, n23547, 
        n23544, n23545, n23124, n11_adj_4433, n23543, n23542, n23548, 
        n13_adj_4434, n23123, n15_adj_4435, n23122, n27_adj_4436, 
        n23121, n22592, n23120, n23119, n9_adj_4437, n23118, n23117, 
        n17_adj_4438, n23116, n23115, n23114, n19_adj_4439, n21_adj_4440, 
        n23113, n29965, n30420, n29956, n23112, n23111, n12_adj_4441, 
        n30_adj_4442, n29828, n4_adj_4443, n29975, n30229, n30225, 
        n30484, n30341, n30508, n6_adj_4444, n30462, n30463, n6_adj_4445;
    wire [3:0]n7707;
    
    wire n16_adj_4446, n24_adj_4447, n29942, n8_adj_4448, n29940, 
        n30347;
    wire [0:0]n5869;
    wire [21:0]n7428;
    
    wire n23110, n23537, n23109, n23108, n30414, n4_adj_4449, n30450, 
        n30444, n22591, n22516, n30451, n29952, n22590, n10_adj_4450, 
        n29950, n30518, n30416;
    wire [1:0]n7718;
    
    wire n4_adj_4451;
    wire [2:0]n7713;
    
    wire n30445, n22589, n12_adj_4452, n8_adj_4453, n11_adj_4454, 
        n30554, n6_adj_4455, n22128, n18_adj_4456, n22588, n22587, 
        n22515, n23107, n30555, n23106, n30541, n23105, n29944, 
        n30474, n40, n30476, duty_23__N_3679, n23361, n23362, n22514, 
        n29918, n22586, n23104, n23103, n22585, n23102, n23101, 
        n23100, n23099, n23098, n23097, n23096, n29916, n30520, 
        n23095, n23094, n23093, n23092, n23091, n23090, n23089, 
        n22513, n22584, n23088, n23087, n23086, n23085, n23084, 
        n23083, n22583, n23082, n23081, n23080, n23079, n23078, 
        n30422, n23077, n13_adj_4457, n4_adj_4458, n23076, n23075, 
        n23074, n23073, n23072, n23071, n23070, n23069, n23068, 
        n30556, n22582, n22581, n22580, n22579, n30557, n22578, 
        n22577;
    wire [8:0]n7959;
    
    wire n23534, n23533, n22576, n39_adj_4460, n30539, n41_adj_4461, 
        n29910, n22575, n22574, n22573, n30480, n40_adj_4462, n30482, 
        n23532, n23531, n23530, n23529, n23528, n23527, n23526, 
        n23525, n22572, n23524, n23523, n23522, n22571, n23521, 
        n22570, n23520, n23519, n22569, n974_adj_4463, n1047_adj_4464, 
        n1120_adj_4465, n101_adj_4466, n32_adj_4467, n174_adj_4468, 
        n247_adj_4469, n320_adj_4470, n393_adj_4471, n22568, n466_adj_4472, 
        n22567, n539_adj_4473, n612_adj_4474, n685_adj_4475, n758_adj_4476, 
        n831_adj_4477, n904_adj_4478, n22566, n977_adj_4479, n1050_adj_4480, 
        n22565, n104_adj_4481, n35_adj_4482, n23535, n177_adj_4483, 
        n23518, n250_adj_4484, n23517, n22564, n323_adj_4485, n22563, 
        n23516;
    wire [23:0]n28;
    
    wire n396_adj_4487, n469_adj_4488, n22562, n542_adj_4489, n615_adj_4490, 
        n688_adj_4491, n761_adj_4492, n834_adj_4493, n907_adj_4494, 
        n980_adj_4495, n22561, n22560, n22559, n107_adj_4496, n38_adj_4497, 
        n180_adj_4498, n253_adj_4499, n326_adj_4500, n399_adj_4501, 
        n472_adj_4502, n545_adj_4503, n618_adj_4504, n691_adj_4505, 
        n764_adj_4506, n837_adj_4507, n910_adj_4508, n110_adj_4509, 
        n41_adj_4510, n183_adj_4511, n256_adj_4512, n329_adj_4515, n23515, 
        n548_adj_4518, n86_adj_4520, n17_adj_4521, n159_adj_4522, n232_adj_4523, 
        n22103, n305_adj_4524, n378_adj_4525, n451_adj_4526, n524_adj_4527, 
        n597_adj_4528, n670_adj_4529, n743_adj_4530, n816_adj_4531, 
        n889_adj_4532, n962_adj_4533, n1035_adj_4534, n1108_adj_4535, 
        n89_adj_4536, n20_adj_4537, n162_adj_4538, n235_adj_4539, n308_adj_4540, 
        n381_adj_4541, n22069, n454_adj_4542, n527_adj_4543, n600_adj_4544, 
        n673_adj_4545, n746_adj_4546, n23511, n819_adj_4547, n892_adj_4548, 
        n4_adj_4549, n22026, n23510, n23509;
    wire [11:0]n7920;
    
    wire n23508, n23507, n23506, n23505, n23504, n23503, n23502, 
        n23501, n23500, n23499, n23498, n22846, n22845, n22844, 
        n22843, n22842, n22841, n22840, n22839, n22838, n22837, 
        n22836, n22835, n22834, n22833, n22832, n22831, n22830, 
        n22829, n22828, n22827, n22826, n22825;
    wire [12:0]n7905;
    
    wire n23497, n22824, n23496, n23495, n23494, n23493, n23492, 
        n23491, n23490, n23489, n23488, n23487, n23486;
    wire [13:0]n7889;
    
    wire n23485, n23484, n23483, n23482, n965_adj_4557, n23481, 
        n23480, n23479, n23478, n23477, n23476, n23475, n23474, 
        n23473;
    wire [14:0]n7872;
    
    wire n23472, n23471, n23470, n4_adj_4558, n901_adj_4559, n23469, 
        n828_adj_4560, n23468, n755_adj_4561, n23467, n682_adj_4562, 
        n23466, n609_adj_4563, n23465, n536_adj_4564, n23464, n463_adj_4565, 
        n23463, n390_adj_4566, n23462, n317_adj_4567, n23461, n244_adj_4568, 
        n23460, n171_adj_4569, n23459, n29_adj_4570, n98_adj_4571;
    wire [15:0]n7854;
    
    wire n23458, n1117_adj_4572, n23457, n1044_adj_4573, n23456, n971_adj_4574, 
        n23455, n898_adj_4575, n23454, n825_adj_4576, n23453, n752_adj_4577, 
        n23452, n679_adj_4578, n23451, n606_adj_4579, n23450, n533_adj_4580, 
        n23449, n460_adj_4581, n23448, n387_adj_4582, n23447, n314_adj_4583, 
        n23446, n22158, n241_adj_4584, n23445, n168_adj_4585, n23444, 
        n26_adj_4586, n95_adj_4587;
    wire [16:0]n7835;
    
    wire n23443, n23442, n1114_adj_4588, n23441, n1041_adj_4589, n23440, 
        n968_adj_4590, n23439, n895_adj_4591, n23438, n822_adj_4592, 
        n23437, n749_adj_4593, n23436, n676_adj_4594, n23435, n603_adj_4595, 
        n23434, n530_adj_4596, n23433, n457_adj_4597, n23432, n1038_adj_4598, 
        n384_adj_4599, n23431, n311_adj_4600, n23430, n238_adj_4601, 
        n23429, n165_adj_4602, n23428, n23_adj_4603, n92_adj_4604;
    wire [17:0]n7815;
    
    wire n23427, n23426, n23425, n1111_adj_4605, n23424, n23423, 
        n22235, n23422, n23421, n23420, n23419, n23418, n23417, 
        n23416, n23415, n23414, n23413, n23412, n23411, n23410, 
        n23409, n23408, n23407, n23406, n23405, n23404, n23403, 
        n23402, n23401, n23400, n23399, n23398, n23397, n23396, 
        n23395, n23394, n23393, n23392, n22488, n22487, n22486;
    
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_9 (.CI(n23338), .I0(n7725[6]), .I1(n585), 
            .CO(n23339));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n7725[5]), .I2(n512), 
            .I3(n23337), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3503_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n23300));
    SB_CARRY mult_11_add_1225_8 (.CI(n23337), .I0(n7725[5]), .I1(n512), 
            .CO(n23338));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n7725[4]), .I2(n439), 
            .I3(n23336), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n23336), .I0(n7725[4]), .I1(n439), 
            .CO(n23337));
    SB_LUT4 add_3502_9_lut (.I0(GND_net), .I1(n7683[6]), .I2(n630), .I3(n23299), 
            .O(n7673[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3502_8_lut (.I0(GND_net), .I1(n7683[5]), .I2(n557), .I3(n23298), 
            .O(n7673[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n7725[3]), .I2(n366), 
            .I3(n23335), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n23335), .I0(n7725[3]), .I1(n366), 
            .CO(n23336));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n7725[2]), .I2(n293), 
            .I3(n23334), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n23334), .I0(n7725[2]), .I1(n293), 
            .CO(n23335));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n7725[1]), .I2(n220), 
            .I3(n23333), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n23333), .I0(n7725[1]), .I1(n220), 
            .CO(n23334));
    SB_CARRY add_3502_8 (.CI(n23298), .I0(n7683[5]), .I1(n557), .CO(n23299));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n7725[0]), .I2(n147), 
            .I3(n23332), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n23332), .I0(n7725[0]), .I1(n147), 
            .CO(n23333));
    SB_LUT4 add_3502_7_lut (.I0(GND_net), .I1(n7683[4]), .I2(n484), .I3(n23297), 
            .O(n7673[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3512_18_lut (.I0(GND_net), .I1(n7794[15]), .I2(GND_net), 
            .I3(n23389), .O(n7772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3502_7 (.CI(n23297), .I0(n7683[4]), .I1(n484), .CO(n23298));
    SB_CARRY add_3512_18 (.CI(n23389), .I0(n7794[15]), .I1(GND_net), .CO(n23390));
    SB_LUT4 add_3512_16_lut (.I0(GND_net), .I1(n7794[13]), .I2(n1105), 
            .I3(n23387), .O(n7772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3502_6_lut (.I0(GND_net), .I1(n7683[3]), .I2(n411), .I3(n23296), 
            .O(n7673[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_16 (.CI(n23387), .I0(n7794[13]), .I1(n1105), .CO(n23388));
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n23332));
    SB_LUT4 add_3512_15_lut (.I0(GND_net), .I1(n7794[12]), .I2(n1032), 
            .I3(n23386), .O(n7772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_15 (.CI(n23386), .I0(n7794[12]), .I1(n1032), .CO(n23387));
    SB_LUT4 add_3510_23_lut (.I0(GND_net), .I1(n7749[20]), .I2(GND_net), 
            .I3(n23331), .O(n7725[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3510_22_lut (.I0(GND_net), .I1(n7749[19]), .I2(GND_net), 
            .I3(n23330), .O(n7725[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3502_6 (.CI(n23296), .I0(n7683[3]), .I1(n411), .CO(n23297));
    SB_LUT4 add_3512_14_lut (.I0(GND_net), .I1(n7794[11]), .I2(n959), 
            .I3(n23385), .O(n7772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_22 (.CI(n23330), .I0(n7749[19]), .I1(GND_net), .CO(n23331));
    SB_LUT4 add_3502_5_lut (.I0(GND_net), .I1(n7683[2]), .I2(n338), .I3(n23295), 
            .O(n7673[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3502_5 (.CI(n23295), .I0(n7683[2]), .I1(n338), .CO(n23296));
    SB_LUT4 add_3502_4_lut (.I0(GND_net), .I1(n7683[1]), .I2(n265), .I3(n23294), 
            .O(n7673[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3502_4 (.CI(n23294), .I0(n7683[1]), .I1(n265), .CO(n23295));
    SB_LUT4 add_3502_3_lut (.I0(GND_net), .I1(n7683[0]), .I2(n192), .I3(n23293), 
            .O(n7673[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_14 (.CI(n23385), .I0(n7794[11]), .I1(n959), .CO(n23386));
    SB_LUT4 add_3510_21_lut (.I0(GND_net), .I1(n7749[18]), .I2(GND_net), 
            .I3(n23329), .O(n7725[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3502_3 (.CI(n23293), .I0(n7683[0]), .I1(n192), .CO(n23294));
    SB_LUT4 add_3512_13_lut (.I0(GND_net), .I1(n7794[10]), .I2(n886), 
            .I3(n23384), .O(n7772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_21 (.CI(n23329), .I0(n7749[18]), .I1(GND_net), .CO(n23330));
    SB_CARRY add_3512_13 (.CI(n23384), .I0(n7794[10]), .I1(n886), .CO(n23385));
    SB_LUT4 add_3510_20_lut (.I0(GND_net), .I1(n7749[17]), .I2(GND_net), 
            .I3(n23328), .O(n7725[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3502_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n7673[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3502_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3512_12_lut (.I0(GND_net), .I1(n7794[9]), .I2(n813), .I3(n23383), 
            .O(n7772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3510_20 (.CI(n23328), .I0(n7749[17]), .I1(GND_net), .CO(n23329));
    SB_LUT4 add_3510_19_lut (.I0(GND_net), .I1(n7749[16]), .I2(GND_net), 
            .I3(n23327), .O(n7725[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_19 (.CI(n23327), .I0(n7749[16]), .I1(GND_net), .CO(n23328));
    SB_LUT4 add_3510_18_lut (.I0(GND_net), .I1(n7749[15]), .I2(GND_net), 
            .I3(n23326), .O(n7725[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_18 (.CI(n23326), .I0(n7749[15]), .I1(GND_net), .CO(n23327));
    SB_LUT4 add_3510_17_lut (.I0(GND_net), .I1(n7749[14]), .I2(GND_net), 
            .I3(n23325), .O(n7725[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_17 (.CI(n23325), .I0(n7749[14]), .I1(GND_net), .CO(n23326));
    SB_LUT4 add_3510_16_lut (.I0(GND_net), .I1(n7749[13]), .I2(n1099), 
            .I3(n23324), .O(n7725[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_16 (.CI(n23324), .I0(n7749[13]), .I1(n1099), .CO(n23325));
    SB_LUT4 add_3510_15_lut (.I0(GND_net), .I1(n7749[12]), .I2(n1026), 
            .I3(n23323), .O(n7725[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_15 (.CI(n23323), .I0(n7749[12]), .I1(n1026), .CO(n23324));
    SB_LUT4 add_3510_14_lut (.I0(GND_net), .I1(n7749[11]), .I2(n953), 
            .I3(n23322), .O(n7725[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_14 (.CI(n23322), .I0(n7749[11]), .I1(n953), .CO(n23323));
    SB_LUT4 add_3510_13_lut (.I0(GND_net), .I1(n7749[10]), .I2(n880), 
            .I3(n23321), .O(n7725[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_13 (.CI(n23321), .I0(n7749[10]), .I1(n880), .CO(n23322));
    SB_LUT4 add_3510_12_lut (.I0(GND_net), .I1(n7749[9]), .I2(n807), .I3(n23320), 
            .O(n7725[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_12 (.CI(n23320), .I0(n7749[9]), .I1(n807), .CO(n23321));
    SB_LUT4 add_3510_11_lut (.I0(GND_net), .I1(n7749[8]), .I2(n734), .I3(n23319), 
            .O(n7725[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_11 (.CI(n23319), .I0(n7749[8]), .I1(n734), .CO(n23320));
    SB_LUT4 add_3510_10_lut (.I0(GND_net), .I1(n7749[7]), .I2(n661), .I3(n23318), 
            .O(n7725[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_10 (.CI(n23318), .I0(n7749[7]), .I1(n661), .CO(n23319));
    SB_LUT4 add_3510_9_lut (.I0(GND_net), .I1(n7749[6]), .I2(n588), .I3(n23317), 
            .O(n7725[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_9 (.CI(n23317), .I0(n7749[6]), .I1(n588), .CO(n23318));
    SB_LUT4 add_3510_8_lut (.I0(GND_net), .I1(n7749[5]), .I2(n515), .I3(n23316), 
            .O(n7725[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_8 (.CI(n23316), .I0(n7749[5]), .I1(n515), .CO(n23317));
    SB_LUT4 add_3510_7_lut (.I0(GND_net), .I1(n7749[4]), .I2(n442), .I3(n23315), 
            .O(n7725[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_7 (.CI(n23315), .I0(n7749[4]), .I1(n442), .CO(n23316));
    SB_LUT4 add_3510_6_lut (.I0(GND_net), .I1(n7749[3]), .I2(n369), .I3(n23314), 
            .O(n7725[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_6 (.CI(n23314), .I0(n7749[3]), .I1(n369), .CO(n23315));
    SB_LUT4 add_3510_5_lut (.I0(GND_net), .I1(n7749[2]), .I2(n296), .I3(n23313), 
            .O(n7725[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_5 (.CI(n23313), .I0(n7749[2]), .I1(n296), .CO(n23314));
    SB_LUT4 add_3510_4_lut (.I0(GND_net), .I1(n7749[1]), .I2(n223), .I3(n23312), 
            .O(n7725[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_4 (.CI(n23312), .I0(n7749[1]), .I1(n223), .CO(n23313));
    SB_LUT4 add_3510_3_lut (.I0(GND_net), .I1(n7749[0]), .I2(n150), .I3(n23311), 
            .O(n7725[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_3 (.CI(n23311), .I0(n7749[0]), .I1(n150), .CO(n23312));
    SB_LUT4 add_3510_2_lut (.I0(GND_net), .I1(n8), .I2(n77), .I3(GND_net), 
            .O(n7725[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3510_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3510_2 (.CI(GND_net), .I0(n8), .I1(n77), .CO(n23311));
    SB_LUT4 add_3504_7_lut (.I0(GND_net), .I1(n28160), .I2(n490), .I3(n23310), 
            .O(n7692[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3504_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3504_6_lut (.I0(GND_net), .I1(n7700[3]), .I2(n417), .I3(n23309), 
            .O(n7692[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3504_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3504_6 (.CI(n23309), .I0(n7700[3]), .I1(n417), .CO(n23310));
    SB_LUT4 add_3504_5_lut (.I0(GND_net), .I1(n7700[2]), .I2(n344), .I3(n23308), 
            .O(n7692[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3504_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3504_5 (.CI(n23308), .I0(n7700[2]), .I1(n344), .CO(n23309));
    SB_LUT4 add_3504_4_lut (.I0(GND_net), .I1(n7700[1]), .I2(n271), .I3(n23307), 
            .O(n7692[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3504_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3504_4 (.CI(n23307), .I0(n7700[1]), .I1(n271), .CO(n23308));
    SB_LUT4 add_3504_3_lut (.I0(GND_net), .I1(n7700[0]), .I2(n198_adj_4178), 
            .I3(n23306), .O(n7692[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3504_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3504_3 (.CI(n23306), .I0(n7700[0]), .I1(n198_adj_4178), 
            .CO(n23307));
    SB_LUT4 add_3504_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n7692[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3504_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3503_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n7683[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3502_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n23293));
    SB_LUT4 add_3501_10_lut (.I0(GND_net), .I1(n7673[7]), .I2(n700), .I3(n23292), 
            .O(n7662[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3501_9_lut (.I0(GND_net), .I1(n7673[6]), .I2(n627), .I3(n23291), 
            .O(n7662[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_9 (.CI(n23291), .I0(n7673[6]), .I1(n627), .CO(n23292));
    SB_LUT4 add_3501_8_lut (.I0(GND_net), .I1(n7673[5]), .I2(n554), .I3(n23290), 
            .O(n7662[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_8 (.CI(n23290), .I0(n7673[5]), .I1(n554), .CO(n23291));
    SB_LUT4 add_3501_7_lut (.I0(GND_net), .I1(n7673[4]), .I2(n481), .I3(n23289), 
            .O(n7662[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n22484), .I0(motor_state[19]), 
            .I1(n1[19]), .CO(n22485));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1[18]), .I3(n22483), .O(\PID_CONTROLLER.err_23__N_3556 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n22483), .I0(motor_state[18]), 
            .I1(n1[18]), .CO(n22484));
    SB_CARRY add_3501_7 (.CI(n23289), .I0(n7673[4]), .I1(n481), .CO(n23290));
    SB_LUT4 add_3501_6_lut (.I0(GND_net), .I1(n7673[3]), .I2(n408), .I3(n23288), 
            .O(n7662[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_6 (.CI(n23288), .I0(n7673[3]), .I1(n408), .CO(n23289));
    SB_LUT4 add_3501_5_lut (.I0(GND_net), .I1(n7673[2]), .I2(n335), .I3(n23287), 
            .O(n7662[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_5 (.CI(n23287), .I0(n7673[2]), .I1(n335), .CO(n23288));
    SB_LUT4 add_3501_4_lut (.I0(GND_net), .I1(n7673[1]), .I2(n262), .I3(n23286), 
            .O(n7662[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_4 (.CI(n23286), .I0(n7673[1]), .I1(n262), .CO(n23287));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1[17]), .I3(n22482), .O(\PID_CONTROLLER.err_23__N_3556 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3503_3 (.CI(n23300), .I0(n7692[0]), .I1(n195), .CO(n23301));
    SB_LUT4 add_3503_3_lut (.I0(GND_net), .I1(n7692[0]), .I2(n195), .I3(n23300), 
            .O(n7683[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3503_4 (.CI(n23301), .I0(n7692[1]), .I1(n268), .CO(n23302));
    SB_LUT4 add_3503_4_lut (.I0(GND_net), .I1(n7692[1]), .I2(n268), .I3(n23301), 
            .O(n7683[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3503_5 (.CI(n23302), .I0(n7692[2]), .I1(n341), .CO(n23303));
    SB_LUT4 add_3503_5_lut (.I0(GND_net), .I1(n7692[2]), .I2(n341), .I3(n23302), 
            .O(n7683[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3504_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n23306));
    SB_LUT4 add_3501_3_lut (.I0(GND_net), .I1(n7673[0]), .I2(n189), .I3(n23285), 
            .O(n7662[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_3 (.CI(n23285), .I0(n7673[0]), .I1(n189), .CO(n23286));
    SB_LUT4 add_3501_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n7662[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n23285));
    SB_LUT4 add_3500_11_lut (.I0(GND_net), .I1(n7662[8]), .I2(n770), .I3(n23284), 
            .O(n7650[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3500_10_lut (.I0(GND_net), .I1(n7662[7]), .I2(n697), .I3(n23283), 
            .O(n7650[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_10 (.CI(n23283), .I0(n7662[7]), .I1(n697), .CO(n23284));
    SB_LUT4 add_3500_9_lut (.I0(GND_net), .I1(n7662[6]), .I2(n624), .I3(n23282), 
            .O(n7650[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_9 (.CI(n23282), .I0(n7662[6]), .I1(n624), .CO(n23283));
    SB_LUT4 add_3500_8_lut (.I0(GND_net), .I1(n7662[5]), .I2(n551), .I3(n23281), 
            .O(n7650[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_8 (.CI(n23281), .I0(n7662[5]), .I1(n551), .CO(n23282));
    SB_LUT4 add_3500_7_lut (.I0(GND_net), .I1(n7662[4]), .I2(n478), .I3(n23280), 
            .O(n7650[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_7 (.CI(n23280), .I0(n7662[4]), .I1(n478), .CO(n23281));
    SB_LUT4 add_3500_6_lut (.I0(GND_net), .I1(n7662[3]), .I2(n405), .I3(n23279), 
            .O(n7650[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_6 (.CI(n23279), .I0(n7662[3]), .I1(n405), .CO(n23280));
    SB_LUT4 add_3500_5_lut (.I0(GND_net), .I1(n7662[2]), .I2(n332), .I3(n23278), 
            .O(n7650[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_5 (.CI(n23278), .I0(n7662[2]), .I1(n332), .CO(n23279));
    SB_LUT4 add_3500_4_lut (.I0(GND_net), .I1(n7662[1]), .I2(n259), .I3(n23277), 
            .O(n7650[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_4 (.CI(n23277), .I0(n7662[1]), .I1(n259), .CO(n23278));
    SB_LUT4 add_3500_3_lut (.I0(GND_net), .I1(n7662[0]), .I2(n186), .I3(n23276), 
            .O(n7650[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_3 (.CI(n23276), .I0(n7662[0]), .I1(n186), .CO(n23277));
    SB_LUT4 add_3500_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n7650[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3500_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3500_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n23276));
    SB_LUT4 add_3499_12_lut (.I0(GND_net), .I1(n7650[9]), .I2(n840), .I3(n23275), 
            .O(n7637[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3499_11_lut (.I0(GND_net), .I1(n7650[8]), .I2(n767), .I3(n23274), 
            .O(n7637[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_11 (.CI(n23274), .I0(n7650[8]), .I1(n767), .CO(n23275));
    SB_LUT4 add_3499_10_lut (.I0(GND_net), .I1(n7650[7]), .I2(n694), .I3(n23273), 
            .O(n7637[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_10 (.CI(n23273), .I0(n7650[7]), .I1(n694), .CO(n23274));
    SB_LUT4 add_3499_9_lut (.I0(GND_net), .I1(n7650[6]), .I2(n621), .I3(n23272), 
            .O(n7637[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_9 (.CI(n23272), .I0(n7650[6]), .I1(n621), .CO(n23273));
    SB_LUT4 add_3499_8_lut (.I0(GND_net), .I1(n7650[5]), .I2(n548), .I3(n23271), 
            .O(n7637[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_8 (.CI(n23271), .I0(n7650[5]), .I1(n548), .CO(n23272));
    SB_LUT4 add_3499_7_lut (.I0(GND_net), .I1(n7650[4]), .I2(n475), .I3(n23270), 
            .O(n7637[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_7 (.CI(n23270), .I0(n7650[4]), .I1(n475), .CO(n23271));
    SB_LUT4 add_3499_6_lut (.I0(GND_net), .I1(n7650[3]), .I2(n402), .I3(n23269), 
            .O(n7637[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_6 (.CI(n23269), .I0(n7650[3]), .I1(n402), .CO(n23270));
    SB_LUT4 add_3499_5_lut (.I0(GND_net), .I1(n7650[2]), .I2(n329), .I3(n23268), 
            .O(n7637[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_5 (.CI(n23268), .I0(n7650[2]), .I1(n329), .CO(n23269));
    SB_LUT4 add_3499_4_lut (.I0(GND_net), .I1(n7650[1]), .I2(n256), .I3(n23267), 
            .O(n7637[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_4 (.CI(n23267), .I0(n7650[1]), .I1(n256), .CO(n23268));
    SB_LUT4 add_3499_3_lut (.I0(GND_net), .I1(n7650[0]), .I2(n183), .I3(n23266), 
            .O(n7637[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_3 (.CI(n23266), .I0(n7650[0]), .I1(n183), .CO(n23267));
    SB_LUT4 add_3499_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n7637[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3499_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3499_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n23266));
    SB_LUT4 add_3498_13_lut (.I0(GND_net), .I1(n7637[10]), .I2(n910), 
            .I3(n23265), .O(n7623[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3498_12_lut (.I0(GND_net), .I1(n7637[9]), .I2(n837), .I3(n23264), 
            .O(n7623[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_12 (.CI(n23264), .I0(n7637[9]), .I1(n837), .CO(n23265));
    SB_LUT4 add_3498_11_lut (.I0(GND_net), .I1(n7637[8]), .I2(n764), .I3(n23263), 
            .O(n7623[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_11 (.CI(n23263), .I0(n7637[8]), .I1(n764), .CO(n23264));
    SB_LUT4 add_3498_10_lut (.I0(GND_net), .I1(n7637[7]), .I2(n691), .I3(n23262), 
            .O(n7623[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_10 (.CI(n23262), .I0(n7637[7]), .I1(n691), .CO(n23263));
    SB_LUT4 add_3498_9_lut (.I0(GND_net), .I1(n7637[6]), .I2(n618), .I3(n23261), 
            .O(n7623[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_9 (.CI(n23261), .I0(n7637[6]), .I1(n618), .CO(n23262));
    SB_LUT4 add_3498_8_lut (.I0(GND_net), .I1(n7637[5]), .I2(n545), .I3(n23260), 
            .O(n7623[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_8 (.CI(n23260), .I0(n7637[5]), .I1(n545), .CO(n23261));
    SB_LUT4 add_3498_7_lut (.I0(GND_net), .I1(n7637[4]), .I2(n472), .I3(n23259), 
            .O(n7623[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_7 (.CI(n23259), .I0(n7637[4]), .I1(n472), .CO(n23260));
    SB_LUT4 add_3498_6_lut (.I0(GND_net), .I1(n7637[3]), .I2(n399), .I3(n23258), 
            .O(n7623[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_6 (.CI(n23258), .I0(n7637[3]), .I1(n399), .CO(n23259));
    SB_LUT4 add_3498_5_lut (.I0(GND_net), .I1(n7637[2]), .I2(n326), .I3(n23257), 
            .O(n7623[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_5 (.CI(n23257), .I0(n7637[2]), .I1(n326), .CO(n23258));
    SB_LUT4 add_3498_4_lut (.I0(GND_net), .I1(n7637[1]), .I2(n253), .I3(n23256), 
            .O(n7623[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3503_7_lut (.I0(GND_net), .I1(n7692[4]), .I2(n487), .I3(n23304), 
            .O(n7683[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3503_6 (.CI(n23303), .I0(n7692[3]), .I1(n414), .CO(n23304));
    SB_CARRY add_3498_4 (.CI(n23256), .I0(n7637[1]), .I1(n253), .CO(n23257));
    SB_LUT4 add_3498_3_lut (.I0(GND_net), .I1(n7637[0]), .I2(n180), .I3(n23255), 
            .O(n7623[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_3 (.CI(n23255), .I0(n7637[0]), .I1(n180), .CO(n23256));
    SB_LUT4 add_3498_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n7623[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3498_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3498_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n23255));
    SB_LUT4 add_3497_14_lut (.I0(GND_net), .I1(n7623[11]), .I2(n980), 
            .I3(n23254), .O(n7608[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3497_13_lut (.I0(GND_net), .I1(n7623[10]), .I2(n907), 
            .I3(n23253), .O(n7608[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_13 (.CI(n23253), .I0(n7623[10]), .I1(n907), .CO(n23254));
    SB_LUT4 add_3497_12_lut (.I0(GND_net), .I1(n7623[9]), .I2(n834), .I3(n23252), 
            .O(n7608[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_12 (.CI(n23252), .I0(n7623[9]), .I1(n834), .CO(n23253));
    SB_LUT4 add_3497_11_lut (.I0(GND_net), .I1(n7623[8]), .I2(n761), .I3(n23251), 
            .O(n7608[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_11 (.CI(n23251), .I0(n7623[8]), .I1(n761), .CO(n23252));
    SB_LUT4 add_3503_6_lut (.I0(GND_net), .I1(n7692[3]), .I2(n414), .I3(n23303), 
            .O(n7683[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3503_7 (.CI(n23304), .I0(n7692[4]), .I1(n487), .CO(n23305));
    SB_LUT4 add_3503_8_lut (.I0(GND_net), .I1(n7692[5]), .I2(n560), .I3(n23305), 
            .O(n7683[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3497_10_lut (.I0(GND_net), .I1(n7623[7]), .I2(n688), .I3(n23250), 
            .O(n7608[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_10 (.CI(n23250), .I0(n7623[7]), .I1(n688), .CO(n23251));
    SB_LUT4 add_3497_9_lut (.I0(GND_net), .I1(n7623[6]), .I2(n615), .I3(n23249), 
            .O(n7608[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_9 (.CI(n23249), .I0(n7623[6]), .I1(n615), .CO(n23250));
    SB_LUT4 add_3497_8_lut (.I0(GND_net), .I1(n7623[5]), .I2(n542), .I3(n23248), 
            .O(n7608[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_8 (.CI(n23248), .I0(n7623[5]), .I1(n542), .CO(n23249));
    SB_LUT4 add_3497_7_lut (.I0(GND_net), .I1(n7623[4]), .I2(n469), .I3(n23247), 
            .O(n7608[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_7 (.CI(n23247), .I0(n7623[4]), .I1(n469), .CO(n23248));
    SB_LUT4 add_3497_6_lut (.I0(GND_net), .I1(n7623[3]), .I2(n396), .I3(n23246), 
            .O(n7608[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_6 (.CI(n23246), .I0(n7623[3]), .I1(n396), .CO(n23247));
    SB_LUT4 add_3497_5_lut (.I0(GND_net), .I1(n7623[2]), .I2(n323), .I3(n23245), 
            .O(n7608[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_5 (.CI(n23245), .I0(n7623[2]), .I1(n323), .CO(n23246));
    SB_LUT4 add_3497_4_lut (.I0(GND_net), .I1(n7623[1]), .I2(n250), .I3(n23244), 
            .O(n7608[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_4 (.CI(n23244), .I0(n7623[1]), .I1(n250), .CO(n23245));
    SB_LUT4 add_3497_3_lut (.I0(GND_net), .I1(n7623[0]), .I2(n177), .I3(n23243), 
            .O(n7608[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_3 (.CI(n23243), .I0(n7623[0]), .I1(n177), .CO(n23244));
    SB_LUT4 add_3497_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n7608[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3497_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3497_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n23243));
    SB_LUT4 add_3496_15_lut (.I0(GND_net), .I1(n7608[12]), .I2(n1050), 
            .I3(n23242), .O(n7592[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3496_14_lut (.I0(GND_net), .I1(n7608[11]), .I2(n977), 
            .I3(n23241), .O(n7592[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_14 (.CI(n23241), .I0(n7608[11]), .I1(n977), .CO(n23242));
    SB_LUT4 add_3496_13_lut (.I0(GND_net), .I1(n7608[10]), .I2(n904), 
            .I3(n23240), .O(n7592[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_13 (.CI(n23240), .I0(n7608[10]), .I1(n904), .CO(n23241));
    SB_LUT4 add_3496_12_lut (.I0(GND_net), .I1(n7608[9]), .I2(n831), .I3(n23239), 
            .O(n7592[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_12 (.CI(n23239), .I0(n7608[9]), .I1(n831), .CO(n23240));
    SB_LUT4 add_3496_11_lut (.I0(GND_net), .I1(n7608[8]), .I2(n758), .I3(n23238), 
            .O(n7592[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_11 (.CI(n23238), .I0(n7608[8]), .I1(n758), .CO(n23239));
    SB_LUT4 add_3496_10_lut (.I0(GND_net), .I1(n7608[7]), .I2(n685), .I3(n23237), 
            .O(n7592[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_10 (.CI(n23237), .I0(n7608[7]), .I1(n685), .CO(n23238));
    SB_LUT4 add_3496_9_lut (.I0(GND_net), .I1(n7608[6]), .I2(n612), .I3(n23236), 
            .O(n7592[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_9 (.CI(n23236), .I0(n7608[6]), .I1(n612), .CO(n23237));
    SB_LUT4 add_3496_8_lut (.I0(GND_net), .I1(n7608[5]), .I2(n539), .I3(n23235), 
            .O(n7592[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_8 (.CI(n23235), .I0(n7608[5]), .I1(n539), .CO(n23236));
    SB_LUT4 add_3496_7_lut (.I0(GND_net), .I1(n7608[4]), .I2(n466), .I3(n23234), 
            .O(n7592[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n22482), .I0(motor_state[17]), 
            .I1(n1[17]), .CO(n22483));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1[16]), .I3(n22481), .O(\PID_CONTROLLER.err_23__N_3556 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_25_lut (.I0(GND_net), .I1(n2908[23]), .I2(n2933[23]), 
            .I3(n22535), .O(duty_23__N_3655[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_24_lut (.I0(GND_net), .I1(n2908[22]), .I2(n2933[22]), 
            .I3(n22534), .O(duty_23__N_3655[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_24 (.CI(n22534), .I0(n2908[22]), .I1(n2933[22]), 
            .CO(n22535));
    SB_CARRY add_3496_7 (.CI(n23234), .I0(n7608[4]), .I1(n466), .CO(n23235));
    SB_LUT4 add_3496_6_lut (.I0(GND_net), .I1(n7608[3]), .I2(n393), .I3(n23233), 
            .O(n7592[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_6 (.CI(n23233), .I0(n7608[3]), .I1(n393), .CO(n23234));
    SB_LUT4 add_3496_5_lut (.I0(GND_net), .I1(n7608[2]), .I2(n320), .I3(n23232), 
            .O(n7592[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_5 (.CI(n23232), .I0(n7608[2]), .I1(n320), .CO(n23233));
    SB_LUT4 add_3496_4_lut (.I0(GND_net), .I1(n7608[1]), .I2(n247), .I3(n23231), 
            .O(n7592[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_4 (.CI(n23231), .I0(n7608[1]), .I1(n247), .CO(n23232));
    SB_LUT4 add_3496_3_lut (.I0(GND_net), .I1(n7608[0]), .I2(n174), .I3(n23230), 
            .O(n7592[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_3 (.CI(n23230), .I0(n7608[0]), .I1(n174), .CO(n23231));
    SB_LUT4 add_3496_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n7592[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3496_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3496_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n23230));
    SB_LUT4 add_3495_16_lut (.I0(GND_net), .I1(n7592[13]), .I2(n1120), 
            .I3(n23229), .O(n7575[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3495_15_lut (.I0(GND_net), .I1(n7592[12]), .I2(n1047), 
            .I3(n23228), .O(n7575[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_15 (.CI(n23228), .I0(n7592[12]), .I1(n1047), .CO(n23229));
    SB_LUT4 add_3495_14_lut (.I0(GND_net), .I1(n7592[11]), .I2(n974), 
            .I3(n23227), .O(n7575[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_14 (.CI(n23227), .I0(n7592[11]), .I1(n974), .CO(n23228));
    SB_LUT4 add_3495_13_lut (.I0(GND_net), .I1(n7592[10]), .I2(n901), 
            .I3(n23226), .O(n7575[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_13 (.CI(n23226), .I0(n7592[10]), .I1(n901), .CO(n23227));
    SB_LUT4 add_3495_12_lut (.I0(GND_net), .I1(n7592[9]), .I2(n828), .I3(n23225), 
            .O(n7575[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_12 (.CI(n23225), .I0(n7592[9]), .I1(n828), .CO(n23226));
    SB_LUT4 add_3495_11_lut (.I0(GND_net), .I1(n7592[8]), .I2(n755), .I3(n23224), 
            .O(n7575[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_11 (.CI(n23224), .I0(n7592[8]), .I1(n755), .CO(n23225));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n22481), .I0(motor_state[16]), 
            .I1(n1[16]), .CO(n22482));
    SB_LUT4 add_616_23_lut (.I0(GND_net), .I1(n2908[21]), .I2(n2933[21]), 
            .I3(n22533), .O(duty_23__N_3655[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1[15]), .I3(n22480), .O(\PID_CONTROLLER.err_23__N_3556 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n22480), .I0(motor_state[15]), 
            .I1(n1[15]), .CO(n22481));
    SB_CARRY add_616_23 (.CI(n22533), .I0(n2908[21]), .I1(n2933[21]), 
            .CO(n22534));
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1[14]), .I3(n22479), .O(\PID_CONTROLLER.err_23__N_3556 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_22_lut (.I0(GND_net), .I1(n2908[20]), .I2(n2933[20]), 
            .I3(n22532), .O(duty_23__N_3655[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_22 (.CI(n22532), .I0(n2908[20]), .I1(n2933[20]), 
            .CO(n22533));
    SB_LUT4 add_616_21_lut (.I0(GND_net), .I1(n2908[19]), .I2(n2933[19]), 
            .I3(n22531), .O(duty_23__N_3655[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n22479), .I0(motor_state[14]), 
            .I1(n1[14]), .CO(n22480));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1[13]), .I3(n22478), .O(\PID_CONTROLLER.err_23__N_3556 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_21 (.CI(n22531), .I0(n2908[19]), .I1(n2933[19]), 
            .CO(n22532));
    SB_LUT4 add_616_20_lut (.I0(GND_net), .I1(n2908[18]), .I2(n2933[18]), 
            .I3(n22530), .O(duty_23__N_3655[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_20 (.CI(n22530), .I0(n2908[18]), .I1(n2933[18]), 
            .CO(n22531));
    SB_CARRY state_23__I_0_add_2_15 (.CI(n22478), .I0(motor_state[13]), 
            .I1(n1[13]), .CO(n22479));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1[12]), .I3(n22477), .O(\PID_CONTROLLER.err_23__N_3556 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_19_lut (.I0(GND_net), .I1(n2908[17]), .I2(n2933[17]), 
            .I3(n22529), .O(duty_23__N_3655[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n22477), .I0(motor_state[12]), 
            .I1(n1[12]), .CO(n22478));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1[11]), .I3(n22476), .O(\PID_CONTROLLER.err_23__N_3556 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n22476), .I0(motor_state[11]), 
            .I1(n1[11]), .CO(n22477));
    SB_CARRY add_616_19 (.CI(n22529), .I0(n2908[17]), .I1(n2933[17]), 
            .CO(n22530));
    SB_LUT4 add_616_18_lut (.I0(GND_net), .I1(n2908[16]), .I2(n2933[16]), 
            .I3(n22528), .O(duty_23__N_3655[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1[10]), .I3(n22475), .O(\PID_CONTROLLER.err_23__N_3556 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1_adj_4607[23]), 
            .I3(n22604), .O(n47_adj_4180)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3495_10_lut (.I0(GND_net), .I1(n7592[7]), .I2(n682), .I3(n23223), 
            .O(n7575[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_10 (.CI(n23223), .I0(n7592[7]), .I1(n682), .CO(n23224));
    SB_LUT4 add_3495_9_lut (.I0(GND_net), .I1(n7592[6]), .I2(n609), .I3(n23222), 
            .O(n7575[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_9 (.CI(n23222), .I0(n7592[6]), .I1(n609), .CO(n23223));
    SB_LUT4 add_3495_8_lut (.I0(GND_net), .I1(n7592[5]), .I2(n536), .I3(n23221), 
            .O(n7575[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_8 (.CI(n23221), .I0(n7592[5]), .I1(n536), .CO(n23222));
    SB_LUT4 add_3495_7_lut (.I0(GND_net), .I1(n7592[4]), .I2(n463), .I3(n23220), 
            .O(n7575[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_7 (.CI(n23220), .I0(n7592[4]), .I1(n463), .CO(n23221));
    SB_LUT4 add_3495_6_lut (.I0(GND_net), .I1(n7592[3]), .I2(n390), .I3(n23219), 
            .O(n7575[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_6 (.CI(n23219), .I0(n7592[3]), .I1(n390), .CO(n23220));
    SB_LUT4 add_3495_5_lut (.I0(GND_net), .I1(n7592[2]), .I2(n317), .I3(n23218), 
            .O(n7575[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_5 (.CI(n23218), .I0(n7592[2]), .I1(n317), .CO(n23219));
    SB_LUT4 add_3495_4_lut (.I0(GND_net), .I1(n7592[1]), .I2(n244), .I3(n23217), 
            .O(n7575[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_4 (.CI(n23217), .I0(n7592[1]), .I1(n244), .CO(n23218));
    SB_LUT4 add_3495_3_lut (.I0(GND_net), .I1(n7592[0]), .I2(n171), .I3(n23216), 
            .O(n7575[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_3 (.CI(n23216), .I0(n7592[0]), .I1(n171), .CO(n23217));
    SB_LUT4 add_3495_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n7575[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3495_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3495_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n23216));
    SB_LUT4 add_3494_17_lut (.I0(GND_net), .I1(n7575[14]), .I2(GND_net), 
            .I3(n23215), .O(n7557[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3494_16_lut (.I0(GND_net), .I1(n7575[13]), .I2(n1117), 
            .I3(n23214), .O(n7557[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_16 (.CI(n23214), .I0(n7575[13]), .I1(n1117), .CO(n23215));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[22]), 
            .I3(n22603), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_18 (.CI(n22528), .I0(n2908[16]), .I1(n2933[16]), 
            .CO(n22529));
    SB_LUT4 add_3494_15_lut (.I0(GND_net), .I1(n7575[12]), .I2(n1044), 
            .I3(n23213), .O(n7557[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n22603), .I0(GND_net), .I1(n1_adj_4607[22]), 
            .CO(n22604));
    SB_CARRY add_3494_15 (.CI(n23213), .I0(n7575[12]), .I1(n1044), .CO(n23214));
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[21]), 
            .I3(n22602), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4182));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n22602), .I0(GND_net), .I1(n1_adj_4607[21]), 
            .CO(n22603));
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[20]), 
            .I3(n22601), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4184));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_616_17_lut (.I0(GND_net), .I1(n2908[15]), .I2(n2933[15]), 
            .I3(n22527), .O(duty_23__N_3655[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3494_14_lut (.I0(GND_net), .I1(n7575[11]), .I2(n971), 
            .I3(n23212), .O(n7557[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24196_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n30048));
    defparam i24196_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_3494_14 (.CI(n23212), .I0(n7575[11]), .I1(n971), .CO(n23213));
    SB_LUT4 i24193_3_lut (.I0(n11_adj_4184), .I1(n9_adj_4182), .I2(n30048), 
            .I3(GND_net), .O(n30045));
    defparam i24193_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 add_3494_13_lut (.I0(GND_net), .I1(n7575[10]), .I2(n898), 
            .I3(n23211), .O(n7557[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_162_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n31459));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_162_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24534_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n31459), 
            .I2(IntegralLimit[7]), .I3(n30045), .O(n30387));
    defparam i24534_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i24438_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n30387), .O(n30291));
    defparam i24438_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_144_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n31441));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_144_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24436_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n9_adj_4182), .O(n30289));
    defparam i24436_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_3494_13 (.CI(n23211), .I0(n7575[10]), .I1(n898), .CO(n23212));
    SB_LUT4 add_3494_12_lut (.I0(GND_net), .I1(n7575[9]), .I2(n825), .I3(n23210), 
            .O(n7557[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24434_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n31441), 
            .I2(IntegralLimit[11]), .I3(n30289), .O(n30287));
    defparam i24434_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_138_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n31435));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_138_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24144_4_lut (.I0(n27), .I1(n15_adj_4185), .I2(n13_adj_4186), 
            .I3(n11_adj_4187), .O(n29996));
    defparam i24144_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24150_4_lut (.I0(n21_adj_4188), .I1(n19), .I2(n17_adj_4189), 
            .I3(n9_adj_4190), .O(n30002));
    defparam i24150_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24125_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n29977));
    defparam i24125_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4189), .I3(GND_net), 
            .O(n8_adj_4191));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_4192));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24160_2_lut (.I0(n7_adj_4193), .I1(n5_adj_4194), .I2(GND_net), 
            .I3(GND_net), .O(n30012));
    defparam i24160_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_3494_12 (.CI(n23210), .I0(n7575[9]), .I1(n825), .CO(n23211));
    SB_LUT4 i24410_4_lut (.I0(n13_adj_4186), .I1(n11_adj_4187), .I2(n9_adj_4190), 
            .I3(n30012), .O(n30263));
    defparam i24410_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_3494_11_lut (.I0(GND_net), .I1(n7575[8]), .I2(n752), .I3(n23209), 
            .O(n7557[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_11 (.CI(n23209), .I0(n7575[8]), .I1(n752), .CO(n23210));
    SB_LUT4 add_3494_10_lut (.I0(GND_net), .I1(n7575[7]), .I2(n679), .I3(n23208), 
            .O(n7557[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24406_4_lut (.I0(n19), .I1(n17_adj_4189), .I2(n15_adj_4185), 
            .I3(n30263), .O(n30259));
    defparam i24406_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24637_4_lut (.I0(n25_c), .I1(n23_adj_4195), .I2(n21_adj_4188), 
            .I3(n30259), .O(n30490));
    defparam i24637_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24512_4_lut (.I0(n31), .I1(n29_adj_4196), .I2(n27), .I3(n30490), 
            .O(n30365));
    defparam i24512_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24661_4_lut (.I0(n37), .I1(n35_adj_4197), .I2(n33), .I3(n30365), 
            .O(n30514));
    defparam i24661_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24440_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n31459), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4184), .O(n30293));
    defparam i24440_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_131_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n31428));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_131_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24428_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n31428), 
            .I2(IntegralLimit[14]), .I3(n30293), .O(n30281));
    defparam i24428_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_126_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n31423));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_126_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4198));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24173_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n30025));
    defparam i24173_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_149_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n31446));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_149_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4199));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4198), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24584_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n31441), 
            .I2(IntegralLimit[11]), .I3(n30291), .O(n30437));
    defparam i24584_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i24181_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n31435), 
            .I2(IntegralLimit[13]), .I3(n30437), .O(n30033));
    defparam i24181_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_129_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n31426));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_129_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24528_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n31426), 
            .I2(IntegralLimit[15]), .I3(n30033), .O(n30381));
    defparam i24528_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_155_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n31452));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_155_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24641_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n31452), 
            .I2(IntegralLimit[17]), .I3(n30381), .O(n30494));
    defparam i24641_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mux_614_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_120_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n31417));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_120_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24683_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n31417), 
            .I2(IntegralLimit[19]), .I3(n30494), .O(n30536));
    defparam i24683_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_117_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n31414));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_117_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4201));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24162_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n30014));
    defparam i24162_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4201), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4202));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4203));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24554_3_lut (.I0(n6_adj_4203), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n30407));   // verilog/motorControl.v(31[10:34])
    defparam i24554_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24555_3_lut (.I0(n30407), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n30408));   // verilog/motorControl.v(31[10:34])
    defparam i24555_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24164_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n31435), 
            .I2(IntegralLimit[21]), .I3(n30287), .O(n30016));
    defparam i24164_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i24490_4_lut (.I0(n24_adj_4202), .I1(n8_adj_4204), .I2(n31412), 
            .I3(n30014), .O(n30343));   // verilog/motorControl.v(31[10:34])
    defparam i24490_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24347_3_lut (.I0(n30408), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n30200));   // verilog/motorControl.v(31[10:34])
    defparam i24347_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3521_6_lut (.I0(GND_net), .I1(n7947[3]), .I2(n402_adj_4205), 
            .I3(n23512), .O(n7934[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3631 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4206), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4207));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i24544_3_lut (.I0(n4_adj_4207), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n30397));   // verilog/motorControl.v(31[38:63])
    defparam i24544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24545_3_lut (.I0(n30397), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4196), .I3(GND_net), .O(n30398));   // verilog/motorControl.v(31[38:63])
    defparam i24545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4208));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24138_2_lut (.I0(n33), .I1(n15_adj_4185), .I2(GND_net), .I3(GND_net), 
            .O(n29990));
    defparam i24138_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4186), .I3(GND_net), 
            .O(n10_adj_4209));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4208), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4197), .I3(GND_net), 
            .O(n30_adj_4210));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_3494_10 (.CI(n23208), .I0(n7575[7]), .I1(n679), .CO(n23209));
    SB_LUT4 add_3494_9_lut (.I0(GND_net), .I1(n7575[6]), .I2(n606), .I3(n23207), 
            .O(n7557[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24140_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4196), .I3(n29996), 
            .O(n29992));
    defparam i24140_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24651_4_lut (.I0(n30_adj_4210), .I1(n10_adj_4209), .I2(n35_adj_4197), 
            .I3(n29990), .O(n30504));   // verilog/motorControl.v(31[38:63])
    defparam i24651_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24359_3_lut (.I0(n30398), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n30212));   // verilog/motorControl.v(31[38:63])
    defparam i24359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24691_4_lut (.I0(n30212), .I1(n30504), .I2(n35_adj_4197), 
            .I3(n29992), .O(n30544));   // verilog/motorControl.v(31[38:63])
    defparam i24691_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24692_3_lut (.I0(n30544), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n30545));   // verilog/motorControl.v(31[38:63])
    defparam i24692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24672_3_lut (.I0(n30545), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n30525));   // verilog/motorControl.v(31[38:63])
    defparam i24672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4193), .I3(GND_net), 
            .O(n6_adj_4211));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24546_3_lut (.I0(n6_adj_4211), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4188), .I3(GND_net), .O(n30399));   // verilog/motorControl.v(31[38:63])
    defparam i24546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24547_3_lut (.I0(n30399), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4195), .I3(GND_net), .O(n30400));   // verilog/motorControl.v(31[38:63])
    defparam i24547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24127_4_lut (.I0(n43), .I1(n25_c), .I2(n23_adj_4195), .I3(n30002), 
            .O(n29979));
    defparam i24127_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24492_4_lut (.I0(n24_adj_4192), .I1(n8_adj_4191), .I2(n45), 
            .I3(n29977), .O(n30345));   // verilog/motorControl.v(31[38:63])
    defparam i24492_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24357_3_lut (.I0(n30400), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_c), .I3(GND_net), .O(n30210));   // verilog/motorControl.v(31[38:63])
    defparam i24357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24130_4_lut (.I0(n43), .I1(n41_adj_4212), .I2(n39), .I3(n30514), 
            .O(n29982));
    defparam i24130_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24617_4_lut (.I0(n30210), .I1(n30345), .I2(n45), .I3(n29979), 
            .O(n30470));   // verilog/motorControl.v(31[38:63])
    defparam i24617_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24365_3_lut (.I0(n30525), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4212), .I3(GND_net), .O(n30218));   // verilog/motorControl.v(31[38:63])
    defparam i24365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24659_4_lut (.I0(n30218), .I1(n30470), .I2(n45), .I3(n29982), 
            .O(n30512));   // verilog/motorControl.v(31[38:63])
    defparam i24659_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4213));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i24552_3_lut (.I0(n4_adj_4213), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n30405));   // verilog/motorControl.v(31[10:34])
    defparam i24552_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24553_3_lut (.I0(n30405), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n30406));   // verilog/motorControl.v(31[10:34])
    defparam i24553_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24175_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n31423), 
            .I2(IntegralLimit[16]), .I3(n30281), .O(n30027));
    defparam i24175_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i24649_4_lut (.I0(n30), .I1(n10_adj_4199), .I2(n31446), .I3(n30025), 
            .O(n30502));   // verilog/motorControl.v(31[10:34])
    defparam i24649_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24349_3_lut (.I0(n30406), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n30202));   // verilog/motorControl.v(31[10:34])
    defparam i24349_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24689_4_lut (.I0(n30202), .I1(n30502), .I2(n31446), .I3(n30027), 
            .O(n30542));   // verilog/motorControl.v(31[10:34])
    defparam i24689_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24690_3_lut (.I0(n30542), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n30543));   // verilog/motorControl.v(31[10:34])
    defparam i24690_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24674_3_lut (.I0(n30543), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n30527));   // verilog/motorControl.v(31[10:34])
    defparam i24674_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24166_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n31414), 
            .I2(IntegralLimit[21]), .I3(n30536), .O(n30018));
    defparam i24166_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_115_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n31412));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_115_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24615_4_lut (.I0(n30200), .I1(n30343), .I2(n31412), .I3(n30016), 
            .O(n30468));   // verilog/motorControl.v(31[10:34])
    defparam i24615_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24355_3_lut (.I0(n30527), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n30208));   // verilog/motorControl.v(31[10:34])
    defparam i24355_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24660_3_lut (.I0(n30512), .I1(\PID_CONTROLLER.integral_23__N_3631 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3630 ));   // verilog/motorControl.v(31[38:63])
    defparam i24660_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24657_4_lut (.I0(n30208), .I1(n30468), .I2(n31412), .I3(n30018), 
            .O(n30510));   // verilog/motorControl.v(31[10:34])
    defparam i24657_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_838_4_lut  (.I0(n30510), .I1(\PID_CONTROLLER.integral_23__N_3630 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3628 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_838_4_lut .LUT_INIT = 16'h80c8;
    SB_CARRY add_616_17 (.CI(n22527), .I0(n2908[15]), .I1(n2933[15]), 
            .CO(n22528));
    SB_CARRY add_3494_9 (.CI(n23207), .I0(n7575[6]), .I1(n606), .CO(n23208));
    SB_LUT4 add_3494_8_lut (.I0(GND_net), .I1(n7575[5]), .I2(n533), .I3(n23206), 
            .O(n7557[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_8 (.CI(n23206), .I0(n7575[5]), .I1(n533), .CO(n23207));
    SB_LUT4 add_3494_7_lut (.I0(GND_net), .I1(n7575[4]), .I2(n460), .I3(n23205), 
            .O(n7557[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_7 (.CI(n23205), .I0(n7575[4]), .I1(n460), .CO(n23206));
    SB_LUT4 add_3494_6_lut (.I0(GND_net), .I1(n7575[3]), .I2(n387), .I3(n23204), 
            .O(n7557[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_16_lut (.I0(GND_net), .I1(n2908[14]), .I2(n2933[14]), 
            .I3(n22526), .O(duty_23__N_3655[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_6 (.CI(n23204), .I0(n7575[3]), .I1(n387), .CO(n23205));
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4214));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3494_5_lut (.I0(GND_net), .I1(n7575[2]), .I2(n314), .I3(n23203), 
            .O(n7557[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4216));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4217));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3494_5 (.CI(n23203), .I0(n7575[2]), .I1(n314), .CO(n23204));
    SB_LUT4 add_3494_4_lut (.I0(GND_net), .I1(n7575[1]), .I2(n241), .I3(n23202), 
            .O(n7557[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_4 (.CI(n23202), .I0(n7575[1]), .I1(n241), .CO(n23203));
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4218));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3494_3_lut (.I0(GND_net), .I1(n7575[0]), .I2(n168), .I3(n23201), 
            .O(n7557[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3494_3 (.CI(n23201), .I0(n7575[0]), .I1(n168), .CO(n23202));
    SB_LUT4 add_3494_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n7557[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3494_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3494_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n23201));
    SB_LUT4 add_3493_18_lut (.I0(GND_net), .I1(n7557[15]), .I2(GND_net), 
            .I3(n23200), .O(n7538[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3493_17_lut (.I0(GND_net), .I1(n7557[14]), .I2(GND_net), 
            .I3(n23199), .O(n7538[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_17 (.CI(n23199), .I0(n7557[14]), .I1(GND_net), .CO(n23200));
    SB_LUT4 add_3493_16_lut (.I0(GND_net), .I1(n7557[13]), .I2(n1114), 
            .I3(n23198), .O(n7538[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_16 (.CI(n23198), .I0(n7557[13]), .I1(n1114), .CO(n23199));
    SB_LUT4 add_3493_15_lut (.I0(GND_net), .I1(n7557[12]), .I2(n1041), 
            .I3(n23197), .O(n7538[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_15 (.CI(n23197), .I0(n7557[12]), .I1(n1041), .CO(n23198));
    SB_LUT4 add_3493_14_lut (.I0(GND_net), .I1(n7557[11]), .I2(n968), 
            .I3(n23196), .O(n7538[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_14 (.CI(n23196), .I0(n7557[11]), .I1(n968), .CO(n23197));
    SB_LUT4 add_3493_13_lut (.I0(GND_net), .I1(n7557[10]), .I2(n895), 
            .I3(n23195), .O(n7538[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_13 (.CI(n23195), .I0(n7557[10]), .I1(n895), .CO(n23196));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n22601), .I0(GND_net), .I1(n1_adj_4607[20]), 
            .CO(n22602));
    SB_LUT4 add_3493_12_lut (.I0(GND_net), .I1(n7557[9]), .I2(n822), .I3(n23194), 
            .O(n7538[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_12 (.CI(n23194), .I0(n7557[9]), .I1(n822), .CO(n23195));
    SB_LUT4 add_3493_11_lut (.I0(GND_net), .I1(n7557[8]), .I2(n749), .I3(n23193), 
            .O(n7538[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n22475), .I0(motor_state[10]), 
            .I1(n1[10]), .CO(n22476));
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4219));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1[9]), .I3(n22474), .O(\PID_CONTROLLER.err_23__N_3556 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n22474), .I0(motor_state[9]), .I1(n1[9]), 
            .CO(n22475));
    SB_CARRY add_616_16 (.CI(n22526), .I0(n2908[14]), .I1(n2933[14]), 
            .CO(n22527));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1[8]), .I3(n22473), .O(\PID_CONTROLLER.err_23__N_3556 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_11 (.CI(n23193), .I0(n7557[8]), .I1(n749), .CO(n23194));
    SB_LUT4 add_3493_10_lut (.I0(GND_net), .I1(n7557[7]), .I2(n676), .I3(n23192), 
            .O(n7538[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_10 (.CI(n23192), .I0(n7557[7]), .I1(n676), .CO(n23193));
    SB_LUT4 add_3493_9_lut (.I0(GND_net), .I1(n7557[6]), .I2(n603), .I3(n23191), 
            .O(n7538[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_9 (.CI(n23191), .I0(n7557[6]), .I1(n603), .CO(n23192));
    SB_LUT4 add_3493_8_lut (.I0(GND_net), .I1(n7557[5]), .I2(n530), .I3(n23190), 
            .O(n7538[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_8 (.CI(n23190), .I0(n7557[5]), .I1(n530), .CO(n23191));
    SB_LUT4 add_3493_7_lut (.I0(GND_net), .I1(n7557[4]), .I2(n457), .I3(n23189), 
            .O(n7538[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_7 (.CI(n23189), .I0(n7557[4]), .I1(n457), .CO(n23190));
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3493_6_lut (.I0(GND_net), .I1(n7557[3]), .I2(n384), .I3(n23188), 
            .O(n7538[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_6 (.CI(n23188), .I0(n7557[3]), .I1(n384), .CO(n23189));
    SB_LUT4 add_3493_5_lut (.I0(GND_net), .I1(n7557[2]), .I2(n311), .I3(n23187), 
            .O(n7538[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_15_lut (.I0(GND_net), .I1(n2908[13]), .I2(n2933[13]), 
            .I3(n22525), .O(duty_23__N_3655[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3493_5 (.CI(n23187), .I0(n7557[2]), .I1(n311), .CO(n23188));
    SB_LUT4 add_3493_4_lut (.I0(GND_net), .I1(n7557[1]), .I2(n238), .I3(n23186), 
            .O(n7538[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3493_4 (.CI(n23186), .I0(n7557[1]), .I1(n238), .CO(n23187));
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3493_3_lut (.I0(GND_net), .I1(n7557[0]), .I2(n165), .I3(n23185), 
            .O(n7538[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4226));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4227));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4228));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4229));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4231));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4233));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4234));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4235));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4237));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4238));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4239));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4240));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3493_3 (.CI(n23185), .I0(n7557[0]), .I1(n165), .CO(n23186));
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4241));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4242));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4243));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4244));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3493_2_lut (.I0(GND_net), .I1(n23_adj_4245), .I2(n92), 
            .I3(GND_net), .O(n7538[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3493_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4246));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3493_2 (.CI(GND_net), .I0(n23_adj_4245), .I1(n92), .CO(n23185));
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4247));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3492_19_lut (.I0(GND_net), .I1(n7538[16]), .I2(GND_net), 
            .I3(n23184), .O(n7518[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4252));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4253));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4254));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4255));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[0]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[1]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_614_i1_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256_adj_4200), .I3(\Ki[0] ), .O(n2933[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i14152_3_lut (.I0(\Kp[0] ), .I1(n256_adj_4200), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n2908[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam i14152_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4263));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4264));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4265));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4266));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4267));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4268));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4269));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4270));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4271));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n22473), .I0(motor_state[8]), .I1(n1[8]), 
            .CO(n22474));
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4272));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4273));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_616_15 (.CI(n22525), .I0(n2908[13]), .I1(n2933[13]), 
            .CO(n22526));
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4274));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4275));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4276));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4277));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4278));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[2]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[3]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_614_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3492_18_lut (.I0(GND_net), .I1(n7538[15]), .I2(GND_net), 
            .I3(n23183), .O(n7518[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4281));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3492_18 (.CI(n23183), .I0(n7538[15]), .I1(GND_net), .CO(n23184));
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4282));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4283));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4284));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4285));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4286));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4287));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4288));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4289));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3492_17_lut (.I0(GND_net), .I1(n7538[14]), .I2(GND_net), 
            .I3(n23182), .O(n7518[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3492_17 (.CI(n23182), .I0(n7538[14]), .I1(GND_net), .CO(n23183));
    SB_LUT4 add_3492_16_lut (.I0(GND_net), .I1(n7538[13]), .I2(n1111), 
            .I3(n23181), .O(n7518[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[4]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[5]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[6]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[7]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[8]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[9]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_614_i5_3_lut (.I0(n155[4]), .I1(PWMLimit[4]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i5_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[10]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14374_1_lut (.I0(n256_adj_4200), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18939));   // verilog/motorControl.v(38[19:35])
    defparam i14374_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4297));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4298));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4299));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4300));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4301));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[11]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4303));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4304));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4305));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4306));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4307));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4308));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4309));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i6_3_lut (.I0(n155[5]), .I1(PWMLimit[5]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4310));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4311));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4312));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4313));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[12]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4315));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4316));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4317));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4318));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4319));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4320));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4321));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4323));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[13]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4325));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4326));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4327));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4328));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4329));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4330));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4331));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4332));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4333));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4334));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4335), .I1(\Ki[4] ), .I2(n8004[2]), .I3(\PID_CONTROLLER.integral [18]), 
            .O(n7997[3]));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4336));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4337));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4339));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4340));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4341));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4342));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4343));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4344));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4345));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4346));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4347));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4348));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4349));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4350));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4351));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4353));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4354));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4355));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4356));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[14]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4359));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17701_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n8015[0]));   // verilog/motorControl.v(34[26:37])
    defparam i17701_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4360));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3492_16 (.CI(n23181), .I0(n7538[13]), .I1(n1111), .CO(n23182));
    SB_LUT4 add_3492_15_lut (.I0(GND_net), .I1(n7538[12]), .I2(n1038), 
            .I3(n23180), .O(n7518[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_15 (.CI(n23180), .I0(n7538[12]), .I1(n1038), .CO(n23181));
    SB_LUT4 add_3492_14_lut (.I0(GND_net), .I1(n7538[11]), .I2(n965), 
            .I3(n23179), .O(n7518[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1483 (.I0(n4_adj_4361), .I1(\Ki[3] ), .I2(n8010[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n8004[2]));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1483.LUT_INIT = 16'h965a;
    SB_CARRY add_3492_14 (.CI(n23179), .I0(n7538[11]), .I1(n965), .CO(n23180));
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4362));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3492_13_lut (.I0(GND_net), .I1(n7538[10]), .I2(n892), 
            .I3(n23178), .O(n7518[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1484 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_4363));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1484.LUT_INIT = 16'h9c50;
    SB_LUT4 i17637_4_lut (.I0(n8004[2]), .I1(\Ki[4] ), .I2(n6_adj_4335), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_4364));   // verilog/motorControl.v(34[26:37])
    defparam i17637_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_4365));   // verilog/motorControl.v(34[26:37])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i17668_4_lut (.I0(n8010[1]), .I1(\Ki[3] ), .I2(n4_adj_4361), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_4366));   // verilog/motorControl.v(34[26:37])
    defparam i17668_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i17703_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n22260));   // verilog/motorControl.v(34[26:37])
    defparam i17703_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4366), .I1(n11_adj_4365), .I2(n8_adj_4364), 
            .I3(n12_adj_4363), .O(n18_adj_4367));   // verilog/motorControl.v(34[26:37])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_4368));   // verilog/motorControl.v(34[26:37])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4368), .I1(n18_adj_4367), .I2(n22260), 
            .I3(n4_adj_4369), .O(n28011));   // verilog/motorControl.v(34[26:37])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4370));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3512_17_lut (.I0(GND_net), .I1(n7794[14]), .I2(GND_net), 
            .I3(n23388), .O(n7772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_13 (.CI(n23178), .I0(n7538[10]), .I1(n892), .CO(n23179));
    SB_LUT4 add_3492_12_lut (.I0(GND_net), .I1(n7538[9]), .I2(n819), .I3(n23177), 
            .O(n7518[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4371));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4372));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3512_12 (.CI(n23383), .I0(n7794[9]), .I1(n813), .CO(n23384));
    SB_CARRY add_3512_11 (.CI(n23382), .I0(n7794[8]), .I1(n740_adj_4373), 
            .CO(n23383));
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4374));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3492_12 (.CI(n23177), .I0(n7538[9]), .I1(n819), .CO(n23178));
    SB_LUT4 add_3512_11_lut (.I0(GND_net), .I1(n7794[8]), .I2(n740_adj_4373), 
            .I3(n23382), .O(n7772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4375));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3492_11_lut (.I0(GND_net), .I1(n7538[8]), .I2(n746), .I3(n23176), 
            .O(n7518[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4376));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[19]), 
            .I3(n22600), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_11 (.CI(n23176), .I0(n7538[8]), .I1(n746), .CO(n23177));
    SB_LUT4 add_616_14_lut (.I0(GND_net), .I1(n2908[12]), .I2(n2933[12]), 
            .I3(n22524), .O(duty_23__N_3655[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_10_lut (.I0(GND_net), .I1(n7538[7]), .I2(n673), .I3(n23175), 
            .O(n7518[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4379));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3492_10 (.CI(n23175), .I0(n7538[7]), .I1(n673), .CO(n23176));
    SB_LUT4 add_3492_9_lut (.I0(GND_net), .I1(n7538[6]), .I2(n600), .I3(n23174), 
            .O(n7518[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_9 (.CI(n23174), .I0(n7538[6]), .I1(n600), .CO(n23175));
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4381));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[15]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_614_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3512_10_lut (.I0(GND_net), .I1(n7794[7]), .I2(n667_adj_4385), 
            .I3(n23381), .O(n7772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3492_8_lut (.I0(GND_net), .I1(n7538[5]), .I2(n527), .I3(n23173), 
            .O(n7518[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3492_8 (.CI(n23173), .I0(n7538[5]), .I1(n527), .CO(n23174));
    SB_LUT4 add_3492_7_lut (.I0(GND_net), .I1(n7538[4]), .I2(n454), .I3(n23172), 
            .O(n7518[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1[7]), .I3(n22472), .O(\PID_CONTROLLER.err_23__N_3556 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_7 (.CI(n23172), .I0(n7538[4]), .I1(n454), .CO(n23173));
    SB_LUT4 add_3492_6_lut (.I0(GND_net), .I1(n7538[3]), .I2(n381), .I3(n23171), 
            .O(n7518[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_6 (.CI(n23171), .I0(n7538[3]), .I1(n381), .CO(n23172));
    SB_CARRY add_3512_10 (.CI(n23381), .I0(n7794[7]), .I1(n667_adj_4385), 
            .CO(n23382));
    SB_CARRY add_3512_19 (.CI(n23390), .I0(n7794[16]), .I1(GND_net), .CO(n23391));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n22600), .I0(GND_net), .I1(n1_adj_4607[19]), 
            .CO(n22601));
    SB_LUT4 add_3512_7_lut (.I0(GND_net), .I1(n7794[4]), .I2(n448_adj_4387), 
            .I3(n23378), .O(n7772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_5_lut (.I0(GND_net), .I1(n7538[2]), .I2(n308), .I3(n23170), 
            .O(n7518[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3532[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_3492_5 (.CI(n23170), .I0(n7538[2]), .I1(n308), .CO(n23171));
    SB_LUT4 add_3492_4_lut (.I0(GND_net), .I1(n7538[1]), .I2(n235), .I3(n23169), 
            .O(n7518[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_4 (.CI(n23169), .I0(n7538[1]), .I1(n235), .CO(n23170));
    SB_LUT4 add_3492_3_lut (.I0(GND_net), .I1(n7538[0]), .I2(n162), .I3(n23168), 
            .O(n7518[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_14 (.CI(n22524), .I0(n2908[12]), .I1(n2933[12]), 
            .CO(n22525));
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3492_3 (.CI(n23168), .I0(n7538[0]), .I1(n162), .CO(n23169));
    SB_LUT4 add_3492_2_lut (.I0(GND_net), .I1(n20_adj_4389), .I2(n89), 
            .I3(GND_net), .O(n7518[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_614_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3492_2 (.CI(GND_net), .I0(n20_adj_4389), .I1(n89), .CO(n23168));
    SB_LUT4 add_3512_2_lut (.I0(GND_net), .I1(n14_adj_4390), .I2(n83_adj_4391), 
            .I3(GND_net), .O(n7772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_9 (.CI(n22472), .I0(motor_state[7]), .I1(n1[7]), 
            .CO(n22473));
    SB_CARRY add_3511_18 (.CI(n23369), .I0(n7772[15]), .I1(GND_net), .CO(n23370));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[18]), 
            .I3(n22599), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_17_lut (.I0(GND_net), .I1(n7772[14]), .I2(GND_net), 
            .I3(n23368), .O(n7749[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_2 (.CI(GND_net), .I0(n14_adj_4390), .I1(n83_adj_4391), 
            .CO(n23374));
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[16]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3491_20_lut (.I0(GND_net), .I1(n7518[17]), .I2(GND_net), 
            .I3(n23167), .O(n7497[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_19_lut (.I0(GND_net), .I1(n7518[16]), .I2(GND_net), 
            .I3(n23166), .O(n7497[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_19 (.CI(n23166), .I0(n7518[16]), .I1(GND_net), .CO(n23167));
    SB_CARRY add_3511_17 (.CI(n23368), .I0(n7772[14]), .I1(GND_net), .CO(n23369));
    SB_LUT4 add_3491_18_lut (.I0(GND_net), .I1(n7518[15]), .I2(GND_net), 
            .I3(n23165), .O(n7497[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_15_lut (.I0(GND_net), .I1(n7772[12]), .I2(n1029_adj_4395), 
            .I3(n23366), .O(n7749[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3491_18 (.CI(n23165), .I0(n7518[15]), .I1(GND_net), .CO(n23166));
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n22599), .I0(GND_net), .I1(n1_adj_4607[18]), 
            .CO(n22600));
    SB_CARRY add_3511_15 (.CI(n23366), .I0(n7772[12]), .I1(n1029_adj_4395), 
            .CO(n23367));
    SB_LUT4 add_616_13_lut (.I0(GND_net), .I1(n2908[11]), .I2(n2933[11]), 
            .I3(n22523), .O(duty_23__N_3655[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_22_lut (.I0(GND_net), .I1(n7772[19]), .I2(GND_net), 
            .I3(n23373), .O(n7749[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_17_lut (.I0(GND_net), .I1(n7518[14]), .I2(GND_net), 
            .I3(n23164), .O(n7497[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3491_17 (.CI(n23164), .I0(n7518[14]), .I1(GND_net), .CO(n23165));
    SB_LUT4 add_3491_16_lut (.I0(GND_net), .I1(n7518[13]), .I2(n1108), 
            .I3(n23163), .O(n7497[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_16 (.CI(n23163), .I0(n7518[13]), .I1(n1108), .CO(n23164));
    SB_CARRY add_616_13 (.CI(n22523), .I0(n2908[11]), .I1(n2933[11]), 
            .CO(n22524));
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[17]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4397));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3491_15_lut (.I0(GND_net), .I1(n7518[12]), .I2(n1035), 
            .I3(n23162), .O(n7497[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_7 (.CI(n23378), .I0(n7794[4]), .I1(n448_adj_4387), 
            .CO(n23379));
    SB_CARRY add_3491_15 (.CI(n23162), .I0(n7518[12]), .I1(n1035), .CO(n23163));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1[6]), .I3(n22471), .O(\PID_CONTROLLER.err_23__N_3556 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_14_lut (.I0(GND_net), .I1(n7518[11]), .I2(n962), 
            .I3(n23161), .O(n7497[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3491_14 (.CI(n23161), .I0(n7518[11]), .I1(n962), .CO(n23162));
    SB_LUT4 add_3491_13_lut (.I0(GND_net), .I1(n7518[10]), .I2(n889), 
            .I3(n23160), .O(n7497[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_13 (.CI(n23160), .I0(n7518[10]), .I1(n889), .CO(n23161));
    SB_LUT4 add_3491_12_lut (.I0(GND_net), .I1(n7518[9]), .I2(n816), .I3(n23159), 
            .O(n7497[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3511_21_lut (.I0(GND_net), .I1(n7772[18]), .I2(GND_net), 
            .I3(n23372), .O(n7749[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_16_lut (.I0(GND_net), .I1(n7772[13]), .I2(n1102_adj_4399), 
            .I3(n23367), .O(n7749[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3511_21 (.CI(n23372), .I0(n7772[18]), .I1(GND_net), .CO(n23373));
    SB_CARRY add_3491_12 (.CI(n23159), .I0(n7518[9]), .I1(n816), .CO(n23160));
    SB_LUT4 add_3512_6_lut (.I0(GND_net), .I1(n7794[3]), .I2(n375_adj_4397), 
            .I3(n23377), .O(n7772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4400));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4401));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n22471), .I0(motor_state[6]), .I1(n1[6]), 
            .CO(n22472));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[17]), 
            .I3(n22598), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_11_lut (.I0(GND_net), .I1(n7518[8]), .I2(n743), .I3(n23158), 
            .O(n7497[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4402));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_616_12_lut (.I0(GND_net), .I1(n2908[10]), .I2(n2933[10]), 
            .I3(n22522), .O(duty_23__N_3655[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1[5]), .I3(n22470), .O(\PID_CONTROLLER.err_23__N_3556 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n22598), .I0(GND_net), .I1(n1_adj_4607[17]), 
            .CO(n22599));
    SB_CARRY add_616_12 (.CI(n22522), .I0(n2908[10]), .I1(n2933[10]), 
            .CO(n22523));
    SB_CARRY add_3491_11 (.CI(n23158), .I0(n7518[8]), .I1(n743), .CO(n23159));
    SB_CARRY state_23__I_0_add_2_7 (.CI(n22470), .I0(motor_state[5]), .I1(n1[5]), 
            .CO(n22471));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[16]), 
            .I3(n22597), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_10_lut (.I0(GND_net), .I1(n7518[7]), .I2(n670), .I3(n23157), 
            .O(n7497[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4404));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_616_11_lut (.I0(GND_net), .I1(n2908[9]), .I2(n2933[9]), 
            .I3(n22521), .O(duty_23__N_3655[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1[4]), .I3(n22469), .O(\PID_CONTROLLER.err_23__N_3556 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_11 (.CI(n22521), .I0(n2908[9]), .I1(n2933[9]), .CO(n22522));
    SB_CARRY state_23__I_0_add_2_6 (.CI(n22469), .I0(motor_state[4]), .I1(n1[4]), 
            .CO(n22470));
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4399));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3491_10 (.CI(n23157), .I0(n7518[7]), .I1(n670), .CO(n23158));
    SB_LUT4 add_3491_9_lut (.I0(GND_net), .I1(n7518[6]), .I2(n597), .I3(n23156), 
            .O(n7497[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1[3]), .I3(n22468), .O(\PID_CONTROLLER.err_23__N_3556 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n22597), .I0(GND_net), .I1(n1_adj_4607[16]), 
            .CO(n22598));
    SB_LUT4 i24076_4_lut (.I0(n21_adj_4404), .I1(n19_adj_4402), .I2(n17_adj_4401), 
            .I3(n9_adj_4400), .O(n29928));
    defparam i24076_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_616_10_lut (.I0(GND_net), .I1(n2908[8]), .I2(n2933[8]), 
            .I3(n22520), .O(duty_23__N_3655[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_9 (.CI(n23156), .I0(n7518[6]), .I1(n597), .CO(n23157));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[15]), 
            .I3(n22596), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_8_lut (.I0(GND_net), .I1(n7518[5]), .I2(n524), .I3(n23155), 
            .O(n7497[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n23339), .I0(n7725[7]), .I1(n658_adj_4379), 
            .CO(n23340));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n7725[7]), .I2(n658_adj_4379), 
            .I3(n23339), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3521_7 (.CI(n23513), .I0(n7947[4]), .I1(n475_adj_4376), 
            .CO(n23514));
    SB_CARRY mult_11_add_1225_11 (.CI(n23340), .I0(n7725[8]), .I1(n731_adj_4375), 
            .CO(n23341));
    SB_LUT4 i24070_4_lut (.I0(n27_adj_4381), .I1(n15_adj_4370), .I2(n13_adj_4360), 
            .I3(n11_adj_4359), .O(n29922));
    defparam i24070_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4353), 
            .I3(GND_net), .O(n12_adj_4405));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3491_8 (.CI(n23155), .I0(n7518[5]), .I1(n524), .CO(n23156));
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4360), 
            .I3(GND_net), .O(n10_adj_4406));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4405), .I1(n257[17]), .I2(n35_adj_4344), 
            .I3(GND_net), .O(n30_adj_4407));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3491_7_lut (.I0(GND_net), .I1(n7518[4]), .I2(n451), .I3(n23154), 
            .O(n7497[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n22596), .I0(GND_net), .I1(n1_adj_4607[15]), 
            .CO(n22597));
    SB_CARRY state_23__I_0_add_2_5 (.CI(n22468), .I0(motor_state[3]), .I1(n1[3]), 
            .CO(n22469));
    SB_LUT4 add_3511_14_lut (.I0(GND_net), .I1(n7772[11]), .I2(n956_adj_4374), 
            .I3(n23365), .O(n7749[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_14 (.CI(n23365), .I0(n7772[11]), .I1(n956_adj_4374), 
            .CO(n23366));
    SB_CARRY add_3512_17 (.CI(n23388), .I0(n7794[14]), .I1(GND_net), .CO(n23389));
    SB_LUT4 add_3511_13_lut (.I0(GND_net), .I1(n7772[10]), .I2(n883_adj_4372), 
            .I3(n23364), .O(n7749[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_13 (.CI(n23364), .I0(n7772[10]), .I1(n883_adj_4372), 
            .CO(n23365));
    SB_LUT4 add_3511_12_lut (.I0(GND_net), .I1(n7772[9]), .I2(n810_adj_4371), 
            .I3(n23363), .O(n7749[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_12 (.CI(n23363), .I0(n7772[9]), .I1(n810_adj_4371), 
            .CO(n23364));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n7725[6]), .I2(n585), 
            .I3(n23338), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n7725[8]), .I2(n731_adj_4375), 
            .I3(n23340), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3526_7_lut (.I0(GND_net), .I1(n28011), .I2(n490_adj_4362), 
            .I3(n23553), .O(n7989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3526_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[14]), 
            .I3(n22595), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_10 (.CI(n22520), .I0(n2908[8]), .I1(n2933[8]), .CO(n22521));
    SB_CARRY add_3491_7 (.CI(n23154), .I0(n7518[4]), .I1(n451), .CO(n23155));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1[2]), .I3(n22467), .O(\PID_CONTROLLER.err_23__N_3556 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_6_lut (.I0(GND_net), .I1(n7518[3]), .I2(n378), .I3(n23153), 
            .O(n7497[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_20_lut (.I0(GND_net), .I1(n7772[17]), .I2(GND_net), 
            .I3(n23371), .O(n7749[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_6 (.CI(n23153), .I0(n7518[3]), .I1(n378), .CO(n23154));
    SB_LUT4 add_3491_5_lut (.I0(GND_net), .I1(n7518[2]), .I2(n305), .I3(n23152), 
            .O(n7497[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_5 (.CI(n23152), .I0(n7518[2]), .I1(n305), .CO(n23153));
    SB_LUT4 add_3525_2_lut (.I0(GND_net), .I1(n53_adj_4356), .I2(n122_adj_4355), 
            .I3(GND_net), .O(n7980[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3524_3_lut (.I0(GND_net), .I1(n7980[0]), .I2(n192_adj_4354), 
            .I3(n23536), .O(n7970[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_4_lut (.I0(GND_net), .I1(n7518[1]), .I2(n232), .I3(n23151), 
            .O(n7497[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_4 (.CI(n23151), .I0(n7518[1]), .I1(n232), .CO(n23152));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n22595), .I0(GND_net), .I1(n1_adj_4607[14]), 
            .CO(n22596));
    SB_CARRY add_3512_6 (.CI(n23377), .I0(n7794[3]), .I1(n375_adj_4397), 
            .CO(n23378));
    SB_LUT4 i24318_4_lut (.I0(n13_adj_4360), .I1(n11_adj_4359), .I2(n9_adj_4400), 
            .I3(n29938), .O(n30171));
    defparam i24318_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24314_4_lut (.I0(n19_adj_4402), .I1(n17_adj_4401), .I2(n15_adj_4370), 
            .I3(n30171), .O(n30167));
    defparam i24314_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24605_4_lut (.I0(n25_adj_4408), .I1(n23_adj_4409), .I2(n21_adj_4404), 
            .I3(n30167), .O(n30458));
    defparam i24605_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_616_9_lut (.I0(GND_net), .I1(n2908[7]), .I2(n2933[7]), 
            .I3(n22519), .O(duty_23__N_3655[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24472_4_lut (.I0(n31_adj_4331), .I1(n29_adj_4410), .I2(n27_adj_4381), 
            .I3(n30458), .O(n30325));
    defparam i24472_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY mult_11_add_1225_12 (.CI(n23341), .I0(n7725[9]), .I1(n804_adj_4351), 
            .CO(n23342));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n7725[11]), .I2(n950_adj_4350), 
            .I3(n23343), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_3_lut (.I0(GND_net), .I1(n7518[0]), .I2(n159), .I3(n23150), 
            .O(n7497[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3512_9_lut (.I0(GND_net), .I1(n7794[6]), .I2(n594_adj_4349), 
            .I3(n23380), .O(n7772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n7725[16]), .I2(GND_net), 
            .I3(n23348), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_4_lut (.I0(GND_net), .I1(n7772[1]), .I2(n226_adj_4348), 
            .I3(n23355), .O(n7749[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24653_4_lut (.I0(n37_adj_4411), .I1(n35_adj_4344), .I2(n33_adj_4353), 
            .I3(n30325), .O(n30506));
    defparam i24653_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3511_5 (.CI(n23356), .I0(n7772[2]), .I1(n299_adj_4347), 
            .CO(n23357));
    SB_CARRY add_3491_3 (.CI(n23150), .I0(n7518[0]), .I1(n159), .CO(n23151));
    SB_LUT4 add_3512_5_lut (.I0(GND_net), .I1(n7794[2]), .I2(n302_adj_4346), 
            .I3(n23376), .O(n7772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_2 (.CI(GND_net), .I0(n11_adj_4345), .I1(n80_adj_4343), 
            .CO(n23354));
    SB_LUT4 add_3511_5_lut (.I0(GND_net), .I1(n7772[2]), .I2(n299_adj_4347), 
            .I3(n23356), .O(n7749[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_20 (.CI(n23371), .I0(n7772[17]), .I1(GND_net), .CO(n23372));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n22467), .I0(motor_state[2]), .I1(n1[2]), 
            .CO(n22468));
    SB_LUT4 add_3511_2_lut (.I0(GND_net), .I1(n11_adj_4345), .I2(n80_adj_4343), 
            .I3(GND_net), .O(n7749[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n23349), .I0(n7725[17]), .I1(GND_net), 
            .CO(n23350));
    SB_CARRY add_3511_3 (.CI(n23354), .I0(n7772[0]), .I1(n153_adj_4342), 
            .CO(n23355));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n7725[17]), .I2(GND_net), 
            .I3(n23349), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n23344), .I0(n7725[12]), .I1(n1023_adj_4341), 
            .CO(n23345));
    SB_CARRY mult_11_add_1225_21 (.CI(n23350), .I0(n7725[18]), .I1(GND_net), 
            .CO(n23351));
    SB_LUT4 add_3511_3_lut (.I0(GND_net), .I1(n7772[0]), .I2(n153_adj_4342), 
            .I3(n23354), .O(n7749[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3491_2_lut (.I0(GND_net), .I1(n17_adj_4340), .I2(n86), 
            .I3(GND_net), .O(n7497[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3491_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4412), 
            .I3(GND_net), .O(n16_adj_4413));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3511_16 (.CI(n23367), .I0(n7772[13]), .I1(n1102_adj_4399), 
            .CO(n23368));
    SB_CARRY add_3511_6 (.CI(n23357), .I0(n7772[3]), .I1(n372_adj_4339), 
            .CO(n23358));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n7725[18]), .I2(GND_net), 
            .I3(n23350), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_19_lut (.I0(GND_net), .I1(n7772[16]), .I2(GND_net), 
            .I3(n23370), .O(n7749[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_5 (.CI(n23376), .I0(n7794[2]), .I1(n302_adj_4346), 
            .CO(n23377));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1[1]), .I3(n22466), .O(\PID_CONTROLLER.err_23__N_3556 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24593_3_lut (.I0(n6_adj_4415), .I1(n257[10]), .I2(n21_adj_4404), 
            .I3(GND_net), .O(n30446));   // verilog/motorControl.v(38[19:35])
    defparam i24593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3511_6_lut (.I0(GND_net), .I1(n7772[3]), .I2(n372_adj_4339), 
            .I3(n23357), .O(n7749[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_7 (.CI(n23358), .I0(n7772[4]), .I1(n445_adj_4337), 
            .CO(n23359));
    SB_LUT4 add_3511_7_lut (.I0(GND_net), .I1(n7772[4]), .I2(n445_adj_4337), 
            .I3(n23358), .O(n7749[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_8 (.CI(n23359), .I0(n7772[5]), .I1(n518_adj_4336), 
            .CO(n23360));
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n7725[12]), .I2(n1023_adj_4341), 
            .I3(n23344), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n23351), .I0(n7725[19]), .I1(GND_net), 
            .CO(n23352));
    SB_LUT4 i24594_3_lut (.I0(n30446), .I1(n257[11]), .I2(n23_adj_4409), 
            .I3(GND_net), .O(n30447));   // verilog/motorControl.v(38[19:35])
    defparam i24594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3526_6_lut (.I0(GND_net), .I1(n7997[3]), .I2(n417_adj_4334), 
            .I3(n23552), .O(n7989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3526_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3491_2 (.CI(GND_net), .I0(n17_adj_4340), .I1(n86), .CO(n23150));
    SB_LUT4 add_3490_21_lut (.I0(GND_net), .I1(n7497[18]), .I2(GND_net), 
            .I3(n23149), .O(n7475[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3511_8_lut (.I0(GND_net), .I1(n7772[5]), .I2(n518_adj_4336), 
            .I3(n23359), .O(n7749[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3490_20_lut (.I0(GND_net), .I1(n7497[17]), .I2(GND_net), 
            .I3(n23148), .O(n7475[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_20 (.CI(n23148), .I0(n7497[17]), .I1(GND_net), .CO(n23149));
    SB_LUT4 add_3490_19_lut (.I0(GND_net), .I1(n7497[16]), .I2(GND_net), 
            .I3(n23147), .O(n7475[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_19 (.CI(n23147), .I0(n7497[16]), .I1(GND_net), .CO(n23148));
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3490_18_lut (.I0(GND_net), .I1(n7497[15]), .I2(GND_net), 
            .I3(n23146), .O(n7475[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4401), 
            .I3(GND_net), .O(n8_adj_4417));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3512_9 (.CI(n23380), .I0(n7794[6]), .I1(n594_adj_4349), 
            .CO(n23381));
    SB_CARRY mult_11_add_1225_16 (.CI(n23345), .I0(n7725[13]), .I1(n1096_adj_4333), 
            .CO(n23346));
    SB_CARRY add_3490_18 (.CI(n23146), .I0(n7497[15]), .I1(GND_net), .CO(n23147));
    SB_LUT4 add_3490_17_lut (.I0(GND_net), .I1(n7497[14]), .I2(GND_net), 
            .I3(n23145), .O(n7475[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n7725[9]), .I2(n804_adj_4351), 
            .I3(n23341), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n7725[13]), .I2(n1096_adj_4333), 
            .I3(n23345), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n7725[19]), .I2(GND_net), 
            .I3(n23351), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_4 (.CI(n23355), .I0(n7772[1]), .I1(n226_adj_4348), 
            .CO(n23356));
    SB_CARRY mult_11_add_1225_23 (.CI(n23352), .I0(n7725[20]), .I1(GND_net), 
            .CO(n23353));
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4413), .I1(n257[22]), .I2(n45_adj_4419), 
            .I3(GND_net), .O(n24_adj_4420));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_11_add_1225_17 (.CI(n23346), .I0(n7725[14]), .I1(GND_net), 
            .CO(n23347));
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n7725[20]), .I2(GND_net), 
            .I3(n23352), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n7725[14]), .I2(GND_net), 
            .I3(n23346), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n23342), .I0(n7725[10]), .I1(n877_adj_4332), 
            .CO(n23343));
    SB_CARRY mult_11_add_1225_18 (.CI(n23347), .I0(n7725[15]), .I1(GND_net), 
            .CO(n23348));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n7725[21]), 
            .I2(GND_net), .I3(n23353), .O(n29838)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n7725[15]), .I2(GND_net), 
            .I3(n23347), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n7725[10]), .I2(n877_adj_4332), 
            .I3(n23342), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n23348), .I0(n7725[16]), .I1(GND_net), 
            .CO(n23349));
    SB_CARRY mult_11_add_1225_14 (.CI(n23343), .I0(n7725[11]), .I1(n950_adj_4350), 
            .CO(n23344));
    SB_LUT4 mux_614_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3490_17 (.CI(n23145), .I0(n7497[14]), .I1(GND_net), .CO(n23146));
    SB_LUT4 add_3490_16_lut (.I0(GND_net), .I1(n7497[13]), .I2(n1105_adj_4330), 
            .I3(n23144), .O(n7475[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_16 (.CI(n23144), .I0(n7497[13]), .I1(n1105_adj_4330), 
            .CO(n23145));
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4395));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3490_15_lut (.I0(GND_net), .I1(n7497[12]), .I2(n1032_adj_4329), 
            .I3(n23143), .O(n7475[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_9 (.CI(n22519), .I0(n2908[7]), .I1(n2933[7]), .CO(n22520));
    SB_CARRY add_3490_15 (.CI(n23143), .I0(n7497[12]), .I1(n1032_adj_4329), 
            .CO(n23144));
    SB_LUT4 add_3490_14_lut (.I0(GND_net), .I1(n7497[11]), .I2(n959_adj_4328), 
            .I3(n23142), .O(n7475[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n22466), .I0(motor_state[1]), .I1(n1[1]), 
            .CO(n22467));
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[18]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4391));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4390));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3490_14 (.CI(n23142), .I0(n7497[11]), .I1(n959_adj_4328), 
            .CO(n23143));
    SB_LUT4 i24056_4_lut (.I0(n43_adj_4412), .I1(n25_adj_4408), .I2(n23_adj_4409), 
            .I3(n29928), .O(n29908));
    defparam i24056_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3490_13_lut (.I0(GND_net), .I1(n7497[10]), .I2(n886_adj_4327), 
            .I3(n23141), .O(n7475[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_4 (.CI(n23375), .I0(n7794[1]), .I1(n229_adj_4326), 
            .CO(n23376));
    SB_CARRY add_3490_13 (.CI(n23141), .I0(n7497[10]), .I1(n886_adj_4327), 
            .CO(n23142));
    SB_LUT4 add_3490_12_lut (.I0(GND_net), .I1(n7497[9]), .I2(n813_adj_4325), 
            .I3(n23140), .O(n7475[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[13]), 
            .I3(n22594), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_12 (.CI(n23140), .I0(n7497[9]), .I1(n813_adj_4325), 
            .CO(n23141));
    SB_LUT4 add_3490_11_lut (.I0(GND_net), .I1(n7497[8]), .I2(n740), .I3(n23139), 
            .O(n7475[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_11 (.CI(n23139), .I0(n7497[8]), .I1(n740), .CO(n23140));
    SB_LUT4 add_3490_10_lut (.I0(GND_net), .I1(n7497[7]), .I2(n667), .I3(n23138), 
            .O(n7475[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3490_10 (.CI(n23138), .I0(n7497[7]), .I1(n667), .CO(n23139));
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3490_9_lut (.I0(GND_net), .I1(n7497[6]), .I2(n594), .I3(n23137), 
            .O(n7475[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n22594), .I0(GND_net), .I1(n1_adj_4607[13]), 
            .CO(n22595));
    SB_CARRY add_3490_9 (.CI(n23137), .I0(n7497[6]), .I1(n594), .CO(n23138));
    SB_LUT4 add_3490_8_lut (.I0(GND_net), .I1(n7497[5]), .I2(n521_adj_4323), 
            .I3(n23136), .O(n7475[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_8 (.CI(n23136), .I0(n7497[5]), .I1(n521_adj_4323), 
            .CO(n23137));
    SB_LUT4 add_3490_7_lut (.I0(GND_net), .I1(n7497[4]), .I2(n448), .I3(n23135), 
            .O(n7475[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_7 (.CI(n23135), .I0(n7497[4]), .I1(n448), .CO(n23136));
    SB_LUT4 add_3490_6_lut (.I0(GND_net), .I1(n7497[3]), .I2(n375), .I3(n23134), 
            .O(n7475[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4389));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3490_6 (.CI(n23134), .I0(n7497[3]), .I1(n375), .CO(n23135));
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_616_8_lut (.I0(GND_net), .I1(n2908[6]), .I2(n2933[6]), 
            .I3(n22518), .O(duty_23__N_3655[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3490_5_lut (.I0(GND_net), .I1(n7497[2]), .I2(n302), .I3(n23133), 
            .O(n7475[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_5 (.CI(n23133), .I0(n7497[2]), .I1(n302), .CO(n23134));
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4422));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3490_4_lut (.I0(GND_net), .I1(n7497[1]), .I2(n229), .I3(n23132), 
            .O(n7475[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_4 (.CI(n23132), .I0(n7497[1]), .I1(n229), .CO(n23133));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3556 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3490_3_lut (.I0(GND_net), .I1(n7497[0]), .I2(n156_adj_4321), 
            .I3(n23131), .O(n7475[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3490_3 (.CI(n23131), .I0(n7497[0]), .I1(n156_adj_4321), 
            .CO(n23132));
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4423));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4424));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4425));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4426));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24496_4_lut (.I0(n24_adj_4420), .I1(n8_adj_4417), .I2(n45_adj_4419), 
            .I3(n29906), .O(n30349));   // verilog/motorControl.v(38[19:35])
    defparam i24496_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3490_2_lut (.I0(GND_net), .I1(n14_adj_4320), .I2(n83), 
            .I3(GND_net), .O(n7475[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3490_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4427));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3526_5_lut (.I0(GND_net), .I1(n7997[2]), .I2(n344_adj_4319), 
            .I3(n23551), .O(n7989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3526_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4428));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3526_4 (.CI(n23550), .I0(n7997[1]), .I1(n271_adj_4318), 
            .CO(n23551));
    SB_CARRY add_3526_6 (.CI(n23552), .I0(n7997[3]), .I1(n417_adj_4334), 
            .CO(n23553));
    SB_LUT4 add_3526_4_lut (.I0(GND_net), .I1(n7997[1]), .I2(n271_adj_4318), 
            .I3(n23550), .O(n7989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3526_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3526_5 (.CI(n23551), .I0(n7997[2]), .I1(n344_adj_4319), 
            .CO(n23552));
    SB_CARRY add_3490_2 (.CI(GND_net), .I0(n14_adj_4320), .I1(n83), .CO(n23131));
    SB_LUT4 add_3489_22_lut (.I0(GND_net), .I1(n7475[19]), .I2(GND_net), 
            .I3(n23130), .O(n7452[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_8 (.CI(n22518), .I0(n2908[6]), .I1(n2933[6]), .CO(n22519));
    SB_LUT4 add_3489_21_lut (.I0(GND_net), .I1(n7475[18]), .I2(GND_net), 
            .I3(n23129), .O(n7452[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_21 (.CI(n23129), .I0(n7475[18]), .I1(GND_net), .CO(n23130));
    SB_LUT4 add_3489_20_lut (.I0(GND_net), .I1(n7475[17]), .I2(GND_net), 
            .I3(n23128), .O(n7452[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_19 (.CI(n23370), .I0(n7772[16]), .I1(GND_net), .CO(n23371));
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4429));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3489_20 (.CI(n23128), .I0(n7475[17]), .I1(GND_net), .CO(n23129));
    SB_LUT4 add_3489_19_lut (.I0(GND_net), .I1(n7475[16]), .I2(GND_net), 
            .I3(n23127), .O(n7452[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_19 (.CI(n23127), .I0(n7475[16]), .I1(GND_net), .CO(n23128));
    SB_LUT4 add_3526_2_lut (.I0(GND_net), .I1(n56_adj_4317), .I2(n125_adj_4316), 
            .I3(GND_net), .O(n7989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3526_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3526_3 (.CI(n23549), .I0(n7997[0]), .I1(n198_adj_4315), 
            .CO(n23550));
    SB_LUT4 add_3526_3_lut (.I0(GND_net), .I1(n7997[0]), .I2(n198_adj_4315), 
            .I3(n23549), .O(n7989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3526_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3489_18_lut (.I0(GND_net), .I1(n7475[15]), .I2(GND_net), 
            .I3(n23126), .O(n7452[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4430));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4431));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3489_18 (.CI(n23126), .I0(n7475[15]), .I1(GND_net), .CO(n23127));
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1[0]), 
            .CO(n22466));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[12]), 
            .I3(n22593), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3489_17_lut (.I0(GND_net), .I1(n7475[14]), .I2(GND_net), 
            .I3(n23125), .O(n7452[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_17 (.CI(n23125), .I0(n7475[14]), .I1(GND_net), .CO(n23126));
    SB_CARRY add_3526_2 (.CI(GND_net), .I0(n56_adj_4317), .I1(n125_adj_4316), 
            .CO(n23549));
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4432));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3524_7 (.CI(n23540), .I0(n7980[4]), .I1(n484_adj_4313), 
            .CO(n23541));
    SB_LUT4 add_3524_7_lut (.I0(GND_net), .I1(n7980[4]), .I2(n484_adj_4313), 
            .I3(n23540), .O(n7970[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3524_5 (.CI(n23538), .I0(n7980[2]), .I1(n338_adj_4312), 
            .CO(n23539));
    SB_LUT4 add_3524_8_lut (.I0(GND_net), .I1(n7980[5]), .I2(n557_adj_4311), 
            .I3(n23541), .O(n7970[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3524_5_lut (.I0(GND_net), .I1(n7980[2]), .I2(n338_adj_4312), 
            .I3(n23538), .O(n7970[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3524_6 (.CI(n23539), .I0(n7980[3]), .I1(n411_adj_4310), 
            .CO(n23540));
    SB_LUT4 add_616_7_lut (.I0(GND_net), .I1(n2908[5]), .I2(n2933[5]), 
            .I3(n22517), .O(duty_23__N_3655[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3525_6 (.CI(n23546), .I0(n7989[3]), .I1(n414_adj_4309), 
            .CO(n23547));
    SB_LUT4 add_3525_4_lut (.I0(GND_net), .I1(n7989[1]), .I2(n268_adj_4308), 
            .I3(n23544), .O(n7980[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3525_5 (.CI(n23545), .I0(n7989[2]), .I1(n341_adj_4307), 
            .CO(n23546));
    SB_LUT4 add_3489_16_lut (.I0(GND_net), .I1(n7475[13]), .I2(n1102), 
            .I3(n23124), .O(n7452[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3525_7_lut (.I0(GND_net), .I1(n7989[4]), .I2(n487_adj_4306), 
            .I3(n23547), .O(n7980[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4433));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3525_3 (.CI(n23543), .I0(n7989[0]), .I1(n195_adj_4305), 
            .CO(n23544));
    SB_CARRY add_3524_8 (.CI(n23541), .I0(n7980[5]), .I1(n557_adj_4311), 
            .CO(n23542));
    SB_LUT4 add_3524_9_lut (.I0(GND_net), .I1(n7980[6]), .I2(n630_adj_4304), 
            .I3(n23542), .O(n7970[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3524_6_lut (.I0(GND_net), .I1(n7980[3]), .I2(n411_adj_4310), 
            .I3(n23539), .O(n7970[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3525_6_lut (.I0(GND_net), .I1(n7989[3]), .I2(n414_adj_4309), 
            .I3(n23546), .O(n7980[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3525_5_lut (.I0(GND_net), .I1(n7989[2]), .I2(n341_adj_4307), 
            .I3(n23545), .O(n7980[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3525_8_lut (.I0(GND_net), .I1(n7989[5]), .I2(n560_adj_4303), 
            .I3(n23548), .O(n7980[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_16 (.CI(n23124), .I0(n7475[13]), .I1(n1102), .CO(n23125));
    SB_LUT4 add_3525_3_lut (.I0(GND_net), .I1(n7989[0]), .I2(n195_adj_4305), 
            .I3(n23543), .O(n7980[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3525_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3525_2 (.CI(GND_net), .I0(n53_adj_4356), .I1(n122_adj_4355), 
            .CO(n23543));
    SB_CARRY add_3525_7 (.CI(n23547), .I0(n7989[4]), .I1(n487_adj_4306), 
            .CO(n23548));
    SB_CARRY add_3525_4 (.CI(n23544), .I0(n7989[1]), .I1(n268_adj_4308), 
            .CO(n23545));
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4434));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3489_15_lut (.I0(GND_net), .I1(n7475[12]), .I2(n1029), 
            .I3(n23123), .O(n7452[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4435));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3489_15 (.CI(n23123), .I0(n7475[12]), .I1(n1029), .CO(n23124));
    SB_CARRY unary_minus_16_add_3_14 (.CI(n22593), .I0(GND_net), .I1(n1_adj_4607[12]), 
            .CO(n22594));
    SB_LUT4 add_3489_14_lut (.I0(GND_net), .I1(n7475[11]), .I2(n956), 
            .I3(n23122), .O(n7452[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4436));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4178));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3489_14 (.CI(n23122), .I0(n7475[11]), .I1(n956), .CO(n23123));
    SB_LUT4 add_3489_13_lut (.I0(GND_net), .I1(n7475[10]), .I2(n883), 
            .I3(n23121), .O(n7452[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_13 (.CI(n23121), .I0(n7475[10]), .I1(n883), .CO(n23122));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[11]), 
            .I3(n22592), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3489_12_lut (.I0(GND_net), .I1(n7475[9]), .I2(n810), .I3(n23120), 
            .O(n7452[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_7 (.CI(n22517), .I0(n2908[5]), .I1(n2933[5]), .CO(n22518));
    SB_CARRY add_3489_12 (.CI(n23120), .I0(n7475[9]), .I1(n810), .CO(n23121));
    SB_LUT4 add_3489_11_lut (.I0(GND_net), .I1(n7475[8]), .I2(n737_adj_4301), 
            .I3(n23119), .O(n7452[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4437));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3489_11 (.CI(n23119), .I0(n7475[8]), .I1(n737_adj_4301), 
            .CO(n23120));
    SB_LUT4 add_3489_10_lut (.I0(GND_net), .I1(n7475[7]), .I2(n664_adj_4300), 
            .I3(n23118), .O(n7452[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_10 (.CI(n23118), .I0(n7475[7]), .I1(n664_adj_4300), 
            .CO(n23119));
    SB_LUT4 add_3489_9_lut (.I0(GND_net), .I1(n7475[6]), .I2(n591_adj_4299), 
            .I3(n23117), .O(n7452[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4438));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3489_9 (.CI(n23117), .I0(n7475[6]), .I1(n591_adj_4299), 
            .CO(n23118));
    SB_LUT4 add_3489_8_lut (.I0(GND_net), .I1(n7475[5]), .I2(n518), .I3(n23116), 
            .O(n7452[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_8 (.CI(n23116), .I0(n7475[5]), .I1(n518), .CO(n23117));
    SB_LUT4 add_3489_7_lut (.I0(GND_net), .I1(n7475[4]), .I2(n445), .I3(n23115), 
            .O(n7452[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_7 (.CI(n23115), .I0(n7475[4]), .I1(n445), .CO(n23116));
    SB_LUT4 add_3489_6_lut (.I0(GND_net), .I1(n7475[3]), .I2(n372), .I3(n23114), 
            .O(n7452[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3489_6 (.CI(n23114), .I0(n7475[3]), .I1(n372), .CO(n23115));
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4439));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4440));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3489_5_lut (.I0(GND_net), .I1(n7475[2]), .I2(n299), .I3(n23113), 
            .O(n7452[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24113_4_lut (.I0(n21_adj_4440), .I1(n19_adj_4439), .I2(n17_adj_4438), 
            .I3(n9_adj_4437), .O(n29965));
    defparam i24113_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24567_3_lut (.I0(n30447), .I1(n257[12]), .I2(n25_adj_4408), 
            .I3(GND_net), .O(n30420));   // verilog/motorControl.v(38[19:35])
    defparam i24567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24104_4_lut (.I0(n27_adj_4436), .I1(n15_adj_4435), .I2(n13_adj_4434), 
            .I3(n11_adj_4433), .O(n29956));
    defparam i24104_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3489_5 (.CI(n23113), .I0(n7475[2]), .I1(n299), .CO(n23114));
    SB_LUT4 add_3489_4_lut (.I0(GND_net), .I1(n7475[1]), .I2(n226), .I3(n23112), 
            .O(n7452[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3489_4 (.CI(n23112), .I0(n7475[1]), .I1(n226), .CO(n23113));
    SB_LUT4 add_3489_3_lut (.I0(GND_net), .I1(n7475[0]), .I2(n153), .I3(n23111), 
            .O(n7452[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_4441), .I1(duty[17]), .I2(n35_adj_4431), 
            .I3(GND_net), .O(n30_adj_4442));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n29828), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_4443));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24376_4_lut (.I0(n13_adj_4434), .I1(n11_adj_4433), .I2(n9_adj_4437), 
            .I3(n29975), .O(n30229));
    defparam i24376_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24372_4_lut (.I0(n19_adj_4439), .I1(n17_adj_4438), .I2(n15_adj_4435), 
            .I3(n30229), .O(n30225));
    defparam i24372_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24631_4_lut (.I0(n25_adj_4428), .I1(n23_adj_4427), .I2(n21_adj_4440), 
            .I3(n30225), .O(n30484));
    defparam i24631_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24488_4_lut (.I0(n31_adj_4430), .I1(n29_adj_4429), .I2(n27_adj_4436), 
            .I3(n30484), .O(n30341));
    defparam i24488_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24655_4_lut (.I0(n37_adj_4425), .I1(n35_adj_4431), .I2(n33_adj_4432), 
            .I3(n30341), .O(n30508));
    defparam i24655_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24609_3_lut (.I0(n6_adj_4444), .I1(duty[10]), .I2(n21_adj_4440), 
            .I3(GND_net), .O(n30462));   // verilog/motorControl.v(36[10:25])
    defparam i24609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24610_3_lut (.I0(n30462), .I1(duty[11]), .I2(n23_adj_4427), 
            .I3(GND_net), .O(n30463));   // verilog/motorControl.v(36[10:25])
    defparam i24610_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3489_3 (.CI(n23111), .I0(n7475[0]), .I1(n153), .CO(n23112));
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1485 (.I0(n6_adj_4445), .I1(\Kp[4] ), .I2(n7707[2]), 
            .I3(\PID_CONTROLLER.err [18]), .O(n7700[3]));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1485.LUT_INIT = 16'h965a;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_4446), .I1(duty[22]), .I2(n45_adj_4424), 
            .I3(GND_net), .O(n24_adj_4447));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24090_4_lut (.I0(n43_adj_4426), .I1(n25_adj_4428), .I2(n23_adj_4427), 
            .I3(n29965), .O(n29942));
    defparam i24090_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3489_2_lut (.I0(GND_net), .I1(n11_adj_4298), .I2(n80), 
            .I3(GND_net), .O(n7452[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3489_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24494_4_lut (.I0(n24_adj_4447), .I1(n8_adj_4448), .I2(n45_adj_4424), 
            .I3(n29940), .O(n30347));   // verilog/motorControl.v(36[10:25])
    defparam i24494_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3489_2 (.CI(GND_net), .I0(n11_adj_4298), .I1(n80), .CO(n23111));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n7428[21]), 
            .I2(GND_net), .I3(n23110), .O(n5869[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3524_4_lut (.I0(GND_net), .I1(n7980[1]), .I2(n265_adj_4297), 
            .I3(n23537), .O(n7970[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n18939), .I1(n7428[20]), .I2(GND_net), 
            .I3(n23109), .O(n2908[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_23 (.CI(n23109), .I0(n7428[20]), .I1(GND_net), 
            .CO(n23110));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n18939), .I1(n7428[19]), .I2(GND_net), 
            .I3(n23108), .O(n2908[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n22592), .I0(GND_net), .I1(n1_adj_4607[11]), 
            .CO(n22593));
    SB_LUT4 i24561_3_lut (.I0(n30463), .I1(duty[12]), .I2(n25_adj_4428), 
            .I3(GND_net), .O(n30414));   // verilog/motorControl.v(36[10:25])
    defparam i24561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4449));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i24597_3_lut (.I0(n4_adj_4449), .I1(duty[13]), .I2(n27_adj_4436), 
            .I3(GND_net), .O(n30450));   // verilog/motorControl.v(36[10:25])
    defparam i24597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24591_3_lut (.I0(n4_adj_4443), .I1(n257[13]), .I2(n27_adj_4381), 
            .I3(GND_net), .O(n30444));   // verilog/motorControl.v(38[19:35])
    defparam i24591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[10]), 
            .I3(n22591), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_6_lut (.I0(GND_net), .I1(n2908[4]), .I2(n2933[4]), 
            .I3(n22516), .O(duty_23__N_3655[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n23108), .I0(n7428[19]), .I1(GND_net), 
            .CO(n23109));
    SB_LUT4 i24598_3_lut (.I0(n30450), .I1(duty[14]), .I2(n29_adj_4429), 
            .I3(GND_net), .O(n30451));   // verilog/motorControl.v(36[10:25])
    defparam i24598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24100_4_lut (.I0(n33_adj_4432), .I1(n31_adj_4430), .I2(n29_adj_4429), 
            .I3(n29956), .O(n29952));
    defparam i24100_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n22591), .I0(GND_net), .I1(n1_adj_4607[10]), 
            .CO(n22592));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[9]), 
            .I3(n22590), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24665_4_lut (.I0(n30_adj_4442), .I1(n10_adj_4450), .I2(n35_adj_4431), 
            .I3(n29950), .O(n30518));   // verilog/motorControl.v(36[10:25])
    defparam i24665_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n22590), .I0(GND_net), .I1(n1_adj_4607[9]), 
            .CO(n22591));
    SB_LUT4 i24563_3_lut (.I0(n30451), .I1(duty[15]), .I2(n31_adj_4430), 
            .I3(GND_net), .O(n30416));   // verilog/motorControl.v(36[10:25])
    defparam i24563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17579_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n7718[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17579_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1486 (.I0(n4_adj_4451), .I1(\Kp[3] ), .I2(n7713[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n7707[2]));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1486.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24592_3_lut (.I0(n30444), .I1(n257[14]), .I2(n29_adj_4410), 
            .I3(GND_net), .O(n30445));   // verilog/motorControl.v(38[19:35])
    defparam i24592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[8]), 
            .I3(n22589), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1487 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_4452));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1487.LUT_INIT = 16'h9c50;
    SB_LUT4 i17515_4_lut (.I0(n7707[2]), .I1(\Kp[4] ), .I2(n6_adj_4445), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_4453));   // verilog/motorControl.v(34[17:23])
    defparam i17515_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1488 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_4454));   // verilog/motorControl.v(34[17:23])
    defparam i1_4_lut_adj_1488.LUT_INIT = 16'h6ca0;
    SB_LUT4 i24701_4_lut (.I0(n30416), .I1(n30518), .I2(n35_adj_4431), 
            .I3(n29952), .O(n30554));   // verilog/motorControl.v(36[10:25])
    defparam i24701_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i17546_4_lut (.I0(n7713[1]), .I1(\Kp[3] ), .I2(n4_adj_4451), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_4455));   // verilog/motorControl.v(34[17:23])
    defparam i17546_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i17581_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n22128));   // verilog/motorControl.v(34[17:23])
    defparam i17581_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1489 (.I0(n6_adj_4455), .I1(n11_adj_4454), .I2(n8_adj_4453), 
            .I3(n12_adj_4452), .O(n18_adj_4456));   // verilog/motorControl.v(34[17:23])
    defparam i8_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 add_3512_4_lut (.I0(GND_net), .I1(n7794[1]), .I2(n229_adj_4326), 
            .I3(n23375), .O(n7772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_6 (.CI(n22516), .I0(n2908[4]), .I1(n2933[4]), .CO(n22517));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n22589), .I0(GND_net), .I1(n1_adj_4607[8]), 
            .CO(n22590));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[7]), 
            .I3(n22588), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n22588), .I0(GND_net), .I1(n1_adj_4607[7]), 
            .CO(n22589));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[6]), 
            .I3(n22587), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_5_lut (.I0(GND_net), .I1(n2908[3]), .I2(n2933[3]), 
            .I3(n22515), .O(duty_23__N_3655[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n18939), .I1(n7428[18]), .I2(GND_net), 
            .I3(n23107), .O(n2908[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_616_5 (.CI(n22515), .I0(n2908[3]), .I1(n2933[3]), .CO(n22516));
    SB_LUT4 i24702_3_lut (.I0(n30554), .I1(duty[18]), .I2(n37_adj_4425), 
            .I3(GND_net), .O(n30555));   // verilog/motorControl.v(36[10:25])
    defparam i24702_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_10_add_1225_21 (.CI(n23107), .I0(n7428[18]), .I1(GND_net), 
            .CO(n23108));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n18939), .I1(n7428[17]), .I2(GND_net), 
            .I3(n23106), .O(n2908[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i24688_3_lut (.I0(n30555), .I1(duty[19]), .I2(n39_adj_4422), 
            .I3(GND_net), .O(n30541));   // verilog/motorControl.v(36[10:25])
    defparam i24688_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_10_add_1225_20 (.CI(n23106), .I0(n7428[17]), .I1(GND_net), 
            .CO(n23107));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n18939), .I1(n7428[16]), .I2(GND_net), 
            .I3(n23105), .O(n2908[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i24092_4_lut (.I0(n43_adj_4426), .I1(n41_adj_4423), .I2(n39_adj_4422), 
            .I3(n30508), .O(n29944));
    defparam i24092_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24621_4_lut (.I0(n30414), .I1(n30347), .I2(n45_adj_4424), 
            .I3(n29942), .O(n30474));   // verilog/motorControl.v(36[10:25])
    defparam i24621_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24678_3_lut (.I0(n30541), .I1(duty[20]), .I2(n41_adj_4423), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(36[10:25])
    defparam i24678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24623_4_lut (.I0(n40), .I1(n30474), .I2(n45_adj_4424), .I3(n29944), 
            .O(n30476));   // verilog/motorControl.v(36[10:25])
    defparam i24623_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24624_3_lut (.I0(n30476), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3679));   // verilog/motorControl.v(36[10:25])
    defparam i24624_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3655[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3511_9 (.CI(n23360), .I0(n7772[6]), .I1(n591), .CO(n23361));
    SB_LUT4 add_3511_9_lut (.I0(GND_net), .I1(n7772[6]), .I2(n591), .I3(n23360), 
            .O(n7749[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_10 (.CI(n23361), .I0(n7772[7]), .I1(n664), .CO(n23362));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n22587), .I0(GND_net), .I1(n1_adj_4607[6]), 
            .CO(n22588));
    SB_LUT4 add_3511_10_lut (.I0(GND_net), .I1(n7772[7]), .I2(n664), .I3(n23361), 
            .O(n7749[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_616_4_lut (.I0(GND_net), .I1(n2908[2]), .I2(n2933[2]), 
            .I3(n22514), .O(duty_23__N_3655[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3511_11 (.CI(n23362), .I0(n7772[8]), .I1(n737), .CO(n23363));
    SB_LUT4 add_3511_11_lut (.I0(GND_net), .I1(n7772[8]), .I2(n737), .I3(n23362), 
            .O(n7749[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24066_4_lut (.I0(n33_adj_4353), .I1(n31_adj_4331), .I2(n29_adj_4410), 
            .I3(n29922), .O(n29918));
    defparam i24066_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[5]), 
            .I3(n22586), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n23105), .I0(n7428[16]), .I1(GND_net), 
            .CO(n23106));
    SB_CARRY unary_minus_16_add_3_7 (.CI(n22586), .I0(GND_net), .I1(n1_adj_4607[5]), 
            .CO(n22587));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n18939), .I1(n7428[15]), .I2(GND_net), 
            .I3(n23104), .O(n2908[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_18 (.CI(n23104), .I0(n7428[15]), .I1(GND_net), 
            .CO(n23105));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n18939), .I1(n7428[14]), .I2(GND_net), 
            .I3(n23103), .O(n2908[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_17 (.CI(n23103), .I0(n7428[14]), .I1(GND_net), 
            .CO(n23104));
    SB_LUT4 add_3511_18_lut (.I0(GND_net), .I1(n7772[15]), .I2(GND_net), 
            .I3(n23369), .O(n7749[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3511_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4387));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[4]), 
            .I3(n22585), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_616_4 (.CI(n22514), .I0(n2908[2]), .I1(n2933[2]), .CO(n22515));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n18939), .I1(n7428[13]), .I2(n1096), 
            .I3(n23102), .O(n2908[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_16 (.CI(n23102), .I0(n7428[13]), .I1(n1096), 
            .CO(n23103));
    SB_LUT4 add_3512_3_lut (.I0(GND_net), .I1(n7794[0]), .I2(n156), .I3(n23374), 
            .O(n7772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3512_8_lut (.I0(GND_net), .I1(n7794[5]), .I2(n521), .I3(n23379), 
            .O(n7772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n18939), .I1(n7428[12]), .I2(n1023), 
            .I3(n23101), .O(n2908[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_15 (.CI(n23101), .I0(n7428[12]), .I1(n1023), 
            .CO(n23102));
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n18939), .I1(n7428[11]), .I2(n950), 
            .I3(n23100), .O(n2908[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_14 (.CI(n23100), .I0(n7428[11]), .I1(n950), 
            .CO(n23101));
    SB_CARRY add_3512_3 (.CI(n23374), .I0(n7794[0]), .I1(n156), .CO(n23375));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n18939), .I1(n7428[10]), .I2(n877), 
            .I3(n23099), .O(n2908[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_13 (.CI(n23099), .I0(n7428[10]), .I1(n877), 
            .CO(n23100));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n18939), .I1(n7428[9]), .I2(n804), 
            .I3(n23098), .O(n2908[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_12 (.CI(n23098), .I0(n7428[9]), .I1(n804), 
            .CO(n23099));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n18939), .I1(n7428[8]), .I2(n731), 
            .I3(n23097), .O(n2908[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3512_8 (.CI(n23379), .I0(n7794[5]), .I1(n521), .CO(n23380));
    SB_CARRY mult_10_add_1225_11 (.CI(n23097), .I0(n7428[8]), .I1(n731), 
            .CO(n23098));
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n18939), .I1(n7428[7]), .I2(n658), 
            .I3(n23096), .O(n2908[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_10 (.CI(n23096), .I0(n7428[7]), .I1(n658), 
            .CO(n23097));
    SB_LUT4 i24667_4_lut (.I0(n30_adj_4407), .I1(n10_adj_4406), .I2(n35_adj_4344), 
            .I3(n29916), .O(n30520));   // verilog/motorControl.v(38[19:35])
    defparam i24667_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n18939), .I1(n7428[6]), .I2(n585_adj_4289), 
            .I3(n23095), .O(n2908[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_9 (.CI(n23095), .I0(n7428[6]), .I1(n585_adj_4289), 
            .CO(n23096));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n18939), .I1(n7428[5]), .I2(n512_adj_4288), 
            .I3(n23094), .O(n2908[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_8 (.CI(n23094), .I0(n7428[5]), .I1(n512_adj_4288), 
            .CO(n23095));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n18939), .I1(n7428[4]), .I2(n439_adj_4287), 
            .I3(n23093), .O(n2908[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_7 (.CI(n23093), .I0(n7428[4]), .I1(n439_adj_4287), 
            .CO(n23094));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n18939), .I1(n7428[3]), .I2(n366_adj_4286), 
            .I3(n23092), .O(n2908[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_6 (.CI(n23092), .I0(n7428[3]), .I1(n366_adj_4286), 
            .CO(n23093));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n18939), .I1(n7428[2]), .I2(n293_adj_4285), 
            .I3(n23091), .O(n2908[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_5 (.CI(n23091), .I0(n7428[2]), .I1(n293_adj_4285), 
            .CO(n23092));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n18939), .I1(n7428[1]), .I2(n220_adj_4284), 
            .I3(n23090), .O(n2908[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_4 (.CI(n23090), .I0(n7428[1]), .I1(n220_adj_4284), 
            .CO(n23091));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n18939), .I1(n7428[0]), .I2(n147_adj_4283), 
            .I3(n23089), .O(n2908[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_3 (.CI(n23089), .I0(n7428[0]), .I1(n147_adj_4283), 
            .CO(n23090));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n18939), .I1(n5_adj_4282), .I2(n74_adj_4281), 
            .I3(GND_net), .O(n2908[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4282), .I1(n74_adj_4281), 
            .CO(n23089));
    SB_LUT4 add_616_3_lut (.I0(GND_net), .I1(n2908[1]), .I2(n2933[1]), 
            .I3(n22513), .O(duty_23__N_3655[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n22585), .I0(GND_net), .I1(n1_adj_4607[4]), 
            .CO(n22586));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[3]), 
            .I3(n22584), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3488_23_lut (.I0(GND_net), .I1(n7452[20]), .I2(GND_net), 
            .I3(n23088), .O(n7428[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3488_22_lut (.I0(GND_net), .I1(n7452[19]), .I2(GND_net), 
            .I3(n23087), .O(n7428[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_22 (.CI(n23087), .I0(n7452[19]), .I1(GND_net), .CO(n23088));
    SB_LUT4 add_3488_21_lut (.I0(GND_net), .I1(n7452[18]), .I2(GND_net), 
            .I3(n23086), .O(n7428[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n22584), .I0(GND_net), .I1(n1_adj_4607[3]), 
            .CO(n22585));
    SB_CARRY add_3488_21 (.CI(n23086), .I0(n7452[18]), .I1(GND_net), .CO(n23087));
    SB_LUT4 add_3488_20_lut (.I0(GND_net), .I1(n7452[17]), .I2(GND_net), 
            .I3(n23085), .O(n7428[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_20 (.CI(n23085), .I0(n7452[17]), .I1(GND_net), .CO(n23086));
    SB_LUT4 add_3488_19_lut (.I0(GND_net), .I1(n7452[16]), .I2(GND_net), 
            .I3(n23084), .O(n7428[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_19 (.CI(n23084), .I0(n7452[16]), .I1(GND_net), .CO(n23085));
    SB_LUT4 add_3488_18_lut (.I0(GND_net), .I1(n7452[15]), .I2(GND_net), 
            .I3(n23083), .O(n7428[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_18 (.CI(n23083), .I0(n7452[15]), .I1(GND_net), .CO(n23084));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[2]), 
            .I3(n22583), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3488_17_lut (.I0(GND_net), .I1(n7452[14]), .I2(GND_net), 
            .I3(n23082), .O(n7428[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_17 (.CI(n23082), .I0(n7452[14]), .I1(GND_net), .CO(n23083));
    SB_LUT4 add_3488_16_lut (.I0(GND_net), .I1(n7452[13]), .I2(n1099_adj_4278), 
            .I3(n23081), .O(n7428[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_16 (.CI(n23081), .I0(n7452[13]), .I1(n1099_adj_4278), 
            .CO(n23082));
    SB_LUT4 add_3488_15_lut (.I0(GND_net), .I1(n7452[12]), .I2(n1026_adj_4277), 
            .I3(n23080), .O(n7428[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_15 (.CI(n23080), .I0(n7452[12]), .I1(n1026_adj_4277), 
            .CO(n23081));
    SB_LUT4 add_3488_14_lut (.I0(GND_net), .I1(n7452[11]), .I2(n953_adj_4276), 
            .I3(n23079), .O(n7428[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_14 (.CI(n23079), .I0(n7452[11]), .I1(n953_adj_4276), 
            .CO(n23080));
    SB_CARRY add_616_3 (.CI(n22513), .I0(n2908[1]), .I1(n2933[1]), .CO(n22514));
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3488_13_lut (.I0(GND_net), .I1(n7452[10]), .I2(n880_adj_4275), 
            .I3(n23078), .O(n7428[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3488_13 (.CI(n23078), .I0(n7452[10]), .I1(n880_adj_4275), 
            .CO(n23079));
    SB_LUT4 i24569_3_lut (.I0(n30445), .I1(n257[15]), .I2(n31_adj_4331), 
            .I3(GND_net), .O(n30422));   // verilog/motorControl.v(38[19:35])
    defparam i24569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3488_12_lut (.I0(GND_net), .I1(n7452[9]), .I2(n807_adj_4274), 
            .I3(n23077), .O(n7428[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1490 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13_adj_4457));   // verilog/motorControl.v(34[17:23])
    defparam i3_4_lut_adj_1490.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1491 (.I0(n13_adj_4457), .I1(n18_adj_4456), .I2(n22128), 
            .I3(n4_adj_4458), .O(n28160));   // verilog/motorControl.v(34[17:23])
    defparam i9_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_CARRY add_3488_12 (.CI(n23077), .I0(n7452[9]), .I1(n807_adj_4274), 
            .CO(n23078));
    SB_LUT4 add_3488_11_lut (.I0(GND_net), .I1(n7452[8]), .I2(n734_adj_4273), 
            .I3(n23076), .O(n7428[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_11 (.CI(n23076), .I0(n7452[8]), .I1(n734_adj_4273), 
            .CO(n23077));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3488_10_lut (.I0(GND_net), .I1(n7452[7]), .I2(n661_adj_4272), 
            .I3(n23075), .O(n7428[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_10 (.CI(n23075), .I0(n7452[7]), .I1(n661_adj_4272), 
            .CO(n23076));
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3488_9_lut (.I0(GND_net), .I1(n7452[6]), .I2(n588_adj_4271), 
            .I3(n23074), .O(n7428[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4385));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i13_3_lut (.I0(n155[12]), .I1(PWMLimit[12]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3488_9 (.CI(n23074), .I0(n7452[6]), .I1(n588_adj_4271), 
            .CO(n23075));
    SB_LUT4 add_3488_8_lut (.I0(GND_net), .I1(n7452[5]), .I2(n515_adj_4270), 
            .I3(n23073), .O(n7428[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_8 (.CI(n23073), .I0(n7452[5]), .I1(n515_adj_4270), 
            .CO(n23074));
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[19]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3488_7_lut (.I0(GND_net), .I1(n7452[4]), .I2(n442_adj_4269), 
            .I3(n23072), .O(n7428[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_7 (.CI(n23072), .I0(n7452[4]), .I1(n442_adj_4269), 
            .CO(n23073));
    SB_LUT4 add_3488_6_lut (.I0(GND_net), .I1(n7452[3]), .I2(n369_adj_4268), 
            .I3(n23071), .O(n7428[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3488_6 (.CI(n23071), .I0(n7452[3]), .I1(n369_adj_4268), 
            .CO(n23072));
    SB_LUT4 add_3488_5_lut (.I0(GND_net), .I1(n7452[2]), .I2(n296_adj_4267), 
            .I3(n23070), .O(n7428[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_5 (.CI(n23070), .I0(n7452[2]), .I1(n296_adj_4267), 
            .CO(n23071));
    SB_LUT4 add_3488_4_lut (.I0(GND_net), .I1(n7452[1]), .I2(n223_adj_4266), 
            .I3(n23069), .O(n7428[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_4 (.CI(n23069), .I0(n7452[1]), .I1(n223_adj_4266), 
            .CO(n23070));
    SB_LUT4 add_3488_3_lut (.I0(GND_net), .I1(n7452[0]), .I2(n150_adj_4265), 
            .I3(n23068), .O(n7428[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_3 (.CI(n23068), .I0(n7452[0]), .I1(n150_adj_4265), 
            .CO(n23069));
    SB_LUT4 add_3488_2_lut (.I0(GND_net), .I1(n8_adj_4264), .I2(n77_adj_4263), 
            .I3(GND_net), .O(n7428[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3488_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3488_2 (.CI(GND_net), .I0(n8_adj_4264), .I1(n77_adj_4263), 
            .CO(n23068));
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4373));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_616_2_lut (.I0(GND_net), .I1(n2908[0]), .I2(n2933[0]), 
            .I3(GND_net), .O(duty_23__N_3655[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_616_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24703_4_lut (.I0(n30422), .I1(n30520), .I2(n35_adj_4344), 
            .I3(n29918), .O(n30556));   // verilog/motorControl.v(38[19:35])
    defparam i24703_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n22583), .I0(GND_net), .I1(n1_adj_4607[2]), 
            .CO(n22584));
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4607[1]), 
            .I3(n22582), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n22582), .I0(GND_net), .I1(n1_adj_4607[1]), 
            .CO(n22583));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1_adj_4607[0]), 
            .I3(VCC_net), .O(n29828)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4607[0]), 
            .CO(n22582));
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_616_2 (.CI(GND_net), .I0(n2908[0]), .I1(n2933[0]), .CO(n22513));
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4606[23]), 
            .I3(n22581), .O(\PID_CONTROLLER.integral_23__N_3631 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4606[22]), .I3(n22580), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n22580), .I0(GND_net), .I1(n1_adj_4606[22]), 
            .CO(n22581));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4606[21]), .I3(n22579), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n22579), .I0(GND_net), .I1(n1_adj_4606[21]), 
            .CO(n22580));
    SB_LUT4 i24704_3_lut (.I0(n30556), .I1(n257[18]), .I2(n37_adj_4411), 
            .I3(GND_net), .O(n30557));   // verilog/motorControl.v(38[19:35])
    defparam i24704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4606[20]), .I3(n22578), .O(n41_adj_4212)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n22578), .I0(GND_net), .I1(n1_adj_4606[20]), 
            .CO(n22579));
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3524_4 (.CI(n23537), .I0(n7980[1]), .I1(n265_adj_4297), 
            .CO(n23538));
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4245));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4606[19]), .I3(n22577), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3524_3 (.CI(n23536), .I0(n7980[0]), .I1(n192_adj_4354), 
            .CO(n23537));
    SB_CARRY add_3524_2 (.CI(GND_net), .I0(n50_adj_4255), .I1(n119_adj_4254), 
            .CO(n23536));
    SB_LUT4 add_3523_9_lut (.I0(GND_net), .I1(n7970[6]), .I2(n627_adj_4253), 
            .I3(n23534), .O(n7959[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n22577), .I0(GND_net), .I1(n1_adj_4606[19]), 
            .CO(n22578));
    SB_LUT4 add_3523_8_lut (.I0(GND_net), .I1(n7970[5]), .I2(n554_adj_4252), 
            .I3(n23533), .O(n7959[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4606[18]), .I3(n22576), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n22576), .I0(GND_net), .I1(n1_adj_4606[18]), 
            .CO(n22577));
    SB_LUT4 mux_614_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i24686_3_lut (.I0(n30557), .I1(n257[19]), .I2(n39_adj_4460), 
            .I3(GND_net), .O(n30539));   // verilog/motorControl.v(38[19:35])
    defparam i24686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24058_4_lut (.I0(n43_adj_4412), .I1(n41_adj_4461), .I2(n39_adj_4460), 
            .I3(n30506), .O(n29910));
    defparam i24058_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4606[17]), .I3(n22575), .O(n35_adj_4197)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n22575), .I0(GND_net), .I1(n1_adj_4606[17]), 
            .CO(n22576));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4606[16]), .I3(n22574), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n22574), .I0(GND_net), .I1(n1_adj_4606[16]), 
            .CO(n22575));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4606[15]), .I3(n22573), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24627_4_lut (.I0(n30420), .I1(n30349), .I2(n45_adj_4419), 
            .I3(n29908), .O(n30480));   // verilog/motorControl.v(38[19:35])
    defparam i24627_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24680_3_lut (.I0(n30539), .I1(n257[20]), .I2(n41_adj_4461), 
            .I3(GND_net), .O(n40_adj_4462));   // verilog/motorControl.v(38[19:35])
    defparam i24680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24629_4_lut (.I0(n40_adj_4462), .I1(n30480), .I2(n45_adj_4419), 
            .I3(n29910), .O(n30482));   // verilog/motorControl.v(38[19:35])
    defparam i24629_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24630_3_lut (.I0(n30482), .I1(duty[23]), .I2(n47_adj_4180), 
            .I3(GND_net), .O(n256_adj_4200));   // verilog/motorControl.v(38[19:35])
    defparam i24630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i24_3_lut (.I0(n29838), .I1(PWMLimit[23]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14397_2_lut (.I0(n5869[0]), .I1(n256_adj_4200), .I2(GND_net), 
            .I3(GND_net), .O(n2908[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam i14397_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3523_8 (.CI(n23533), .I0(n7970[5]), .I1(n554_adj_4252), 
            .CO(n23534));
    SB_LUT4 add_3523_7_lut (.I0(GND_net), .I1(n7970[4]), .I2(n481_adj_4247), 
            .I3(n23532), .O(n7959[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3523_7 (.CI(n23532), .I0(n7970[4]), .I1(n481_adj_4247), 
            .CO(n23533));
    SB_LUT4 add_3523_6_lut (.I0(GND_net), .I1(n7970[3]), .I2(n408_adj_4246), 
            .I3(n23531), .O(n7959[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3523_6 (.CI(n23531), .I0(n7970[3]), .I1(n408_adj_4246), 
            .CO(n23532));
    SB_LUT4 add_3523_5_lut (.I0(GND_net), .I1(n7970[2]), .I2(n335_adj_4244), 
            .I3(n23530), .O(n7959[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3523_5 (.CI(n23530), .I0(n7970[2]), .I1(n335_adj_4244), 
            .CO(n23531));
    SB_LUT4 add_3523_4_lut (.I0(GND_net), .I1(n7970[1]), .I2(n262_adj_4243), 
            .I3(n23529), .O(n7959[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3523_4 (.CI(n23529), .I0(n7970[1]), .I1(n262_adj_4243), 
            .CO(n23530));
    SB_LUT4 add_3523_3_lut (.I0(GND_net), .I1(n7970[0]), .I2(n189_adj_4242), 
            .I3(n23528), .O(n7959[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3523_3 (.CI(n23528), .I0(n7970[0]), .I1(n189_adj_4242), 
            .CO(n23529));
    SB_LUT4 add_3523_2_lut (.I0(GND_net), .I1(n47_adj_4241), .I2(n116_adj_4240), 
            .I3(GND_net), .O(n7959[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3523_2 (.CI(GND_net), .I0(n47_adj_4241), .I1(n116_adj_4240), 
            .CO(n23528));
    SB_LUT4 add_3522_11_lut (.I0(GND_net), .I1(n7959[8]), .I2(n770_adj_4239), 
            .I3(n23527), .O(n7947[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3522_10_lut (.I0(GND_net), .I1(n7959[7]), .I2(n697_adj_4238), 
            .I3(n23526), .O(n7947[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n22573), .I0(GND_net), .I1(n1_adj_4606[15]), 
            .CO(n22574));
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3522_10 (.CI(n23526), .I0(n7959[7]), .I1(n697_adj_4238), 
            .CO(n23527));
    SB_CARRY add_3522_9 (.CI(n23525), .I0(n7959[6]), .I1(n624_adj_4237), 
            .CO(n23526));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4606[14]), .I3(n22572), .O(n29_adj_4196)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3522_8_lut (.I0(GND_net), .I1(n7959[5]), .I2(n551_adj_4235), 
            .I3(n23524), .O(n7947[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_8 (.CI(n23524), .I0(n7959[5]), .I1(n551_adj_4235), 
            .CO(n23525));
    SB_LUT4 add_3522_7_lut (.I0(GND_net), .I1(n7959[4]), .I2(n478_adj_4234), 
            .I3(n23523), .O(n7947[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_7 (.CI(n23523), .I0(n7959[4]), .I1(n478_adj_4234), 
            .CO(n23524));
    SB_LUT4 add_3522_6_lut (.I0(GND_net), .I1(n7959[3]), .I2(n405_adj_4233), 
            .I3(n23522), .O(n7947[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_6 (.CI(n23522), .I0(n7959[3]), .I1(n405_adj_4233), 
            .CO(n23523));
    SB_CARRY unary_minus_5_add_3_16 (.CI(n22572), .I0(GND_net), .I1(n1_adj_4606[14]), 
            .CO(n22573));
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4606[13]), .I3(n22571), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3522_5_lut (.I0(GND_net), .I1(n7959[2]), .I2(n332_adj_4231), 
            .I3(n23521), .O(n7947[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_5 (.CI(n23521), .I0(n7959[2]), .I1(n332_adj_4231), 
            .CO(n23522));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n22571), .I0(GND_net), .I1(n1_adj_4606[13]), 
            .CO(n22572));
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4205));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4606[12]), .I3(n22570), .O(n25_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3522_4_lut (.I0(GND_net), .I1(n7959[1]), .I2(n259_adj_4229), 
            .I3(n23520), .O(n7947[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_4 (.CI(n23520), .I0(n7959[1]), .I1(n259_adj_4229), 
            .CO(n23521));
    SB_LUT4 add_3522_3_lut (.I0(GND_net), .I1(n7959[0]), .I2(n186_adj_4228), 
            .I3(n23519), .O(n7947[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_3 (.CI(n23519), .I0(n7959[0]), .I1(n186_adj_4228), 
            .CO(n23520));
    SB_LUT4 add_3522_2_lut (.I0(GND_net), .I1(n44_adj_4227), .I2(n113_adj_4226), 
            .I3(GND_net), .O(n7947[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n22570), .I0(GND_net), .I1(n1_adj_4606[12]), 
            .CO(n22571));
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4606[11]), .I3(n22569), .O(n23_adj_4195)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_614_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n22569), .I0(GND_net), .I1(n1_adj_4606[11]), 
            .CO(n22570));
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[20]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[21]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4463));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4464));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4465));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4466));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4467));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4468));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4469));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4470));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4471));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4606[10]), .I3(n22568), .O(n21_adj_4188)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4472));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n22568), .I0(GND_net), .I1(n1_adj_4606[10]), 
            .CO(n22569));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4606[9]), .I3(n22567), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n22567), .I0(GND_net), .I1(n1_adj_4606[9]), 
            .CO(n22568));
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4473));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4474));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4475));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4476));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4477));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4478));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4606[8]), .I3(n22566), .O(n17_adj_4189)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n22566), .I0(GND_net), .I1(n1_adj_4606[8]), 
            .CO(n22567));
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4479));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4480));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4606[7]), .I3(n22565), .O(n15_adj_4185)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4481));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4482));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3523_9 (.CI(n23534), .I0(n7970[6]), .I1(n627_adj_4253), 
            .CO(n23535));
    SB_LUT4 add_3523_10_lut (.I0(GND_net), .I1(n7970[7]), .I2(n700_adj_4218), 
            .I3(n23535), .O(n7959[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3523_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4483));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3524_2_lut (.I0(GND_net), .I1(n50_adj_4255), .I2(n119_adj_4254), 
            .I3(GND_net), .O(n7970[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3524_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3522_2 (.CI(GND_net), .I0(n44_adj_4227), .I1(n113_adj_4226), 
            .CO(n23519));
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[22]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3521_12_lut (.I0(GND_net), .I1(n7947[9]), .I2(n840_adj_4217), 
            .I3(n23518), .O(n7934[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4484));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3521_11_lut (.I0(GND_net), .I1(n7947[8]), .I2(n767_adj_4216), 
            .I3(n23517), .O(n7934[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n22565), .I0(GND_net), .I1(n1_adj_4606[7]), 
            .CO(n22566));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4606[6]), .I3(n22564), .O(n13_adj_4186)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4485));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n22564), .I0(GND_net), .I1(n1_adj_4606[6]), 
            .CO(n22565));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4606[5]), .I3(n22563), .O(n11_adj_4187)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3521_11 (.CI(n23517), .I0(n7947[8]), .I1(n767_adj_4216), 
            .CO(n23518));
    SB_LUT4 add_3521_10_lut (.I0(GND_net), .I1(n7947[7]), .I2(n694_adj_4214), 
            .I3(n23516), .O(n7934[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3521_10 (.CI(n23516), .I0(n7947[7]), .I1(n694_adj_4214), 
            .CO(n23517));
    SB_DFFE \PID_CONTROLLER.integral_1209__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[0]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4487));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4488));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n22563), .I0(GND_net), .I1(n1_adj_4606[5]), 
            .CO(n22564));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4606[4]), .I3(n22562), .O(n9_adj_4190)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n22562), .I0(GND_net), .I1(n1_adj_4606[4]), 
            .CO(n22563));
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4489));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4490));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4491));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4492));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4493));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4494));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4495));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4607[23]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4606[3]), .I3(n22561), .O(n7_adj_4193)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n22561), .I0(GND_net), .I1(n1_adj_4606[3]), 
            .CO(n22562));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4606[2]), .I3(n22560), .O(n5_adj_4194)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_614_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n22560), .I0(GND_net), .I1(n1_adj_4606[2]), 
            .CO(n22561));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4606[1]), .I3(n22559), .O(n3_adj_4206)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i18_3_lut (.I0(n155[17]), .I1(PWMLimit[17]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_614_i19_3_lut (.I0(n155[18]), .I1(PWMLimit[18]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4496));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4497));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4498));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4499));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4500));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4501));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4502));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4503));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i20_3_lut (.I0(n155[19]), .I1(PWMLimit[19]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4504));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i21_3_lut (.I0(n155[20]), .I1(PWMLimit[20]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4505));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4506));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4507));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4508));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4509));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4510));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4511));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4512));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_614_i22_3_lut (.I0(n155[21]), .I1(PWMLimit[21]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24782_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30633));   // verilog/motorControl.v(29[14] 48[8])
    defparam i24782_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n22559), .I0(GND_net), .I1(n1_adj_4606[1]), 
            .CO(n22560));
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3655[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3655[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3655[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3655[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3655[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3655[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3655[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3655[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3655[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3655[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3655[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_614_i23_3_lut (.I0(n155[22]), .I1(PWMLimit[22]), .I2(n256_adj_4200), 
            .I3(GND_net), .O(n2933[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_614_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3655[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3655[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3655[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3655[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3655[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3655[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3655[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3655[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3655[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3655[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4515));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3521_9_lut (.I0(GND_net), .I1(n7947[6]), .I2(n621_adj_4219), 
            .I3(n23515), .O(n7934[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3521_9 (.CI(n23515), .I0(n7947[6]), .I1(n621_adj_4219), 
            .CO(n23516));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3532[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4606[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3631 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4606[0]), 
            .CO(n22559));
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4461));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3655[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4518));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3522_9_lut (.I0(GND_net), .I1(n7959[6]), .I2(n624_adj_4237), 
            .I3(n23525), .O(n7947[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3522_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(30[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3521_8 (.CI(n23514), .I0(n7947[5]), .I1(n548_adj_4518), 
            .CO(n23515));
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4606[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4460));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4520));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4521));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4522));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4523));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3532[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i17569_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n22103), .I3(n7718[0]), .O(n4_adj_4458));   // verilog/motorControl.v(34[17:23])
    defparam i17569_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4524));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3521_8_lut (.I0(GND_net), .I1(n7947[5]), .I2(n548_adj_4518), 
            .I3(n23514), .O(n7934[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n7718[0]), .I3(n22103), .O(n7713[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 add_3521_7_lut (.I0(GND_net), .I1(n7947[4]), .I2(n475_adj_4376), 
            .I3(n23513), .O(n7934[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4525));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4526));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17558_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n22103));   // verilog/motorControl.v(34[17:23])
    defparam i17558_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4527));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17556_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n7713[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17556_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4528));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3655[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3679), .I3(GND_net), .O(duty_23__N_3532[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4529));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4530));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4531));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4532));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4533));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4534));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4535));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4536));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4537));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4538));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4539));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4540));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4541));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17538_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n22069), .I3(n7713[0]), .O(n4_adj_4451));   // verilog/motorControl.v(34[17:23])
    defparam i17538_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4542));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3521_6 (.CI(n23512), .I0(n7947[3]), .I1(n402_adj_4205), 
            .CO(n23513));
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4543));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4544));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4545));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4546));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3521_5_lut (.I0(GND_net), .I1(n7947[2]), .I2(n329_adj_4515), 
            .I3(n23511), .O(n7934[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1492 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n7713[0]), .I3(n22069), .O(n7707[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1492.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4547));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17525_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n7707[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17525_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i17527_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n22069));   // verilog/motorControl.v(34[17:23])
    defparam i17527_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4548));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3532[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3532[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3532[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3532[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3532[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3532[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3532[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3532[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3532[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3532[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3532[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3532[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3532[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3532[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3532[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3532[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3532[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3532[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3532[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3532[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3532[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3556 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i17507_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_4549), .I3(n7707[1]), .O(n6_adj_4445));   // verilog/motorControl.v(34[17:23])
    defparam i17507_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1493 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n7707[1]), .I3(n4_adj_4549), .O(n7700[2]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1493.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1494 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n7707[0]), .I3(n22026), .O(n7700[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1494.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17499_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n22026), .I3(n7707[0]), .O(n4_adj_4549));   // verilog/motorControl.v(34[17:23])
    defparam i17499_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17486_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n7700[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17486_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i17488_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n22026));   // verilog/motorControl.v(34[17:23])
    defparam i17488_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_3521_5 (.CI(n23511), .I0(n7947[2]), .I1(n329_adj_4515), 
            .CO(n23512));
    SB_LUT4 add_3521_4_lut (.I0(GND_net), .I1(n7947[1]), .I2(n256_adj_4512), 
            .I3(n23510), .O(n7934[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3521_4 (.CI(n23510), .I0(n7947[1]), .I1(n256_adj_4512), 
            .CO(n23511));
    SB_LUT4 add_3521_3_lut (.I0(GND_net), .I1(n7947[0]), .I2(n183_adj_4511), 
            .I3(n23509), .O(n7934[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3521_3 (.CI(n23509), .I0(n7947[0]), .I1(n183_adj_4511), 
            .CO(n23510));
    SB_LUT4 add_3521_2_lut (.I0(GND_net), .I1(n41_adj_4510), .I2(n110_adj_4509), 
            .I3(GND_net), .O(n7934[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3521_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3521_2 (.CI(GND_net), .I0(n41_adj_4510), .I1(n110_adj_4509), 
            .CO(n23509));
    SB_LUT4 add_3520_13_lut (.I0(GND_net), .I1(n7934[10]), .I2(n910_adj_4508), 
            .I3(n23508), .O(n7920[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3520_12_lut (.I0(GND_net), .I1(n7934[9]), .I2(n837_adj_4507), 
            .I3(n23507), .O(n7920[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_12 (.CI(n23507), .I0(n7934[9]), .I1(n837_adj_4507), 
            .CO(n23508));
    SB_LUT4 add_3520_11_lut (.I0(GND_net), .I1(n7934[8]), .I2(n764_adj_4506), 
            .I3(n23506), .O(n7920[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_11 (.CI(n23506), .I0(n7934[8]), .I1(n764_adj_4506), 
            .CO(n23507));
    SB_LUT4 add_3520_10_lut (.I0(GND_net), .I1(n7934[7]), .I2(n691_adj_4505), 
            .I3(n23505), .O(n7920[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_10 (.CI(n23505), .I0(n7934[7]), .I1(n691_adj_4505), 
            .CO(n23506));
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4419));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24123_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n29975));   // verilog/motorControl.v(36[10:25])
    defparam i24123_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_4444));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_3520_9_lut (.I0(GND_net), .I1(n7934[6]), .I2(n618_adj_4504), 
            .I3(n23504), .O(n7920[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_9 (.CI(n23504), .I0(n7934[6]), .I1(n618_adj_4504), 
            .CO(n23505));
    SB_LUT4 add_3520_8_lut (.I0(GND_net), .I1(n7934[5]), .I2(n545_adj_4503), 
            .I3(n23503), .O(n7920[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_8 (.CI(n23503), .I0(n7934[5]), .I1(n545_adj_4503), 
            .CO(n23504));
    SB_LUT4 add_3520_7_lut (.I0(GND_net), .I1(n7934[4]), .I2(n472_adj_4502), 
            .I3(n23502), .O(n7920[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_7 (.CI(n23502), .I0(n7934[4]), .I1(n472_adj_4502), 
            .CO(n23503));
    SB_LUT4 add_3520_6_lut (.I0(GND_net), .I1(n7934[3]), .I2(n399_adj_4501), 
            .I3(n23501), .O(n7920[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_6 (.CI(n23501), .I0(n7934[3]), .I1(n399_adj_4501), 
            .CO(n23502));
    SB_LUT4 add_3520_5_lut (.I0(GND_net), .I1(n7934[2]), .I2(n326_adj_4500), 
            .I3(n23500), .O(n7920[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_5 (.CI(n23500), .I0(n7934[2]), .I1(n326_adj_4500), 
            .CO(n23501));
    SB_LUT4 add_3520_4_lut (.I0(GND_net), .I1(n7934[1]), .I2(n253_adj_4499), 
            .I3(n23499), .O(n7920[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_4 (.CI(n23499), .I0(n7934[1]), .I1(n253_adj_4499), 
            .CO(n23500));
    SB_LUT4 add_3520_3_lut (.I0(GND_net), .I1(n7934[0]), .I2(n180_adj_4498), 
            .I3(n23498), .O(n7920[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3520_3 (.CI(n23498), .I0(n7934[0]), .I1(n180_adj_4498), 
            .CO(n23499));
    SB_LUT4 add_3520_2_lut (.I0(GND_net), .I1(n38_adj_4497), .I2(n107_adj_4496), 
            .I3(GND_net), .O(n7920[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3520_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4411));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3520_2 (.CI(GND_net), .I0(n38_adj_4497), .I1(n107_adj_4496), 
            .CO(n23498));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n22846), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n22845), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_24  (.CI(n22845), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n22846));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n22844), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_23  (.CI(n22844), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n22845));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n22843), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_22  (.CI(n22843), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n22844));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n22842), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_21  (.CI(n22842), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n22843));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n22841), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_20  (.CI(n22841), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n22842));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n22840), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_19  (.CI(n22840), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n22841));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n22839), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_18  (.CI(n22839), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n22840));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n22838), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_17  (.CI(n22838), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n22839));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n22837), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_16  (.CI(n22837), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n22838));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n22836), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_15  (.CI(n22836), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n22837));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n22835), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_14  (.CI(n22835), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n22836));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n22834), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_13  (.CI(n22834), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n22835));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n22833), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_12  (.CI(n22833), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n22834));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n22832), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_11  (.CI(n22832), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n22833));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n22831), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_10  (.CI(n22831), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n22832));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n22830), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_9  (.CI(n22830), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n22831));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n22829), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_8  (.CI(n22829), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n22830));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n22828), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_7  (.CI(n22828), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n22829));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n22827), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_6  (.CI(n22827), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n22828));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n22826), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_5  (.CI(n22826), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n22827));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n22825), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3519_14_lut (.I0(GND_net), .I1(n7920[11]), .I2(n980_adj_4495), 
            .I3(n23497), .O(n7905[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_4  (.CI(n22825), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n22826));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n22824), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3519_13_lut (.I0(GND_net), .I1(n7920[10]), .I2(n907_adj_4494), 
            .I3(n23496), .O(n7905[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_3  (.CI(n22824), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n22825));
    SB_LUT4 \PID_CONTROLLER.integral_1209_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1209_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1209_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n22824));
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4412));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4409));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4408));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3519_13 (.CI(n23496), .I0(n7920[10]), .I1(n907_adj_4494), 
            .CO(n23497));
    SB_LUT4 add_3519_12_lut (.I0(GND_net), .I1(n7920[9]), .I2(n834_adj_4493), 
            .I3(n23495), .O(n7905[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_12 (.CI(n23495), .I0(n7920[9]), .I1(n834_adj_4493), 
            .CO(n23496));
    SB_LUT4 add_3519_11_lut (.I0(GND_net), .I1(n7920[8]), .I2(n761_adj_4492), 
            .I3(n23494), .O(n7905[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_11 (.CI(n23494), .I0(n7920[8]), .I1(n761_adj_4492), 
            .CO(n23495));
    SB_LUT4 add_3519_10_lut (.I0(GND_net), .I1(n7920[7]), .I2(n688_adj_4491), 
            .I3(n23493), .O(n7905[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_10 (.CI(n23493), .I0(n7920[7]), .I1(n688_adj_4491), 
            .CO(n23494));
    SB_LUT4 add_3519_9_lut (.I0(GND_net), .I1(n7920[6]), .I2(n615_adj_4490), 
            .I3(n23492), .O(n7905[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_9 (.CI(n23492), .I0(n7920[6]), .I1(n615_adj_4490), 
            .CO(n23493));
    SB_LUT4 add_3519_8_lut (.I0(GND_net), .I1(n7920[5]), .I2(n542_adj_4489), 
            .I3(n23491), .O(n7905[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_8 (.CI(n23491), .I0(n7920[5]), .I1(n542_adj_4489), 
            .CO(n23492));
    SB_LUT4 add_3519_7_lut (.I0(GND_net), .I1(n7920[4]), .I2(n469_adj_4488), 
            .I3(n23490), .O(n7905[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_7 (.CI(n23490), .I0(n7920[4]), .I1(n469_adj_4488), 
            .CO(n23491));
    SB_LUT4 add_3519_6_lut (.I0(GND_net), .I1(n7920[3]), .I2(n396_adj_4487), 
            .I3(n23489), .O(n7905[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_6 (.CI(n23489), .I0(n7920[3]), .I1(n396_adj_4487), 
            .CO(n23490));
    SB_LUT4 add_3519_5_lut (.I0(GND_net), .I1(n7920[2]), .I2(n323_adj_4485), 
            .I3(n23488), .O(n7905[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_5 (.CI(n23488), .I0(n7920[2]), .I1(n323_adj_4485), 
            .CO(n23489));
    SB_LUT4 add_3519_4_lut (.I0(GND_net), .I1(n7920[1]), .I2(n250_adj_4484), 
            .I3(n23487), .O(n7905[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_4 (.CI(n23487), .I0(n7920[1]), .I1(n250_adj_4484), 
            .CO(n23488));
    SB_LUT4 add_3519_3_lut (.I0(GND_net), .I1(n7920[0]), .I2(n177_adj_4483), 
            .I3(n23486), .O(n7905[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_3 (.CI(n23486), .I0(n7920[0]), .I1(n177_adj_4483), 
            .CO(n23487));
    SB_LUT4 add_3519_2_lut (.I0(GND_net), .I1(n35_adj_4482), .I2(n104_adj_4481), 
            .I3(GND_net), .O(n7905[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3519_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3519_2 (.CI(GND_net), .I0(n35_adj_4482), .I1(n104_adj_4481), 
            .CO(n23486));
    SB_LUT4 add_3518_15_lut (.I0(GND_net), .I1(n7905[12]), .I2(n1050_adj_4480), 
            .I3(n23485), .O(n7889[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3518_14_lut (.I0(GND_net), .I1(n7905[11]), .I2(n977_adj_4479), 
            .I3(n23484), .O(n7889[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_14 (.CI(n23484), .I0(n7905[11]), .I1(n977_adj_4479), 
            .CO(n23485));
    SB_LUT4 add_3518_13_lut (.I0(GND_net), .I1(n7905[10]), .I2(n904_adj_4478), 
            .I3(n23483), .O(n7889[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_13 (.CI(n23483), .I0(n7905[10]), .I1(n904_adj_4478), 
            .CO(n23484));
    SB_LUT4 add_3518_12_lut (.I0(GND_net), .I1(n7905[9]), .I2(n831_adj_4477), 
            .I3(n23482), .O(n7889[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_12 (.CI(n23482), .I0(n7905[9]), .I1(n831_adj_4477), 
            .CO(n23483));
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4557));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3518_11_lut (.I0(GND_net), .I1(n7905[8]), .I2(n758_adj_4476), 
            .I3(n23481), .O(n7889[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_11 (.CI(n23481), .I0(n7905[8]), .I1(n758_adj_4476), 
            .CO(n23482));
    SB_LUT4 add_3518_10_lut (.I0(GND_net), .I1(n7905[7]), .I2(n685_adj_4475), 
            .I3(n23480), .O(n7889[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_10 (.CI(n23480), .I0(n7905[7]), .I1(n685_adj_4475), 
            .CO(n23481));
    SB_LUT4 add_3518_9_lut (.I0(GND_net), .I1(n7905[6]), .I2(n612_adj_4474), 
            .I3(n23479), .O(n7889[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_9 (.CI(n23479), .I0(n7905[6]), .I1(n612_adj_4474), 
            .CO(n23480));
    SB_LUT4 add_3518_8_lut (.I0(GND_net), .I1(n7905[5]), .I2(n539_adj_4473), 
            .I3(n23478), .O(n7889[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_8 (.CI(n23478), .I0(n7905[5]), .I1(n539_adj_4473), 
            .CO(n23479));
    SB_LUT4 add_3518_7_lut (.I0(GND_net), .I1(n7905[4]), .I2(n466_adj_4472), 
            .I3(n23477), .O(n7889[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_7 (.CI(n23477), .I0(n7905[4]), .I1(n466_adj_4472), 
            .CO(n23478));
    SB_LUT4 add_3518_6_lut (.I0(GND_net), .I1(n7905[3]), .I2(n393_adj_4471), 
            .I3(n23476), .O(n7889[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_6 (.CI(n23476), .I0(n7905[3]), .I1(n393_adj_4471), 
            .CO(n23477));
    SB_LUT4 add_3518_5_lut (.I0(GND_net), .I1(n7905[2]), .I2(n320_adj_4470), 
            .I3(n23475), .O(n7889[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_5 (.CI(n23475), .I0(n7905[2]), .I1(n320_adj_4470), 
            .CO(n23476));
    SB_LUT4 add_3518_4_lut (.I0(GND_net), .I1(n7905[1]), .I2(n247_adj_4469), 
            .I3(n23474), .O(n7889[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_4 (.CI(n23474), .I0(n7905[1]), .I1(n247_adj_4469), 
            .CO(n23475));
    SB_LUT4 add_3518_3_lut (.I0(GND_net), .I1(n7905[0]), .I2(n174_adj_4468), 
            .I3(n23473), .O(n7889[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_3 (.CI(n23473), .I0(n7905[0]), .I1(n174_adj_4468), 
            .CO(n23474));
    SB_LUT4 add_3518_2_lut (.I0(GND_net), .I1(n32_adj_4467), .I2(n101_adj_4466), 
            .I3(GND_net), .O(n7889[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3518_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3518_2 (.CI(GND_net), .I0(n32_adj_4467), .I1(n101_adj_4466), 
            .CO(n23473));
    SB_LUT4 add_3517_16_lut (.I0(GND_net), .I1(n7889[13]), .I2(n1120_adj_4465), 
            .I3(n23472), .O(n7872[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3517_15_lut (.I0(GND_net), .I1(n7889[12]), .I2(n1047_adj_4464), 
            .I3(n23471), .O(n7872[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_15 (.CI(n23471), .I0(n7889[12]), .I1(n1047_adj_4464), 
            .CO(n23472));
    SB_LUT4 add_3517_14_lut (.I0(GND_net), .I1(n7889[11]), .I2(n974_adj_4463), 
            .I3(n23470), .O(n7872[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_14 (.CI(n23470), .I0(n7889[11]), .I1(n974_adj_4463), 
            .CO(n23471));
    SB_LUT4 i17629_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_4558), .I3(n8004[1]), .O(n6_adj_4335));   // verilog/motorControl.v(34[26:37])
    defparam i17629_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1495 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8004[1]), .I3(n4_adj_4558), .O(n7997[2]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1495.LUT_INIT = 16'h8778;
    SB_LUT4 add_3517_13_lut (.I0(GND_net), .I1(n7889[10]), .I2(n901_adj_4559), 
            .I3(n23469), .O(n7872[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_13 (.CI(n23469), .I0(n7889[10]), .I1(n901_adj_4559), 
            .CO(n23470));
    SB_LUT4 add_3517_12_lut (.I0(GND_net), .I1(n7889[9]), .I2(n828_adj_4560), 
            .I3(n23468), .O(n7872[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_12 (.CI(n23468), .I0(n7889[9]), .I1(n828_adj_4560), 
            .CO(n23469));
    SB_LUT4 add_3517_11_lut (.I0(GND_net), .I1(n7889[8]), .I2(n755_adj_4561), 
            .I3(n23467), .O(n7872[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_11 (.CI(n23467), .I0(n7889[8]), .I1(n755_adj_4561), 
            .CO(n23468));
    SB_LUT4 add_3517_10_lut (.I0(GND_net), .I1(n7889[7]), .I2(n682_adj_4562), 
            .I3(n23466), .O(n7872[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_10 (.CI(n23466), .I0(n7889[7]), .I1(n682_adj_4562), 
            .CO(n23467));
    SB_LUT4 add_3517_9_lut (.I0(GND_net), .I1(n7889[6]), .I2(n609_adj_4563), 
            .I3(n23465), .O(n7872[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_9 (.CI(n23465), .I0(n7889[6]), .I1(n609_adj_4563), 
            .CO(n23466));
    SB_LUT4 add_3517_8_lut (.I0(GND_net), .I1(n7889[5]), .I2(n536_adj_4564), 
            .I3(n23464), .O(n7872[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_8 (.CI(n23464), .I0(n7889[5]), .I1(n536_adj_4564), 
            .CO(n23465));
    SB_LUT4 add_3517_7_lut (.I0(GND_net), .I1(n7889[4]), .I2(n463_adj_4565), 
            .I3(n23463), .O(n7872[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_7 (.CI(n23463), .I0(n7889[4]), .I1(n463_adj_4565), 
            .CO(n23464));
    SB_LUT4 add_3517_6_lut (.I0(GND_net), .I1(n7889[3]), .I2(n390_adj_4566), 
            .I3(n23462), .O(n7872[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_6 (.CI(n23462), .I0(n7889[3]), .I1(n390_adj_4566), 
            .CO(n23463));
    SB_LUT4 add_3517_5_lut (.I0(GND_net), .I1(n7889[2]), .I2(n317_adj_4567), 
            .I3(n23461), .O(n7872[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_5 (.CI(n23461), .I0(n7889[2]), .I1(n317_adj_4567), 
            .CO(n23462));
    SB_LUT4 add_3517_4_lut (.I0(GND_net), .I1(n7889[1]), .I2(n244_adj_4568), 
            .I3(n23460), .O(n7872[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_4 (.CI(n23460), .I0(n7889[1]), .I1(n244_adj_4568), 
            .CO(n23461));
    SB_LUT4 add_3517_3_lut (.I0(GND_net), .I1(n7889[0]), .I2(n171_adj_4569), 
            .I3(n23459), .O(n7872[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_3 (.CI(n23459), .I0(n7889[0]), .I1(n171_adj_4569), 
            .CO(n23460));
    SB_LUT4 add_3517_2_lut (.I0(GND_net), .I1(n29_adj_4570), .I2(n98_adj_4571), 
            .I3(GND_net), .O(n7872[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_2 (.CI(GND_net), .I0(n29_adj_4570), .I1(n98_adj_4571), 
            .CO(n23459));
    SB_LUT4 add_3516_17_lut (.I0(GND_net), .I1(n7872[14]), .I2(GND_net), 
            .I3(n23458), .O(n7854[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_16_lut (.I0(GND_net), .I1(n7872[13]), .I2(n1117_adj_4572), 
            .I3(n23457), .O(n7854[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_16 (.CI(n23457), .I0(n7872[13]), .I1(n1117_adj_4572), 
            .CO(n23458));
    SB_LUT4 add_3516_15_lut (.I0(GND_net), .I1(n7872[12]), .I2(n1044_adj_4573), 
            .I3(n23456), .O(n7854[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_15 (.CI(n23456), .I0(n7872[12]), .I1(n1044_adj_4573), 
            .CO(n23457));
    SB_LUT4 add_3516_14_lut (.I0(GND_net), .I1(n7872[11]), .I2(n971_adj_4574), 
            .I3(n23455), .O(n7854[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_14 (.CI(n23455), .I0(n7872[11]), .I1(n971_adj_4574), 
            .CO(n23456));
    SB_LUT4 add_3516_13_lut (.I0(GND_net), .I1(n7872[10]), .I2(n898_adj_4575), 
            .I3(n23454), .O(n7854[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_13 (.CI(n23454), .I0(n7872[10]), .I1(n898_adj_4575), 
            .CO(n23455));
    SB_LUT4 add_3516_12_lut (.I0(GND_net), .I1(n7872[9]), .I2(n825_adj_4576), 
            .I3(n23453), .O(n7854[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_12 (.CI(n23453), .I0(n7872[9]), .I1(n825_adj_4576), 
            .CO(n23454));
    SB_LUT4 add_3516_11_lut (.I0(GND_net), .I1(n7872[8]), .I2(n752_adj_4577), 
            .I3(n23452), .O(n7854[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_11 (.CI(n23452), .I0(n7872[8]), .I1(n752_adj_4577), 
            .CO(n23453));
    SB_LUT4 add_3516_10_lut (.I0(GND_net), .I1(n7872[7]), .I2(n679_adj_4578), 
            .I3(n23451), .O(n7854[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_10 (.CI(n23451), .I0(n7872[7]), .I1(n679_adj_4578), 
            .CO(n23452));
    SB_LUT4 add_3516_9_lut (.I0(GND_net), .I1(n7872[6]), .I2(n606_adj_4579), 
            .I3(n23450), .O(n7854[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_9 (.CI(n23450), .I0(n7872[6]), .I1(n606_adj_4579), 
            .CO(n23451));
    SB_LUT4 add_3516_8_lut (.I0(GND_net), .I1(n7872[5]), .I2(n533_adj_4580), 
            .I3(n23449), .O(n7854[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_4448));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3516_8 (.CI(n23449), .I0(n7872[5]), .I1(n533_adj_4580), 
            .CO(n23450));
    SB_LUT4 add_3516_7_lut (.I0(GND_net), .I1(n7872[4]), .I2(n460_adj_4581), 
            .I3(n23448), .O(n7854[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_7 (.CI(n23448), .I0(n7872[4]), .I1(n460_adj_4581), 
            .CO(n23449));
    SB_LUT4 add_3516_6_lut (.I0(GND_net), .I1(n7872[3]), .I2(n387_adj_4582), 
            .I3(n23447), .O(n7854[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_6 (.CI(n23447), .I0(n7872[3]), .I1(n387_adj_4582), 
            .CO(n23448));
    SB_LUT4 add_3516_5_lut (.I0(GND_net), .I1(n7872[2]), .I2(n314_adj_4583), 
            .I3(n23446), .O(n7854[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_5 (.CI(n23446), .I0(n7872[2]), .I1(n314_adj_4583), 
            .CO(n23447));
    SB_LUT4 i2_3_lut_4_lut_adj_1496 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8004[0]), .I3(n22158), .O(n7997[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1496.LUT_INIT = 16'h8778;
    SB_LUT4 i17621_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n22158), .I3(n8004[0]), .O(n4_adj_4558));   // verilog/motorControl.v(34[26:37])
    defparam i17621_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_3516_4_lut (.I0(GND_net), .I1(n7872[1]), .I2(n241_adj_4584), 
            .I3(n23445), .O(n7854[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_4 (.CI(n23445), .I0(n7872[1]), .I1(n241_adj_4584), 
            .CO(n23446));
    SB_LUT4 i17610_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n22158));   // verilog/motorControl.v(34[26:37])
    defparam i17610_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3516_3_lut (.I0(GND_net), .I1(n7872[0]), .I2(n168_adj_4585), 
            .I3(n23444), .O(n7854[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17608_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n7997[0]));   // verilog/motorControl.v(34[26:37])
    defparam i17608_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_3516_3 (.CI(n23444), .I0(n7872[0]), .I1(n168_adj_4585), 
            .CO(n23445));
    SB_LUT4 add_3516_2_lut (.I0(GND_net), .I1(n26_adj_4586), .I2(n95_adj_4587), 
            .I3(GND_net), .O(n7854[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_2 (.CI(GND_net), .I0(n26_adj_4586), .I1(n95_adj_4587), 
            .CO(n23444));
    SB_LUT4 i24088_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n29940));
    defparam i24088_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_3515_18_lut (.I0(GND_net), .I1(n7854[15]), .I2(GND_net), 
            .I3(n23443), .O(n7835[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3515_17_lut (.I0(GND_net), .I1(n7854[14]), .I2(GND_net), 
            .I3(n23442), .O(n7835[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_4446));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3515_17 (.CI(n23442), .I0(n7854[14]), .I1(GND_net), .CO(n23443));
    SB_LUT4 add_3515_16_lut (.I0(GND_net), .I1(n7854[13]), .I2(n1114_adj_4588), 
            .I3(n23441), .O(n7835[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_16 (.CI(n23441), .I0(n7854[13]), .I1(n1114_adj_4588), 
            .CO(n23442));
    SB_LUT4 add_3515_15_lut (.I0(GND_net), .I1(n7854[12]), .I2(n1041_adj_4589), 
            .I3(n23440), .O(n7835[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_15 (.CI(n23440), .I0(n7854[12]), .I1(n1041_adj_4589), 
            .CO(n23441));
    SB_LUT4 add_3515_14_lut (.I0(GND_net), .I1(n7854[11]), .I2(n968_adj_4590), 
            .I3(n23439), .O(n7835[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_4450));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3515_14 (.CI(n23439), .I0(n7854[11]), .I1(n968_adj_4590), 
            .CO(n23440));
    SB_LUT4 add_3515_13_lut (.I0(GND_net), .I1(n7854[10]), .I2(n895_adj_4591), 
            .I3(n23438), .O(n7835[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_13 (.CI(n23438), .I0(n7854[10]), .I1(n895_adj_4591), 
            .CO(n23439));
    SB_LUT4 add_3515_12_lut (.I0(GND_net), .I1(n7854[9]), .I2(n822_adj_4592), 
            .I3(n23437), .O(n7835[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_12 (.CI(n23437), .I0(n7854[9]), .I1(n822_adj_4592), 
            .CO(n23438));
    SB_LUT4 add_3515_11_lut (.I0(GND_net), .I1(n7854[8]), .I2(n749_adj_4593), 
            .I3(n23436), .O(n7835[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_11 (.CI(n23436), .I0(n7854[8]), .I1(n749_adj_4593), 
            .CO(n23437));
    SB_LUT4 add_3515_10_lut (.I0(GND_net), .I1(n7854[7]), .I2(n676_adj_4594), 
            .I3(n23435), .O(n7835[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_10 (.CI(n23435), .I0(n7854[7]), .I1(n676_adj_4594), 
            .CO(n23436));
    SB_LUT4 add_3515_9_lut (.I0(GND_net), .I1(n7854[6]), .I2(n603_adj_4595), 
            .I3(n23434), .O(n7835[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_9 (.CI(n23434), .I0(n7854[6]), .I1(n603_adj_4595), 
            .CO(n23435));
    SB_LUT4 add_3515_8_lut (.I0(GND_net), .I1(n7854[5]), .I2(n530_adj_4596), 
            .I3(n23433), .O(n7835[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_8 (.CI(n23433), .I0(n7854[5]), .I1(n530_adj_4596), 
            .CO(n23434));
    SB_LUT4 add_3515_7_lut (.I0(GND_net), .I1(n7854[4]), .I2(n457_adj_4597), 
            .I3(n23432), .O(n7835[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4598));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3515_7 (.CI(n23432), .I0(n7854[4]), .I1(n457_adj_4597), 
            .CO(n23433));
    SB_LUT4 add_3515_6_lut (.I0(GND_net), .I1(n7854[3]), .I2(n384_adj_4599), 
            .I3(n23431), .O(n7835[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_6 (.CI(n23431), .I0(n7854[3]), .I1(n384_adj_4599), 
            .CO(n23432));
    SB_LUT4 add_3515_5_lut (.I0(GND_net), .I1(n7854[2]), .I2(n311_adj_4600), 
            .I3(n23430), .O(n7835[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24098_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n29950));
    defparam i24098_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_3515_5 (.CI(n23430), .I0(n7854[2]), .I1(n311_adj_4600), 
            .CO(n23431));
    SB_LUT4 add_3515_4_lut (.I0(GND_net), .I1(n7854[1]), .I2(n238_adj_4601), 
            .I3(n23429), .O(n7835[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_4 (.CI(n23429), .I0(n7854[1]), .I1(n238_adj_4601), 
            .CO(n23430));
    SB_LUT4 add_3515_3_lut (.I0(GND_net), .I1(n7854[0]), .I2(n165_adj_4602), 
            .I3(n23428), .O(n7835[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_3 (.CI(n23428), .I0(n7854[0]), .I1(n165_adj_4602), 
            .CO(n23429));
    SB_LUT4 add_3515_2_lut (.I0(GND_net), .I1(n23_adj_4603), .I2(n92_adj_4604), 
            .I3(GND_net), .O(n7835[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3515_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3515_2 (.CI(GND_net), .I0(n23_adj_4603), .I1(n92_adj_4604), 
            .CO(n23428));
    SB_LUT4 add_3514_19_lut (.I0(GND_net), .I1(n7835[16]), .I2(GND_net), 
            .I3(n23427), .O(n7815[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3514_18_lut (.I0(GND_net), .I1(n7835[15]), .I2(GND_net), 
            .I3(n23426), .O(n7815[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_18 (.CI(n23426), .I0(n7835[15]), .I1(GND_net), .CO(n23427));
    SB_LUT4 add_3514_17_lut (.I0(GND_net), .I1(n7835[14]), .I2(GND_net), 
            .I3(n23425), .O(n7815[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_17 (.CI(n23425), .I0(n7835[14]), .I1(GND_net), .CO(n23426));
    SB_LUT4 add_3514_16_lut (.I0(GND_net), .I1(n7835[13]), .I2(n1111_adj_4605), 
            .I3(n23424), .O(n7815[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_16 (.CI(n23424), .I0(n7835[13]), .I1(n1111_adj_4605), 
            .CO(n23425));
    SB_LUT4 add_3514_15_lut (.I0(GND_net), .I1(n7835[12]), .I2(n1038_adj_4598), 
            .I3(n23423), .O(n7815[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_15 (.CI(n23423), .I0(n7835[12]), .I1(n1038_adj_4598), 
            .CO(n23424));
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_4441));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4605));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24054_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n29906));
    defparam i24054_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i24064_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n29916));
    defparam i24064_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i17691_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n22235), .I3(n8015[0]), .O(n4_adj_4369));   // verilog/motorControl.v(34[26:37])
    defparam i17691_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4604));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4603));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4602));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17647_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral [19]), .O(n8004[0]));   // verilog/motorControl.v(34[26:37])
    defparam i17647_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i2_3_lut_4_lut_adj_1497 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n8015[0]), .I3(n22235), .O(n8010[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1497.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4601));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1498 (.I0(n62), .I1(n131), .I2(n8010[0]), 
            .I3(n204), .O(n8004[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1498.LUT_INIT = 16'h8778;
    SB_LUT4 add_3514_14_lut (.I0(GND_net), .I1(n7835[11]), .I2(n965_adj_4557), 
            .I3(n23422), .O(n7815[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4600));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4599));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17660_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n8010[0]), 
            .O(n4_adj_4361));   // verilog/motorControl.v(34[26:37])
    defparam i17660_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i17680_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n22235));   // verilog/motorControl.v(34[26:37])
    defparam i17680_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i17678_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n8010[0]));   // verilog/motorControl.v(34[26:37])
    defparam i17678_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4410));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24086_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n29938));   // verilog/motorControl.v(38[19:35])
    defparam i24086_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4597));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_4415));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4596));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4595));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4594));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4593));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4592));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4591));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4590));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4589));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4588));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4587));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4586));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4585));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4584));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4583));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4582));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE \PID_CONTROLLER.integral_1209__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[1]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[2]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[3]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[4]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[5]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[6]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[7]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[8]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[9]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[10]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[11]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[12]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[13]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[14]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[15]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[16]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[17]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[18]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[19]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[20]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[21]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[22]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1209__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3628 ), .D(n28[23]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4581));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3514_14 (.CI(n23422), .I0(n7835[11]), .I1(n965_adj_4557), 
            .CO(n23423));
    SB_LUT4 add_3514_13_lut (.I0(GND_net), .I1(n7835[10]), .I2(n892_adj_4548), 
            .I3(n23421), .O(n7815[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_13 (.CI(n23421), .I0(n7835[10]), .I1(n892_adj_4548), 
            .CO(n23422));
    SB_LUT4 add_3514_12_lut (.I0(GND_net), .I1(n7835[9]), .I2(n819_adj_4547), 
            .I3(n23420), .O(n7815[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4580));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3514_12 (.CI(n23420), .I0(n7835[9]), .I1(n819_adj_4547), 
            .CO(n23421));
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4579));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3514_11_lut (.I0(GND_net), .I1(n7835[8]), .I2(n746_adj_4546), 
            .I3(n23419), .O(n7815[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_11 (.CI(n23419), .I0(n7835[8]), .I1(n746_adj_4546), 
            .CO(n23420));
    SB_LUT4 add_3514_10_lut (.I0(GND_net), .I1(n7835[7]), .I2(n673_adj_4545), 
            .I3(n23418), .O(n7815[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_10 (.CI(n23418), .I0(n7835[7]), .I1(n673_adj_4545), 
            .CO(n23419));
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4578));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3514_9_lut (.I0(GND_net), .I1(n7835[6]), .I2(n600_adj_4544), 
            .I3(n23417), .O(n7815[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_9 (.CI(n23417), .I0(n7835[6]), .I1(n600_adj_4544), 
            .CO(n23418));
    SB_LUT4 add_3514_8_lut (.I0(GND_net), .I1(n7835[5]), .I2(n527_adj_4543), 
            .I3(n23416), .O(n7815[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4577));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3514_8 (.CI(n23416), .I0(n7835[5]), .I1(n527_adj_4543), 
            .CO(n23417));
    SB_LUT4 add_3514_7_lut (.I0(GND_net), .I1(n7835[4]), .I2(n454_adj_4542), 
            .I3(n23415), .O(n7815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_7 (.CI(n23415), .I0(n7835[4]), .I1(n454_adj_4542), 
            .CO(n23416));
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4576));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3514_6_lut (.I0(GND_net), .I1(n7835[3]), .I2(n381_adj_4541), 
            .I3(n23414), .O(n7815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_6 (.CI(n23414), .I0(n7835[3]), .I1(n381_adj_4541), 
            .CO(n23415));
    SB_LUT4 add_3514_5_lut (.I0(GND_net), .I1(n7835[2]), .I2(n308_adj_4540), 
            .I3(n23413), .O(n7815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_5 (.CI(n23413), .I0(n7835[2]), .I1(n308_adj_4540), 
            .CO(n23414));
    SB_LUT4 add_3514_4_lut (.I0(GND_net), .I1(n7835[1]), .I2(n235_adj_4539), 
            .I3(n23412), .O(n7815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_4 (.CI(n23412), .I0(n7835[1]), .I1(n235_adj_4539), 
            .CO(n23413));
    SB_LUT4 add_3514_3_lut (.I0(GND_net), .I1(n7835[0]), .I2(n162_adj_4538), 
            .I3(n23411), .O(n7815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_3 (.CI(n23411), .I0(n7835[0]), .I1(n162_adj_4538), 
            .CO(n23412));
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4575));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3514_2_lut (.I0(GND_net), .I1(n20_adj_4537), .I2(n89_adj_4536), 
            .I3(GND_net), .O(n7815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3514_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3514_2 (.CI(GND_net), .I0(n20_adj_4537), .I1(n89_adj_4536), 
            .CO(n23411));
    SB_LUT4 add_3513_20_lut (.I0(GND_net), .I1(n7815[17]), .I2(GND_net), 
            .I3(n23410), .O(n7794[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4574));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3513_19_lut (.I0(GND_net), .I1(n7815[16]), .I2(GND_net), 
            .I3(n23409), .O(n7794[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_19 (.CI(n23409), .I0(n7815[16]), .I1(GND_net), .CO(n23410));
    SB_LUT4 add_3513_18_lut (.I0(GND_net), .I1(n7815[15]), .I2(GND_net), 
            .I3(n23408), .O(n7794[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_18 (.CI(n23408), .I0(n7815[15]), .I1(GND_net), .CO(n23409));
    SB_LUT4 add_3513_17_lut (.I0(GND_net), .I1(n7815[14]), .I2(GND_net), 
            .I3(n23407), .O(n7794[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_17 (.CI(n23407), .I0(n7815[14]), .I1(GND_net), .CO(n23408));
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4573));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3513_16_lut (.I0(GND_net), .I1(n7815[13]), .I2(n1108_adj_4535), 
            .I3(n23406), .O(n7794[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_16 (.CI(n23406), .I0(n7815[13]), .I1(n1108_adj_4535), 
            .CO(n23407));
    SB_LUT4 add_3513_15_lut (.I0(GND_net), .I1(n7815[12]), .I2(n1035_adj_4534), 
            .I3(n23405), .O(n7794[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_15 (.CI(n23405), .I0(n7815[12]), .I1(n1035_adj_4534), 
            .CO(n23406));
    SB_LUT4 add_3513_14_lut (.I0(GND_net), .I1(n7815[11]), .I2(n962_adj_4533), 
            .I3(n23404), .O(n7794[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4572));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3513_14 (.CI(n23404), .I0(n7815[11]), .I1(n962_adj_4533), 
            .CO(n23405));
    SB_LUT4 add_3513_13_lut (.I0(GND_net), .I1(n7815[10]), .I2(n889_adj_4532), 
            .I3(n23403), .O(n7794[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_13 (.CI(n23403), .I0(n7815[10]), .I1(n889_adj_4532), 
            .CO(n23404));
    SB_LUT4 add_3513_12_lut (.I0(GND_net), .I1(n7815[9]), .I2(n816_adj_4531), 
            .I3(n23402), .O(n7794[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_12 (.CI(n23402), .I0(n7815[9]), .I1(n816_adj_4531), 
            .CO(n23403));
    SB_LUT4 add_3513_11_lut (.I0(GND_net), .I1(n7815[8]), .I2(n743_adj_4530), 
            .I3(n23401), .O(n7794[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_11 (.CI(n23401), .I0(n7815[8]), .I1(n743_adj_4530), 
            .CO(n23402));
    SB_LUT4 add_3513_10_lut (.I0(GND_net), .I1(n7815[7]), .I2(n670_adj_4529), 
            .I3(n23400), .O(n7794[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_10 (.CI(n23400), .I0(n7815[7]), .I1(n670_adj_4529), 
            .CO(n23401));
    SB_LUT4 add_3513_9_lut (.I0(GND_net), .I1(n7815[6]), .I2(n597_adj_4528), 
            .I3(n23399), .O(n7794[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_9 (.CI(n23399), .I0(n7815[6]), .I1(n597_adj_4528), 
            .CO(n23400));
    SB_LUT4 add_3513_8_lut (.I0(GND_net), .I1(n7815[5]), .I2(n524_adj_4527), 
            .I3(n23398), .O(n7794[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_8 (.CI(n23398), .I0(n7815[5]), .I1(n524_adj_4527), 
            .CO(n23399));
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4571));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3513_7_lut (.I0(GND_net), .I1(n7815[4]), .I2(n451_adj_4526), 
            .I3(n23397), .O(n7794[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4570));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3513_7 (.CI(n23397), .I0(n7815[4]), .I1(n451_adj_4526), 
            .CO(n23398));
    SB_LUT4 add_3513_6_lut (.I0(GND_net), .I1(n7815[3]), .I2(n378_adj_4525), 
            .I3(n23396), .O(n7794[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_6 (.CI(n23396), .I0(n7815[3]), .I1(n378_adj_4525), 
            .CO(n23397));
    SB_LUT4 add_3513_5_lut (.I0(GND_net), .I1(n7815[2]), .I2(n305_adj_4524), 
            .I3(n23395), .O(n7794[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_5 (.CI(n23395), .I0(n7815[2]), .I1(n305_adj_4524), 
            .CO(n23396));
    SB_LUT4 add_3513_4_lut (.I0(GND_net), .I1(n7815[1]), .I2(n232_adj_4523), 
            .I3(n23394), .O(n7794[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4569));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3513_4 (.CI(n23394), .I0(n7815[1]), .I1(n232_adj_4523), 
            .CO(n23395));
    SB_LUT4 add_3513_3_lut (.I0(GND_net), .I1(n7815[0]), .I2(n159_adj_4522), 
            .I3(n23393), .O(n7794[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3513_3 (.CI(n23393), .I0(n7815[0]), .I1(n159_adj_4522), 
            .CO(n23394));
    SB_LUT4 add_3513_2_lut (.I0(GND_net), .I1(n17_adj_4521), .I2(n86_adj_4520), 
            .I3(GND_net), .O(n7794[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3513_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4568));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4567));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4566));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3513_2 (.CI(GND_net), .I0(n17_adj_4521), .I1(n86_adj_4520), 
            .CO(n23393));
    SB_LUT4 add_3512_21_lut (.I0(GND_net), .I1(n7794[18]), .I2(GND_net), 
            .I3(n23392), .O(n7772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3512_20_lut (.I0(GND_net), .I1(n7794[17]), .I2(GND_net), 
            .I3(n23391), .O(n7772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3512_20 (.CI(n23391), .I0(n7794[17]), .I1(GND_net), .CO(n23392));
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4565));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1[23]), .I3(n22488), .O(\PID_CONTROLLER.err_23__N_3556 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4564));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4563));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4204));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4562));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1[22]), .I3(n22487), .O(\PID_CONTROLLER.err_23__N_3556 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3512_19_lut (.I0(GND_net), .I1(n7794[16]), .I2(GND_net), 
            .I3(n23390), .O(n7772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3512_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4561));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n22487), .I0(motor_state[22]), 
            .I1(n1[22]), .CO(n22488));
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4560));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4559));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1[21]), .I3(n22486), .O(\PID_CONTROLLER.err_23__N_3556 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n22486), .I0(motor_state[21]), 
            .I1(n1[21]), .CO(n22487));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1[20]), .I3(n22485), .O(\PID_CONTROLLER.err_23__N_3556 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n22485), .I0(motor_state[20]), 
            .I1(n1[20]), .CO(n22486));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1[19]), .I3(n22484), .O(\PID_CONTROLLER.err_23__N_3556 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (data_o, GND_net, encoder1_position, 
            clk32MHz, n28888, reg_B, ENCODER1_A_c_1, VCC_net, ENCODER1_B_c_0, 
            n16185, n15699) /* synthesis syn_module_defined=1 */ ;
    output [1:0]data_o;
    input GND_net;
    output [23:0]encoder1_position;
    input clk32MHz;
    output n28888;
    output [1:0]reg_B;
    input ENCODER1_A_c_1;
    input VCC_net;
    input ENCODER1_B_c_0;
    input n16185;
    input n15699;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire B_delayed, count_direction;
    wire [23:0]n2806;
    
    wire count_enable, A_delayed, n2791, n22512, n22511, n22510, 
        n22509, n22508, n22507, n22506, n22505, n22504, n22503, 
        n22502, n22501, n22500, n22499, n22498, n22497, n22496, 
        n22495, n22494, n22493, n22492, n22491, n22490, n22489;
    
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_584_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2791), 
            .I3(n22512), .O(n2806[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_584_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2791), 
            .I3(n22511), .O(n2806[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_24 (.CI(n22511), .I0(encoder1_position[22]), .I1(n2791), 
            .CO(n22512));
    SB_LUT4 add_584_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2791), 
            .I3(n22510), .O(n2806[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_23 (.CI(n22510), .I0(encoder1_position[21]), .I1(n2791), 
            .CO(n22511));
    SB_LUT4 add_584_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2791), 
            .I3(n22509), .O(n2806[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_22 (.CI(n22509), .I0(encoder1_position[20]), .I1(n2791), 
            .CO(n22510));
    SB_LUT4 add_584_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2791), 
            .I3(n22508), .O(n2806[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_21 (.CI(n22508), .I0(encoder1_position[19]), .I1(n2791), 
            .CO(n22509));
    SB_LUT4 add_584_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2791), 
            .I3(n22507), .O(n2806[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_20 (.CI(n22507), .I0(encoder1_position[18]), .I1(n2791), 
            .CO(n22508));
    SB_LUT4 add_584_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2791), 
            .I3(n22506), .O(n2806[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_19 (.CI(n22506), .I0(encoder1_position[17]), .I1(n2791), 
            .CO(n22507));
    SB_LUT4 add_584_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2791), 
            .I3(n22505), .O(n2806[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_18 (.CI(n22505), .I0(encoder1_position[16]), .I1(n2791), 
            .CO(n22506));
    SB_LUT4 add_584_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2791), 
            .I3(n22504), .O(n2806[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_17 (.CI(n22504), .I0(encoder1_position[15]), .I1(n2791), 
            .CO(n22505));
    SB_LUT4 add_584_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2791), 
            .I3(n22503), .O(n2806[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_16 (.CI(n22503), .I0(encoder1_position[14]), .I1(n2791), 
            .CO(n22504));
    SB_LUT4 add_584_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2791), 
            .I3(n22502), .O(n2806[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_15 (.CI(n22502), .I0(encoder1_position[13]), .I1(n2791), 
            .CO(n22503));
    SB_LUT4 add_584_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2791), 
            .I3(n22501), .O(n2806[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_14 (.CI(n22501), .I0(encoder1_position[12]), .I1(n2791), 
            .CO(n22502));
    SB_LUT4 add_584_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2791), 
            .I3(n22500), .O(n2806[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_13 (.CI(n22500), .I0(encoder1_position[11]), .I1(n2791), 
            .CO(n22501));
    SB_LUT4 add_584_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2791), 
            .I3(n22499), .O(n2806[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_12 (.CI(n22499), .I0(encoder1_position[10]), .I1(n2791), 
            .CO(n22500));
    SB_LUT4 add_584_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2791), 
            .I3(n22498), .O(n2806[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_11 (.CI(n22498), .I0(encoder1_position[9]), .I1(n2791), 
            .CO(n22499));
    SB_LUT4 add_584_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2791), 
            .I3(n22497), .O(n2806[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_10 (.CI(n22497), .I0(encoder1_position[8]), .I1(n2791), 
            .CO(n22498));
    SB_LUT4 add_584_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2791), 
            .I3(n22496), .O(n2806[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2806[23]));   // quad.v(35[10] 41[6])
    SB_CARRY add_584_9 (.CI(n22496), .I0(encoder1_position[7]), .I1(n2791), 
            .CO(n22497));
    SB_LUT4 add_584_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2791), 
            .I3(n22495), .O(n2806[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_8 (.CI(n22495), .I0(encoder1_position[6]), .I1(n2791), 
            .CO(n22496));
    SB_LUT4 add_584_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2791), 
            .I3(n22494), .O(n2806[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_7 (.CI(n22494), .I0(encoder1_position[5]), .I1(n2791), 
            .CO(n22495));
    SB_LUT4 add_584_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2791), 
            .I3(n22493), .O(n2806[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_6 (.CI(n22493), .I0(encoder1_position[4]), .I1(n2791), 
            .CO(n22494));
    SB_LUT4 add_584_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2791), 
            .I3(n22492), .O(n2806[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_5 (.CI(n22492), .I0(encoder1_position[3]), .I1(n2791), 
            .CO(n22493));
    SB_LUT4 add_584_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2791), 
            .I3(n22491), .O(n2806[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_4 (.CI(n22491), .I0(encoder1_position[2]), .I1(n2791), 
            .CO(n22492));
    SB_LUT4 add_584_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2791), 
            .I3(n22490), .O(n2806[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_3 (.CI(n22490), .I0(encoder1_position[1]), .I1(n2791), 
            .CO(n22491));
    SB_LUT4 add_584_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n22489), .O(n2806[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_584_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_584_2 (.CI(n22489), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n22490));
    SB_LUT4 i912_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2791));   // quad.v(37[5] 40[8])
    defparam i912_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_584_1 (.CI(GND_net), .I0(n2791), .I1(n2791), .CO(n22489));
    \grp_debouncer(2,100)  debounce (.n28888(n28888), .reg_B({reg_B}), .GND_net(GND_net), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .ENCODER1_B_c_0(ENCODER1_B_c_0), .n16185(n16185), .data_o({data_o}), 
            .n15699(n15699));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (n28888, reg_B, GND_net, ENCODER1_A_c_1, 
            clk32MHz, VCC_net, ENCODER1_B_c_0, n16185, data_o, n15699);
    output n28888;
    output [1:0]reg_B;
    input GND_net;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input VCC_net;
    input ENCODER1_B_c_0;
    input n16185;
    output [1:0]data_o;
    input n15699;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3740;
    wire [6:0]n33;
    
    wire n22873, n22872, n22871, n22870, n22869, n22868;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n28888));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n28888), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1215__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 cnt_reg_1215_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n22873), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1215_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n22872), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1215_add_4_7 (.CI(n22872), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n22873));
    SB_LUT4 cnt_reg_1215_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n22871), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1215_add_4_6 (.CI(n22871), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n22872));
    SB_LUT4 cnt_reg_1215_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n22870), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1215_add_4_5 (.CI(n22870), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n22871));
    SB_LUT4 cnt_reg_1215_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n22869), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1215_add_4_4 (.CI(n22869), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n22870));
    SB_LUT4 cnt_reg_1215_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n22868), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1215_add_4_3 (.CI(n22868), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n22869));
    SB_LUT4 cnt_reg_1215_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1215_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1215_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n22868));
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n16185));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n15699));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1215__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1215__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1215__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1215__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1215__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1215__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3740));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,8000000,23,1) 
//

module \pwm(32000000,20000,8000000,23,1)  (INHA_c_0, clk32MHz, \half_duty_new[0] , 
            n15460, \half_duty[0][0] , GND_net, \half_duty[0][1] , \half_duty[0][2] , 
            \half_duty[0][3] , \half_duty[0][4] , \half_duty[0][5] , \half_duty[0][6] , 
            \half_duty[0][7] , VCC_net, pwm_setpoint, \half_duty_new[1] , 
            \half_duty_new[2] , \half_duty_new[3] , \half_duty_new[4] , 
            \half_duty_new[5] , \half_duty_new[6] , \half_duty_new[7] , 
            n16195, n16194, n16193, n16192, n16191, n16190, n16189, 
            n15700);
    output INHA_c_0;
    input clk32MHz;
    output \half_duty_new[0] ;
    output n15460;
    output \half_duty[0][0] ;
    input GND_net;
    output \half_duty[0][1] ;
    output \half_duty[0][2] ;
    output \half_duty[0][3] ;
    output \half_duty[0][4] ;
    output \half_duty[0][5] ;
    output \half_duty[0][6] ;
    output \half_duty[0][7] ;
    input VCC_net;
    input [22:0]pwm_setpoint;
    output \half_duty_new[1] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[5] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n16195;
    input n16194;
    input n16193;
    input n16192;
    input n16191;
    input n16190;
    input n16189;
    input n15700;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n18721, n15462;
    wire [9:0]half_duty_new_9__N_678;
    wire [10:0]n49;
    
    wire pwm_out_0__N_621;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    wire [2:0]n125;
    
    wire n15430;
    wire [2:0]\pause_counter[0] ;   // vhdl/pwm.vhd(52[11:24])
    
    wire n15602;
    wire [10:0]pwm_out_0__N_597;
    
    wire n22351, pwm_out_0__N_596, n22350, n10, n22349, n9, n22348, 
        n8, n22347, n7, n22346, n6, n22345, n5, n22344;
    wire [2:0]pause_counter_0__2__N_672;
    
    wire n4, n22343;
    wire [22:0]n5413;
    
    wire n22682, n22681, n22680, n22679, n22678, n3, n22342, n22677, 
        n22676, n2, n22341, n22675, n22674, n22673, n22672, n22671, 
        n22670, n22669, n12, n28931, n10_adj_4176, n22668, n22667, 
        n22666, n22665, n22664, n22663, n22662, n22661, n22660, 
        n22659, n22658, n1, n22657, n22656, n22655, n22654, n22653, 
        n22652, n22651, n22650, n21, n22649, n22648, n22647, n22646, 
        n22645, n22644, n22643, n22642, n22641, n22640, n15582, 
        n22823, n22822, n22821, n22820, n22819, n22818, n22817, 
        n22816, n22815, n22814, n15, n14, n13, n17, n19, n29009, 
        n29069, n21_adj_4177, n23;
    
    SB_DFFE pwm_out_0__40 (.Q(INHA_c_0), .C(clk32MHz), .E(n15462), .D(n18721));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(clk32MHz), .D(half_duty_new_9__N_678[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1208__i10 (.Q(\count[0] [10]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[10]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i9 (.Q(\count[0] [9]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[9]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i8 (.Q(\count[0] [8]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[8]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i7 (.Q(\count[0] [7]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[7]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i6 (.Q(\count[0] [6]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[6]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i5 (.Q(\count[0] [5]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[5]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i4 (.Q(\count[0] [4]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[4]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i3 (.Q(\count[0] [3]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[3]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i2 (.Q(\count[0] [2]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[2]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1208__i1 (.Q(\count[0] [1]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[1]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR pause_counter_0__i2 (.Q(\pause_counter[0] [2]), .C(clk32MHz), 
            .E(n15430), .D(n125[2]), .R(n15602));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR pause_counter_0__i1 (.Q(\pause_counter[0] [1]), .C(clk32MHz), 
            .E(n15430), .D(n125[1]), .R(n15602));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0][5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i7_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[6]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_597[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY pwm_out_0__I_20_13 (.CI(n22351), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_596));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n22350), .I0(VCC_net), .I1(VCC_net), 
            .CO(n22351));
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n22349), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n22349), .I0(VCC_net), .I1(VCC_net), 
            .CO(n22350));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n22348), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_10 (.CI(n22348), .I0(GND_net), .I1(VCC_net), 
            .CO(n22349));
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_597[7]), 
            .I3(n22347), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_9 (.CI(n22347), .I0(GND_net), .I1(pwm_out_0__N_597[7]), 
            .CO(n22348));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_597[6]), 
            .I3(n22346), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n22346), .I0(VCC_net), .I1(pwm_out_0__N_597[6]), 
            .CO(n22347));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_597[5]), 
            .I3(n22345), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_DFFESR count_0__1208__i0 (.Q(\count[0] [0]), .C(clk32MHz), .E(pwm_out_0__N_621), 
            .D(n49[0]), .R(n15460));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY pwm_out_0__I_20_7 (.CI(n22345), .I0(GND_net), .I1(pwm_out_0__N_597[5]), 
            .CO(n22346));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_597[4]), 
            .I3(n22344), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n22344), .I0(GND_net), .I1(pwm_out_0__N_597[4]), 
            .CO(n22345));
    SB_LUT4 i14076_3_lut_3_lut (.I0(\pause_counter[0] [0]), .I1(\pause_counter[0] [1]), 
            .I2(\pause_counter[0] [2]), .I3(GND_net), .O(pause_counter_0__2__N_672[0]));   // vhdl/pwm.vhd(72[7:27])
    defparam i14076_3_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i24742_2_lut_3_lut (.I0(\pause_counter[0] [0]), .I1(\pause_counter[0] [1]), 
            .I2(\pause_counter[0] [2]), .I3(GND_net), .O(pwm_out_0__N_621));   // vhdl/pwm.vhd(72[7:27])
    defparam i24742_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_597[3]), 
            .I3(n22343), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_1670_24_lut (.I0(GND_net), .I1(n5413[22]), .I2(pwm_setpoint[22]), 
            .I3(n22682), .O(half_duty_new_9__N_678[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1670_23_lut (.I0(GND_net), .I1(n5413[21]), .I2(pwm_setpoint[21]), 
            .I3(n22681), .O(half_duty_new_9__N_678[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1670_23 (.CI(n22681), .I0(n5413[21]), .I1(pwm_setpoint[21]), 
            .CO(n22682));
    SB_LUT4 add_1670_22_lut (.I0(GND_net), .I1(n5413[20]), .I2(pwm_setpoint[20]), 
            .I3(n22680), .O(half_duty_new_9__N_678[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1670_22 (.CI(n22680), .I0(n5413[20]), .I1(pwm_setpoint[20]), 
            .CO(n22681));
    SB_CARRY pwm_out_0__I_20_5 (.CI(n22343), .I0(GND_net), .I1(pwm_out_0__N_597[3]), 
            .CO(n22344));
    SB_LUT4 add_1670_21_lut (.I0(GND_net), .I1(n5413[19]), .I2(pwm_setpoint[19]), 
            .I3(n22679), .O(half_duty_new_9__N_678[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1670_21 (.CI(n22679), .I0(n5413[19]), .I1(pwm_setpoint[19]), 
            .CO(n22680));
    SB_LUT4 add_1670_20_lut (.I0(GND_net), .I1(n5413[18]), .I2(pwm_setpoint[18]), 
            .I3(n22678), .O(half_duty_new_9__N_678[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1670_20 (.CI(n22678), .I0(n5413[18]), .I1(pwm_setpoint[18]), 
            .CO(n22679));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_597[2]), 
            .I3(n22342), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_1670_19_lut (.I0(GND_net), .I1(n5413[17]), .I2(pwm_setpoint[17]), 
            .I3(n22677), .O(half_duty_new_9__N_678[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1670_19 (.CI(n22677), .I0(n5413[17]), .I1(pwm_setpoint[17]), 
            .CO(n22678));
    SB_CARRY pwm_out_0__I_20_4 (.CI(n22342), .I0(GND_net), .I1(pwm_out_0__N_597[2]), 
            .CO(n22343));
    SB_LUT4 add_1670_18_lut (.I0(GND_net), .I1(n5413[16]), .I2(pwm_setpoint[16]), 
            .I3(n22676), .O(half_duty_new_9__N_678[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_597[1]), 
            .I3(n22341), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_1670_18 (.CI(n22676), .I0(n5413[16]), .I1(pwm_setpoint[16]), 
            .CO(n22677));
    SB_LUT4 add_1670_17_lut (.I0(GND_net), .I1(n5413[15]), .I2(pwm_setpoint[15]), 
            .I3(n22675), .O(half_duty_new_9__N_678[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1670_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1670_17 (.CI(n22675), .I0(n5413[15]), .I1(pwm_setpoint[15]), 
            .CO(n22676));
    SB_CARRY add_1670_16 (.CI(n22674), .I0(n5413[14]), .I1(pwm_setpoint[14]), 
            .CO(n22675));
    SB_CARRY add_1670_15 (.CI(n22673), .I0(n5413[13]), .I1(pwm_setpoint[13]), 
            .CO(n22674));
    SB_CARRY add_1670_14 (.CI(n22672), .I0(n5413[12]), .I1(pwm_setpoint[12]), 
            .CO(n22673));
    SB_CARRY add_1670_13 (.CI(n22671), .I0(n5413[11]), .I1(pwm_setpoint[11]), 
            .CO(n22672));
    SB_CARRY add_1670_12 (.CI(n22670), .I0(n5413[10]), .I1(pwm_setpoint[10]), 
            .CO(n22671));
    SB_CARRY pwm_out_0__I_20_3 (.CI(n22341), .I0(GND_net), .I1(pwm_out_0__N_597[1]), 
            .CO(n22342));
    SB_CARRY add_1670_11 (.CI(n22669), .I0(n5413[9]), .I1(pwm_setpoint[9]), 
            .CO(n22670));
    SB_LUT4 i5_4_lut (.I0(\count[0] [10]), .I1(\count[0] [6]), .I2(\count[0] [7]), 
            .I3(\count[0] [0]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i6_4_lut (.I0(\count[0] [3]), .I1(n12), .I2(\count[0] [8]), 
            .I3(\count[0] [4]), .O(n28931));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i4_4_lut (.I0(pwm_out_0__N_621), .I1(n28931), .I2(\count[0] [1]), 
            .I3(\count[0] [5]), .O(n10_adj_4176));
    defparam i4_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i24744_3_lut (.I0(\count[0] [2]), .I1(n10_adj_4176), .I2(\count[0] [9]), 
            .I3(GND_net), .O(n15460));
    defparam i24744_3_lut.LUT_INIT = 16'h2020;
    SB_CARRY add_1670_10 (.CI(n22668), .I0(n5413[8]), .I1(pwm_setpoint[8]), 
            .CO(n22669));
    SB_CARRY add_1670_9 (.CI(n22667), .I0(n5413[7]), .I1(pwm_setpoint[7]), 
            .CO(n22668));
    SB_CARRY add_1670_8 (.CI(n22666), .I0(n5413[6]), .I1(pwm_setpoint[6]), 
            .CO(n22667));
    SB_CARRY add_1670_7 (.CI(n22665), .I0(n5413[5]), .I1(pwm_setpoint[5]), 
            .CO(n22666));
    SB_CARRY add_1670_6 (.CI(n22664), .I0(n5413[4]), .I1(pwm_setpoint[4]), 
            .CO(n22665));
    SB_CARRY add_1670_5 (.CI(n22663), .I0(n5413[3]), .I1(pwm_setpoint[3]), 
            .CO(n22664));
    SB_CARRY add_1670_4 (.CI(n22662), .I0(n5413[2]), .I1(pwm_setpoint[2]), 
            .CO(n22663));
    SB_CARRY add_1670_3 (.CI(n22661), .I0(n5413[1]), .I1(pwm_setpoint[1]), 
            .CO(n22662));
    SB_CARRY add_1670_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n22661));
    SB_LUT4 add_1677_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n22660), .O(n5413[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1677_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n22659), .O(n5413[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_22 (.CI(n22659), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n22660));
    SB_LUT4 add_1677_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n22658), .O(n5413[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_597[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_1677_21 (.CI(n22658), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n22659));
    SB_LUT4 add_1677_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n22657), .O(n5413[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_597[0]), 
            .CO(n22341));
    SB_CARRY add_1677_20 (.CI(n22657), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n22658));
    SB_LUT4 add_1677_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n22656), .O(n5413[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_19 (.CI(n22656), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n22657));
    SB_LUT4 add_1677_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n22655), .O(n5413[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_18 (.CI(n22655), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n22656));
    SB_LUT4 add_1677_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n22654), .O(n5413[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_17 (.CI(n22654), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n22655));
    SB_LUT4 add_1677_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n22653), .O(n5413[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_16 (.CI(n22653), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n22654));
    SB_LUT4 add_1677_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n22652), .O(n5413[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_15 (.CI(n22652), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n22653));
    SB_LUT4 add_1677_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n22651), .O(n5413[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_14 (.CI(n22651), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n22652));
    SB_LUT4 add_1677_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n22650), .O(n5413[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1280_2_lut (.I0(\pause_counter[0] [1]), .I1(\pause_counter[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n125[1]));   // vhdl/pwm.vhd(89[25:41])
    defparam i1280_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(n21), .I1(pwm_out_0__N_621), .I2(GND_net), .I3(GND_net), 
            .O(n15430));
    defparam i1_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1287_3_lut (.I0(\pause_counter[0] [2]), .I1(\pause_counter[0] [1]), 
            .I2(\pause_counter[0] [0]), .I3(GND_net), .O(n125[2]));   // vhdl/pwm.vhd(89[25:41])
    defparam i1287_3_lut.LUT_INIT = 16'h6a6a;
    SB_CARRY add_1677_13 (.CI(n22650), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n22651));
    SB_LUT4 add_1677_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n22649), .O(n5413[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_12 (.CI(n22649), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n22650));
    SB_LUT4 add_1677_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n22648), .O(n5413[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_11 (.CI(n22648), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n22649));
    SB_LUT4 add_1677_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n22647), .O(n5413[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_10 (.CI(n22647), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n22648));
    SB_LUT4 add_1677_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n22646), .O(n5413[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_9 (.CI(n22646), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n22647));
    SB_LUT4 add_1677_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n22645), .O(n5413[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_8 (.CI(n22645), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n22646));
    SB_LUT4 add_1677_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n22644), .O(n5413[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_7 (.CI(n22644), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n22645));
    SB_LUT4 add_1677_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n22643), .O(n5413[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_6 (.CI(n22643), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n22644));
    SB_LUT4 add_1677_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n22642), .O(n5413[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_5 (.CI(n22642), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n22643));
    SB_LUT4 add_1677_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n22641), .O(n5413[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_4 (.CI(n22641), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n22642));
    SB_LUT4 add_1677_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n22640), .O(n5413[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_3 (.CI(n22640), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n22641));
    SB_LUT4 add_1677_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5413[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1677_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1677_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n22640));
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(clk32MHz), .D(half_duty_new_9__N_678[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(clk32MHz), .D(half_duty_new_9__N_678[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(clk32MHz), .D(half_duty_new_9__N_678[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(clk32MHz), .D(half_duty_new_9__N_678[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(\half_duty_new[5] ), .C(clk32MHz), .D(half_duty_new_9__N_678[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(clk32MHz), .D(half_duty_new_9__N_678[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(clk32MHz), .D(half_duty_new_9__N_678[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESS pause_counter_0__i0 (.Q(\pause_counter[0] [0]), .C(clk32MHz), 
            .E(n15430), .D(pause_counter_0__2__N_672[0]), .S(n15582));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i21460_1_lut_2_lut (.I0(n21), .I1(pwm_out_0__N_621), .I2(GND_net), 
            .I3(GND_net), .O(n15582));
    defparam i21460_1_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 count_0__1208_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n22823), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1208_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n22822), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_11 (.CI(n22822), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n22823));
    SB_LUT4 count_0__1208_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n22821), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_10 (.CI(n22821), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n22822));
    SB_LUT4 count_0__1208_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n22820), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_9 (.CI(n22820), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n22821));
    SB_LUT4 count_0__1208_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n22819), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_8 (.CI(n22819), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n22820));
    SB_LUT4 count_0__1208_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n22818), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_7 (.CI(n22818), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n22819));
    SB_LUT4 count_0__1208_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n22817), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_6 (.CI(n22817), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n22818));
    SB_LUT4 count_0__1208_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n22816), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_5 (.CI(n22816), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n22817));
    SB_LUT4 count_0__1208_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n22815), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_4 (.CI(n22815), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n22816));
    SB_LUT4 count_0__1208_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n22814), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_3 (.CI(n22814), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n22815));
    SB_LUT4 count_0__1208_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1208_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1208_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n22814));
    SB_LUT4 i4_4_lut_adj_1479 (.I0(\half_duty[0][3] ), .I1(\half_duty[0][5] ), 
            .I2(\count[0] [3]), .I3(\count[0] [5]), .O(n15));   // vhdl/pwm.vhd(80[8:31])
    defparam i4_4_lut_adj_1479.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(\half_duty[0][2] ), .I1(\half_duty[0][4] ), .I2(\count[0] [2]), 
            .I3(\count[0] [4]), .O(n14));   // vhdl/pwm.vhd(80[8:31])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut (.I0(\half_duty[0][7] ), .I1(\half_duty[0][1] ), .I2(\count[0] [7]), 
            .I3(\count[0] [1]), .O(n13));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i6_4_lut_adj_1480 (.I0(\count[0] [10]), .I1(\count[0] [9]), 
            .I2(\half_duty[0][0] ), .I3(\count[0] [0]), .O(n17));   // vhdl/pwm.vhd(80[8:31])
    defparam i6_4_lut_adj_1480.LUT_INIT = 16'heffe;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(\half_duty[0][6] ), .I2(\count[0] [8]), 
            .I3(\count[0] [6]), .O(n19));   // vhdl/pwm.vhd(80[8:31])
    defparam i8_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i10_4_lut (.I0(n19), .I1(n17), .I2(n13), .I3(n14), .O(n21));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23158_2_lut (.I0(n1), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n29009));
    defparam i23158_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23217_4_lut (.I0(n4), .I1(n7), .I2(n5), .I3(n10), .O(n29069));
    defparam i23217_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1481 (.I0(\count[0] [10]), .I1(n9), .I2(n8), 
            .I3(n2), .O(n21_adj_4177));
    defparam i8_4_lut_adj_1481.LUT_INIT = 16'h0002;
    SB_LUT4 i10_4_lut_adj_1482 (.I0(n29009), .I1(pwm_out_0__N_596), .I2(n6), 
            .I3(pwm_out_0__N_621), .O(n23));
    defparam i10_4_lut_adj_1482.LUT_INIT = 16'h0400;
    SB_LUT4 i1_4_lut (.I0(n23), .I1(n18721), .I2(n21_adj_4177), .I3(n29069), 
            .O(n15462));
    defparam i1_4_lut.LUT_INIT = 16'h33b3;
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(clk32MHz), .D(n16195));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(clk32MHz), .D(n16194));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0][5] ), .C(clk32MHz), .D(n16193));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(clk32MHz), .D(n16192));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(clk32MHz), .D(n16191));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(clk32MHz), .D(n16190));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(clk32MHz), .D(n16189));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i11027_2_lut_3_lut_4_lut (.I0(\pause_counter[0] [0]), .I1(\pause_counter[0] [1]), 
            .I2(n21), .I3(pwm_out_0__N_621), .O(n15602));   // vhdl/pwm.vhd(72[7:27])
    defparam i11027_2_lut_3_lut_4_lut.LUT_INIT = 16'h0111;
    SB_LUT4 i14156_2_lut (.I0(n21), .I1(pwm_out_0__N_621), .I2(GND_net), 
            .I3(GND_net), .O(n18721));
    defparam i14156_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(clk32MHz), .D(n15700));   // vhdl/pwm.vhd(59[5] 95[12])
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_out_frame[16] , \data_out_frame[17] , GND_net, \data_out_frame[18] , 
            \data_out_frame[19] , \data_out_frame[23] , n15762, \data_in[3] , 
            clk32MHz, \data_out_frame[24] , \data_out_frame[20] , n15761, 
            \data_out_frame[13] , \data_out_frame[15] , n15760, \data_in[2] , 
            \data_out_frame[25] , setpoint, n15759, \data_out_frame[5] , 
            \data_out_frame[6] , \data_out_frame[7] , n15758, n15757, 
            \data_out_frame[14] , \data_out_frame[12] , \data_out_frame[10] , 
            \data_out_frame[11] , \data_out_frame[9] , \data_out_frame[8] , 
            n15756, n15755, rx_data, \data_in_frame[9] , n15754, n15753, 
            \data_in_frame[1] , \data_in_frame[2] , \data_in_frame[3] , 
            n15752, \data_in[1] , \data_in_frame[4] , \data_in_frame[5] , 
            \data_in_frame[8] , \data_in_frame[6] , n15751, rx_data_ready, 
            n15750, n15749, n15748, n15747, n14288, n771, n9520, 
            n4609, \FRAME_MATCHER.state[0] , n14253, n123, n63, n26561, 
            n14291, n4677, n14254, \FRAME_MATCHER.state[3] , \data_in_frame[12] , 
            \data_in_frame[13] , \data_in_frame[10] , n15746, \FRAME_MATCHER.state_31__N_2672[1] , 
            n8595, n122, \FRAME_MATCHER.state_31__N_2672[2] , n4452, 
            n7, n2649, n8, n14279, n15745, \data_in_frame[11] , 
            tx_active, n15744, \data_in[0] , n15743, n15742, n27362, 
            n4772, n15741, LED_c, n27374, n15740, n15739, n15738, 
            n15737, IntegralLimit, n15736, n15735, n15734, n15733, 
            n15732, n15731, n15730, n15729, n15728, n15727, n15726, 
            n15725, n15724, n15723, n15722, n15721, n15720, n15719, 
            n15718, n15717, n15716, n15715, n63_adj_3, n27965, n25997, 
            DE_c, n31238, n31239, n16178, PWMLimit, n16177, n16176, 
            n16175, n16174, n16173, n16172, n16171, n16170, n16169, 
            n16168, n16167, n16166, n16165, n16164, n16163, n16162, 
            n16161, n16160, n16159, n16158, n16157, n16156, n16155, 
            control_mode, n16154, n16153, n16152, n16151, n16150, 
            n16149, n15973, neopxl_color, n15972, n15971, n15970, 
            n15969, n15968, n15967, n15966, n15965, n15964, n15963, 
            n15962, n15961, n15960, n15959, n15958, n15957, n15956, 
            n15955, n15954, n15953, n15952, n15951, n15950, n15949, 
            n15948, n15947, n15946, n15945, n15944, n15943, n15942, 
            n15941, n15940, n15939, n15938, n15937, n15936, n15935, 
            n15934, n15933, n15932, n15931, n15930, n15929, n15928, 
            n15927, n15926, n15925, n15924, n15923, n15922, n15921, 
            n15920, n15919, n15918, n15917, n15916, n15915, n15914, 
            n15913, n15912, n15911, n15910, n15909, n15908, n15907, 
            n15906, n15905, n15904, n15903, n15902, n15901, n15900, 
            n15899, n15898, n15897, n15896, n15895, n15894, n15893, 
            n15892, n15891, n15890, n15889, n15888, n15887, n15886, 
            n15885, n15884, n15883, n15882, n15881, n25861, n15695, 
            n15880, n15879, n15878, n15877, n15876, n15875, n15874, 
            n15873, n15872, n15871, n15870, n15869, n15868, n15867, 
            n15866, n15865, n15864, n15863, n15862, n15861, n15860, 
            n15859, n15858, n15857, n15856, n15855, n15854, n15853, 
            n15852, n15851, n15850, n15849, n15848, n15694, n15692, 
            n15691, \Ki[0] , n15690, \Kp[0] , n15689, n15847, n15846, 
            n15845, n15844, n15843, n15842, n15841, n15682, n15840, 
            n15839, n15838, n15837, n15836, n15835, n15834, n15833, 
            n15832, n15831, n15830, n15829, n15828, n15827, n15826, 
            n15825, n15824, n15823, n15822, n15821, n15820, n15819, 
            n15818, n15817, n11648, n4774, n15816, n15815, n15814, 
            n15813, n15812, n15811, n15810, n15809, n15808, n15807, 
            n15806, n15805, n15804, n15803, n15802, n15801, n15800, 
            n15799, n15798, \Ki[15] , n15797, \Ki[14] , n15796, 
            \Ki[13] , n15795, \Ki[12] , n15794, \Ki[11] , n15793, 
            \Ki[10] , n15792, \Ki[9] , n15791, \Ki[8] , n15790, 
            \Ki[7] , n15789, \Ki[6] , n15788, \Ki[5] , n15787, \Ki[4] , 
            n15786, \Ki[3] , n15785, \Ki[2] , n15784, \Ki[1] , n15783, 
            \Kp[15] , n15782, \Kp[14] , n15781, \Kp[13] , n15780, 
            \Kp[12] , n15779, \Kp[11] , n15778, \Kp[10] , n15777, 
            \Kp[9] , n15776, \Kp[8] , n15775, \Kp[7] , n15774, \Kp[6] , 
            n15773, \Kp[5] , n15772, \Kp[4] , n15771, \Kp[3] , n15770, 
            \Kp[2] , n15769, \Kp[1] , n15768, n15767, n15766, n15765, 
            n15764, n15763, \r_Bit_Index[0] , tx_o, r_SM_Main, \r_SM_Main_2__N_3497[1] , 
            n27464, n27476, n4, VCC_net, n15704, n8439, n31237, 
            n15698, tx_enable, \r_SM_Main_2__N_3426[2] , r_SM_Main_adj_11, 
            n26557, \r_Bit_Index[0]_adj_7 , r_Rx_Data, RX_N_2, n14264, 
            n18753, n14259, n4_adj_8, n15508, n15619, n4_adj_9, 
            n4_adj_10, n15711, n16227, n15707, n26153, n15686, n15685, 
            n15684, n15683, n15681, n15680) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    input GND_net;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[23] ;
    input n15762;
    output [7:0]\data_in[3] ;
    input clk32MHz;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_out_frame[20] ;
    input n15761;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[15] ;
    input n15760;
    output [7:0]\data_in[2] ;
    output [7:0]\data_out_frame[25] ;
    output [23:0]setpoint;
    input n15759;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    input n15758;
    input n15757;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[8] ;
    input n15756;
    input n15755;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[9] ;
    input n15754;
    input n15753;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[3] ;
    input n15752;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[6] ;
    input n15751;
    output rx_data_ready;
    input n15750;
    input n15749;
    input n15748;
    input n15747;
    output n14288;
    output n771;
    output n9520;
    output n4609;
    output \FRAME_MATCHER.state[0] ;
    output n14253;
    output n123;
    output n63;
    output n26561;
    output n14291;
    output n4677;
    output n14254;
    output \FRAME_MATCHER.state[3] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[10] ;
    input n15746;
    output \FRAME_MATCHER.state_31__N_2672[1] ;
    output n8595;
    output n122;
    output \FRAME_MATCHER.state_31__N_2672[2] ;
    output n4452;
    output n7;
    output n2649;
    output n8;
    output n14279;
    input n15745;
    output [7:0]\data_in_frame[11] ;
    output tx_active;
    input n15744;
    output [7:0]\data_in[0] ;
    input n15743;
    input n15742;
    input n27362;
    output n4772;
    input n15741;
    output LED_c;
    output n27374;
    input n15740;
    input n15739;
    input n15738;
    input n15737;
    output [23:0]IntegralLimit;
    input n15736;
    input n15735;
    input n15734;
    input n15733;
    input n15732;
    input n15731;
    input n15730;
    input n15729;
    input n15728;
    input n15727;
    input n15726;
    input n15725;
    input n15724;
    input n15723;
    input n15722;
    input n15721;
    input n15720;
    input n15719;
    input n15718;
    input n15717;
    input n15716;
    input n15715;
    input n63_adj_3;
    output n27965;
    input n25997;
    output DE_c;
    input n31238;
    input n31239;
    input n16178;
    output [23:0]PWMLimit;
    input n16177;
    input n16176;
    input n16175;
    input n16174;
    input n16173;
    input n16172;
    input n16171;
    input n16170;
    input n16169;
    input n16168;
    input n16167;
    input n16166;
    input n16165;
    input n16164;
    input n16163;
    input n16162;
    input n16161;
    input n16160;
    input n16159;
    input n16158;
    input n16157;
    input n16156;
    input n16155;
    output [7:0]control_mode;
    input n16154;
    input n16153;
    input n16152;
    input n16151;
    input n16150;
    input n16149;
    input n15973;
    output [23:0]neopxl_color;
    input n15972;
    input n15971;
    input n15970;
    input n15969;
    input n15968;
    input n15967;
    input n15966;
    input n15965;
    input n15964;
    input n15963;
    input n15962;
    input n15961;
    input n15960;
    input n15959;
    input n15958;
    input n15957;
    input n15956;
    input n15955;
    input n15954;
    input n15953;
    input n15952;
    input n15951;
    input n15950;
    input n15949;
    input n15948;
    input n15947;
    input n15946;
    input n15945;
    input n15944;
    input n15943;
    input n15942;
    input n15941;
    input n15940;
    input n15939;
    input n15938;
    input n15937;
    input n15936;
    input n15935;
    input n15934;
    input n15933;
    input n15932;
    input n15931;
    input n15930;
    input n15929;
    input n15928;
    input n15927;
    input n15926;
    input n15925;
    input n15924;
    input n15923;
    input n15922;
    input n15921;
    input n15920;
    input n15919;
    input n15918;
    input n15917;
    input n15916;
    input n15915;
    input n15914;
    input n15913;
    input n15912;
    input n15911;
    input n15910;
    input n15909;
    input n15908;
    input n15907;
    input n15906;
    input n15905;
    input n15904;
    input n15903;
    input n15902;
    input n15901;
    input n15900;
    input n15899;
    input n15898;
    input n15897;
    input n15896;
    input n15895;
    input n15894;
    input n15893;
    input n15892;
    input n15891;
    input n15890;
    input n15889;
    input n15888;
    input n15887;
    input n15886;
    input n15885;
    input n15884;
    input n15883;
    input n15882;
    input n15881;
    input n25861;
    input n15695;
    input n15880;
    input n15879;
    input n15878;
    input n15877;
    input n15876;
    input n15875;
    input n15874;
    input n15873;
    input n15872;
    input n15871;
    input n15870;
    input n15869;
    input n15868;
    input n15867;
    input n15866;
    input n15865;
    input n15864;
    input n15863;
    input n15862;
    input n15861;
    input n15860;
    input n15859;
    input n15858;
    input n15857;
    input n15856;
    input n15855;
    input n15854;
    input n15853;
    input n15852;
    input n15851;
    input n15850;
    input n15849;
    input n15848;
    input n15694;
    input n15692;
    input n15691;
    output \Ki[0] ;
    input n15690;
    output \Kp[0] ;
    input n15689;
    input n15847;
    input n15846;
    input n15845;
    input n15844;
    input n15843;
    input n15842;
    input n15841;
    input n15682;
    input n15840;
    input n15839;
    input n15838;
    input n15837;
    input n15836;
    input n15835;
    input n15834;
    input n15833;
    input n15832;
    input n15831;
    input n15830;
    input n15829;
    input n15828;
    input n15827;
    input n15826;
    input n15825;
    input n15824;
    input n15823;
    input n15822;
    input n15821;
    input n15820;
    input n15819;
    input n15818;
    input n15817;
    output n11648;
    output n4774;
    input n15816;
    input n15815;
    input n15814;
    input n15813;
    input n15812;
    input n15811;
    input n15810;
    input n15809;
    input n15808;
    input n15807;
    input n15806;
    input n15805;
    input n15804;
    input n15803;
    input n15802;
    input n15801;
    input n15800;
    input n15799;
    input n15798;
    output \Ki[15] ;
    input n15797;
    output \Ki[14] ;
    input n15796;
    output \Ki[13] ;
    input n15795;
    output \Ki[12] ;
    input n15794;
    output \Ki[11] ;
    input n15793;
    output \Ki[10] ;
    input n15792;
    output \Ki[9] ;
    input n15791;
    output \Ki[8] ;
    input n15790;
    output \Ki[7] ;
    input n15789;
    output \Ki[6] ;
    input n15788;
    output \Ki[5] ;
    input n15787;
    output \Ki[4] ;
    input n15786;
    output \Ki[3] ;
    input n15785;
    output \Ki[2] ;
    input n15784;
    output \Ki[1] ;
    input n15783;
    output \Kp[15] ;
    input n15782;
    output \Kp[14] ;
    input n15781;
    output \Kp[13] ;
    input n15780;
    output \Kp[12] ;
    input n15779;
    output \Kp[11] ;
    input n15778;
    output \Kp[10] ;
    input n15777;
    output \Kp[9] ;
    input n15776;
    output \Kp[8] ;
    input n15775;
    output \Kp[7] ;
    input n15774;
    output \Kp[6] ;
    input n15773;
    output \Kp[5] ;
    input n15772;
    output \Kp[4] ;
    input n15771;
    output \Kp[3] ;
    input n15770;
    output \Kp[2] ;
    input n15769;
    output \Kp[1] ;
    input n15768;
    input n15767;
    input n15766;
    input n15765;
    input n15764;
    input n15763;
    output \r_Bit_Index[0] ;
    output tx_o;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3497[1] ;
    output n27464;
    output n27476;
    output n4;
    input VCC_net;
    input n15704;
    output n8439;
    input n31237;
    input n15698;
    output tx_enable;
    output \r_SM_Main_2__N_3426[2] ;
    output [2:0]r_SM_Main_adj_11;
    input n26557;
    output \r_Bit_Index[0]_adj_7 ;
    output r_Rx_Data;
    input RX_N_2;
    output n14264;
    output n18753;
    output n14259;
    output n4_adj_8;
    output n15508;
    output n15619;
    output n4_adj_9;
    output n4_adj_10;
    input n15711;
    input n16227;
    input n15707;
    input n26153;
    input n15686;
    input n15685;
    input n15684;
    input n15683;
    input n15681;
    input n15680;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n16, n17, n29802, n25220, n26701, n27063, n15095, n6, 
        n28624, n29801, n16_adj_3883, n17_adj_3884, n29799, n26631, 
        n14751, n6_adj_3885, n14715, n28728, n24228, n26920, n24198, 
        n25156, n29798, n26831, n24287, n24578, n4572, n15432, 
        n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n6_adj_3886, n5, n29727, n7_c, n27124, n25217, n27282, 
        n26872, n30886, n30874, n14, n30664, n29791, n26797, n25249, 
        n24154, n6_adj_3887, n6_adj_3888, n5_adj_3889, n7_adj_3890, 
        n24240, n27199, n14577, n14_adj_3891, n1312, n26690, n15, 
        n14061, n27049, n27165, n26951, n10, n30868, n30856, n14_adj_3892, 
        n30670, n29794, n27019, n16_adj_3893, n26728, n27208, n27056, 
        n26941, n11, n17_adj_3894, n29796, n29795, n27264, n13, 
        n14762, n25128, n6_adj_3895, n26634, n6_adj_3896, n26945, 
        n25120, n15084, n5_adj_3897, n7_adj_3898, n26975, n30862, 
        n30898, n14_adj_3899, n30676, n29797, n16_adj_3900, n27205, 
        n17_adj_3901, n27053, n15275, n26847, n25182, n29793, n29792, 
        n14370, n27190, n24202, n12, n14784, n27013, n26724, n15290, 
        n26790, n27098, n10_adj_3902, n27148, n26907, n28593, n6_adj_3903, 
        n5_adj_3904, n7_adj_3905, n30850, n30712, n14_adj_3906, n30682, 
        n29800, n15110, n26900, n30083, n5_adj_3907, n7_adj_3908, 
        n15114, n27178, n27824, n14730, n14_adj_3909, n9, n12556, 
        n12515, n15162, n30844, n30928, n14_adj_3910, n30688, n29803, 
        n30077, n5_adj_3911, n27202, n15105, n27228, n1427, n24, 
        n7_adj_3912, n14755, n26, n27270, n26772, n25, n30838, 
        n30946, n14_adj_3913, n27060, n27285, n27, n30694, n29806, 
        n6_adj_3914, n27022, n28861, n30070, n5_adj_3915, n27091, 
        n26750, n7_adj_3916, n12513, n26753, n12559, n14313, n27066, 
        n10_adj_3917, n30832, n30814, n14_adj_3918, n30700, n29809, 
        n26706, n25096, n15266, n6_adj_3919, n5_adj_3920, n7_adj_3921, 
        n27069, n30892, n30802, n14_adj_3922, n30706, n29812;
    wire [7:0]n8825;
    
    wire n22434, n26646, n22433, n26794, n22432, n22431, n22430, 
        n22429, n22358, n22359, n2_adj_3923, n22357, n2034, n22428, 
        n17_adj_3924, n15439, n15586, n27016, n14390, n21, n24_adj_3925, 
        n26695, n20, n14911, n14422, n15127, n26628, n25_adj_3926, 
        n33, n22, n2_adj_3927, n22356, n25253, n38, n36, n37, 
        tx_transmit_N_3397, n27101, n35, n25098, n27126, n24627, 
        n24109, n6_adj_3928, n26669, n14868, n27095, n14400, n25143, 
        n26718, n14822, n1265, n24178, n15_adj_3929, n14_adj_3930, 
        n26625, n6_adj_3931, n27246, n6_adj_3932, n27225, n27123, 
        n25207, n26933, n12650, n26636, n6_adj_3933, n28020, n8_c, 
        n26601, n16045, n2656, n3_adj_3934, n3_adj_3935, n3_adj_3936, 
        n3_adj_3937, n3_adj_3938, n3_adj_3939, n3_adj_3940, n3_adj_3941, 
        n3_adj_3942, n3_adj_3943, n3_adj_3944, n3_adj_3945, n3_adj_3946, 
        n3_adj_3947, n3_adj_3948, n3_adj_3949, n3_adj_3950, n16046, 
        n3_adj_3951, n3_adj_3952, n3_adj_3953, n3_adj_3954, n3_adj_3955, 
        n3_adj_3956, n3_adj_3957, n3_adj_3958, n3_adj_3959, n3_adj_3960, 
        n3_adj_3961, n3_adj_3962, n16_adj_3963, n17_adj_3964, n3_adj_3965, 
        n3_adj_3966;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n4571, n4595, n4594, n4593, n4592, n4591, n4590, n4589, 
        n4588;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n4587, n4586, n4585, n4584, n4583, n4582, n4581, n4580;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n4579, n16047, n4578, n4577, n4576, n4575, n4574, n4573, 
        n26592, n15981, n29824, n29823, n16_adj_3967, n17_adj_3968, 
        n29811, n29810, n16_adj_3969, n17_adj_3970, n29808, n29807, 
        n16_adj_3971, n17_adj_3972, n29805, n27037, n6_adj_3973, n14827, 
        n31, n31_adj_3974;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n11503, n16048, Kp_23__N_877;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n28581, Kp_23__N_980, n26676;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n14506, n12_adj_3975, n15190, n27040, n15022, n16049, n14324, 
        n26763, n10_adj_3976, Kp_23__N_814, n12_adj_3977, n14586;
    wire [0:0]n3512;
    wire [2:0]r_SM_Main_2__N_3500;
    
    wire n27430, n16050, n26743, Kp_23__N_974, n14613, n16051, n16052, 
        n26682, \FRAME_MATCHER.rx_data_ready_prev , n161, n26994, n14500, 
        n2_adj_3978, n22355, n8_adj_3979, n16037, n16038, n16039, 
        n25175, n24366, n15263, n2_adj_3980, n22354, n2_adj_3981, 
        n22353, n2_adj_3982, n22383, n2_adj_3983, n22382, n25139, 
        n2_adj_3984, n22381, n27134, n1862, n15693, n16040, n15974, 
        n15975, n15976, n15977, n15978, n15979, n2_adj_3985, n22380, 
        n15980, n2_adj_3986, n22379, Kp_23__N_977, n24238, n28631, 
        n16041, n14637, n12_adj_3987, Kp_23__N_1067, n14_adj_3988, 
        n26735, n26809, n12_adj_3989, n14745, n27139, n29039, n27104, 
        n14806, n26936, n28926, n27043, n10_adj_3990, n27696, n27154, 
        n26987, n15982, n24234, n24273, n28568, n26827, n4_c, 
        n10_adj_3991, n26928, n27163, n2_adj_3992, n22378, n25245, 
        n27132, n11580, n26569, n25811, n19259, n25903, n2_adj_3993, 
        n22377, n16042, n25907, n8_adj_3994, n20_adj_3995, n16043, 
        n8_adj_3996, n49, n37_adj_3997, n28216, n16044, n14553, 
        n15036, n15_adj_3998, n2_adj_3999, n22376, n8_adj_4000, n5_adj_4001, 
        n63_c, n63_adj_4002, n2_adj_4003, n22375, n2_adj_4005, n22374, 
        n14_adj_4006, n18698, n26585, n18667, n11603, n14304, n2_adj_4007, 
        n22373, n11608, n25951, n18692, n26001, n18650, n26015, 
        n26041, n26039, n18690, n26035, n15983, n11991, n26033, 
        n26031, n26029, n26013, n2_adj_4008, n22372, n26011, n26009, 
        n16_adj_4009, n25955, n26027, n26025, n2_adj_4010, n22371, 
        n7_adj_4011, n11544, n13_adj_4012, n4_adj_4013, n26023, n19325, 
        n5_adj_4014, n19260, n27959, n29049, n19295, n16029, n16030, 
        n6_adj_4015, n7_adj_4016, n7_adj_4017, n2_adj_4018, n22370, 
        n7_adj_4019, n15984, n26019, n26021, n26037, n16031, n16032, 
        n26017, n8_adj_4020, n25853, n14120, n14285, n16033, n2_adj_4021, 
        n22369, n14284, n48, n46, n47, n45, n44, n43, n54, 
        n49_adj_4022, n26866, n25179, n26613, n27005, n12843, n27072;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n14_adj_4023;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n25122, n27025, n27168, n15_adj_4024, n26643, Kp_23__N_1194, 
        n26709, n14671, n26657, n12_adj_4025, n27028, n14908, n26666, 
        n27255, n6_adj_4026, n26966, n15199, n16034, n3303, n8_adj_4027, 
        n16035, n16036, n8_adj_4030, n2_adj_4031, n22368, n19293, 
        n14277, Kp_23__N_1079, n27291, n26821, n27151, n12_adj_4032, 
        n27249, n14665, n27107, n26981, n27075, n12_adj_4033, n27217, 
        n15202, n26948, n10_adj_4034, n27288, n27849, n26654, n26972, 
        n26984, n10_adj_4035, n27034, n25169, n14_adj_4036, n25132, 
        Kp_23__N_1382, n27276, n6_adj_4037, n14654, n6_adj_4038, n15058, 
        n26679, n25161, n10_adj_4039, n26880, n26877, n26978, n14526, 
        n14682, n26957, n27294, n16021, n12_adj_4040, n26769, n25187, 
        n12_adj_4041, n27214, n16022, n6_adj_4042, n26664, n27184, 
        n13948, n28209, n27002, n16023, n2_adj_4043, n22367, n16024, 
        n2_adj_4044, n22366, n14_adj_4045, n10_adj_4046, n25171, n25134, 
        n10_adj_4047, n27234, n26903, n14627, n52, n60, n26712, 
        n58, Kp_23__N_1190, n59, n27231, n27187, n26910, n57, 
        n38_adj_4048, n16025, n27279, n54_adj_4049, n27258, n56, 
        n26863, n55, n66, n61, n26860, n14582, n15074, n14455, 
        n27273, n14982, n22_adj_4050, n15302, n16_adj_4051, n24_adj_4052, 
        n20_adj_4053, n27120, n2_adj_4054, n22365, n27171, n6_adj_4055, 
        n12757, n10_adj_4056, n26637, n6_adj_4057, n26766, n16026, 
        n16027, n25136, Kp_23__N_1214, n15317, n10_adj_4058, n16_adj_4059, 
        n15046, n15_adj_4060, n16028, Kp_23__N_804, n14411, n15047, 
        n15_adj_4061, n14515, n14_adj_4062, n15985, n19276, n26482, 
        n27116, n28, n28485, n32, n27046, n26732, n30, n14882, 
        n14327, n31_adj_4063, n25231, n29, n6_adj_4064, n26651, 
        n27145, n5_adj_4065, n25102, n8_adj_4066;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n27667;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n28499, n31308, n14_adj_4067, n14308, n15_adj_4068, n31309, 
        n31310, n10_adj_4069, n28716, n10_adj_4070, n28060, n6_adj_4071, 
        n27883, n10_adj_4072, n28849, n12_adj_4073, n10_adj_4074, 
        n11_adj_4075, n9_adj_4076, n28014, n28808, n28793, n27726, 
        n12_adj_4077, n11_adj_4078, n28789, n13_adj_4079, n30943, 
        n14975, n26890, n10_adj_4080, n30718, n30931;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n26815, n26778, Kp_23__N_904, n6_adj_4081, n27087, n18, 
        n26738, n26775, n26617, n27010, n28235, n30925, n15077, 
        n15244, n30724, n30919, n30730, n30913, Kp_23__N_820, n30736, 
        n30907, n30742, n30901, n26721, n30895, n30889, n30883, 
        n27084, n10_adj_4082, n14550, Kp_23__N_948, n26784, n14332, 
        n30871, n6_adj_4083, n30865, n30859, n30853, n30847, n30841, 
        n30835, n30829, Kp_23__N_872, n8_adj_4084, n16013, n30811, 
        n30799, n27031, n30775, n30173, n30748, n30769, n30763, 
        n30183, n30757, n30751, n30745, n30739, n29804, n30733, 
        n26969, n30727, n26661, n30721, n30715, n16014, n10_adj_4085, 
        n16015, n16016, n16017, n16018, n15986, n15987, n16019, 
        n16020, n30709, n27196;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n30703, n26758, n30697, n8_adj_4086, n16005, n16006, n2_adj_4087, 
        n2_adj_4088, n2_adj_4089, n2_adj_4090, n2_adj_4091, n2_adj_4092, 
        n2_adj_4093, n15474, n2279, n28646, n25148, n10_adj_4094, 
        n26803, n26804, n6_adj_4095, n6_adj_4096, n27243, n17_adj_4097, 
        n26835, n27113, n27240, n27142, n16007, n28402, n28641, 
        n26761, n27629, n15282, n24570, n28404, n26828, n27679, 
        n16008, n30_adj_4098, n26954, n6_adj_4099, n24121, n27160, 
        n10_adj_4100, n25116, n26005, n25855, n25927, n25925, n25909, 
        n25923, n25921, n25919, n25873, n25947, n25937, n25935, 
        n25917, n25915, n25913, n25911, n25797, n25933, n25845, 
        n25843, n25899, n25841, n15577, n26510, n28091, n15988, 
        n26844, n22364, n14292, n4_adj_4101, n16009, n26565, n24254, 
        n26818, n16010, n27452, n13981, n27181, n24115, n5_adj_4102, 
        n6_adj_4103, n16141, n16142, n16143, n16144, n16145, n13_adj_4104, 
        n16011, n28283, n14243, n5_adj_4105, n16146, n16147, n16148, 
        n16012, n6_adj_4106, n1;
    wire [31:0]\FRAME_MATCHER.state_31__N_2608 ;
    
    wire n22363, n14_adj_4107, n8_adj_4108, n15997, n16133, n22362, 
        n16134, n16135, n16136, n26787, n16137, n16138, n16139, 
        n16140, n16125, n14117, n16126, n16127, n16128, n10_adj_4110, 
        n16129, n28313, n30691, n30685, n24_adj_4111, n30679, n22_adj_4112, 
        n30673, n26_adj_4113, n30667, n30661, n15998, n13_adj_4114, 
        n16130, n29021, n30_adj_4115, n15999, n28_adj_4116, n29_adj_4117, 
        n27_adj_4118, n16131, n22361, n16132, n16000, n8_adj_4119, 
        n44_adj_4120, n42, n16117, n16118, n16119, n16120, n16121, 
        n43_adj_4121, n41, n16122, n40, n39, n16123, n16124, n50, 
        n45_adj_4122, n16109, n16110, n16111, n16112, n16113, n16001, 
        n29071, n15_adj_4123, n14293, n14129, n10_adj_4124, n16114, 
        n14_adj_4125, n9_adj_4126, n14296, n16_adj_4127, n17_adj_4128, 
        n14269, n29053, n18_adj_4129, n19, n16_adj_4130, n17_adj_4131, 
        n16115, n16116, n16002, n16108, n16107, n16106, n16105, 
        n16104, n16103, n16102, n16101, n16100, n16099, n16098, 
        n16097, n16096, n16095, n16094, n16093, n16092, n16091, 
        n16090, n16089, n16088, n16087, n16086, n16085, n16084, 
        n16083, n16082, n16081, n16080, n16079, n16078, n16077, 
        n16076, n16075, n16074, n16073, n16072, n16071, n16070, 
        n16069, n16068, n20_adj_4132, n16003, n19_adj_4133, n29075, 
        n16004, n16067, n16066, n16065, n16064, n16063, n16062, 
        n16061, n16060, n16059, n16058, n16057, n16056, n16055, 
        n16054, n16053, n15996, n15995, n15994, n15993, n15992, 
        n15991, n15990, n15989, n26924, n27254, n12_adj_4134, n27237, 
        n26915, n15138, n25094, n10_adj_4135, n24210, n26963, n26869, 
        n26850, n14387, n27778, n27220, n27081, n26715, n14899, 
        n26897, n22_adj_4136, n20_adj_4137, n27261, n24_adj_4138, 
        n14894, n13_adj_4139, n15_adj_4140, n26857, n37_adj_4141, 
        n27136, n28_adj_4142, n36_adj_4143, n42_adj_4144, n40_adj_4145, 
        n41_adj_4146, n26960, n39_adj_4147, n27936, n32_adj_4148, 
        n27078, n30_adj_4149, n31_adj_4150, n29_adj_4151, n14_adj_4152, 
        n15_adj_4153, n10_adj_4154, n18_adj_4155, n26781, n19_adj_4156, 
        n24_adj_4157, n27_adj_4158, n26938, n25204, n26_adj_4159, 
        n30_adj_4160, n25_adj_4161, n10_adj_4162, n14_adj_4163, n27110, 
        n14776, n24200, n22360, n12_adj_4164, n26886, n27532, n6_adj_4165, 
        n7_adj_4166;
    
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24234_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29802));
    defparam i24234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(n25220), .I1(n26701), .I2(\data_out_frame[19] [6]), 
            .I3(n27063), .O(n15095));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n15762));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [0]), 
            .I2(n15095), .I3(n6), .O(n28624));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24236_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29801));
    defparam i24236_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3883));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n15761));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3884));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24239_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29799));
    defparam i24239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_847 (.I0(\data_out_frame[13] [2]), .I1(n26631), 
            .I2(n14751), .I3(n6_adj_3885), .O(n14715));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_847.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n14715), .I1(n28728), .I2(\data_out_frame[15] [3]), 
            .I3(GND_net), .O(n24228));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut (.I0(n24228), .I1(\data_out_frame[19] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n26920));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n15760));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_848 (.I0(n24198), .I1(n26920), .I2(\data_out_frame[17] [3]), 
            .I3(\data_out_frame[17] [4]), .O(n25156));
    defparam i3_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i24241_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29798));
    defparam i24241_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_849 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[24] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26831));
    defparam i1_2_lut_adj_849.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_850 (.I0(\data_out_frame[23] [7]), .I1(n25220), 
            .I2(n24287), .I3(n25156), .O(n24578));
    defparam i3_4_lut_adj_850.LUT_INIT = 16'h9669;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n15432), .D(n4572));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n15759));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i6_3_lut (.I0(\data_out_frame[5] [1]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n6_adj_3886));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut (.I0(n5), .I1(n6_adj_3886), 
            .I2(n29727), .I3(GND_net), .O(n7_c));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_851 (.I0(n27124), .I1(\data_out_frame[23] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25217));
    defparam i1_2_lut_adj_851.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_852 (.I0(\data_out_frame[17] [0]), .I1(n27282), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n26872));
    defparam i2_3_lut_adj_852.LUT_INIT = 16'h9696;
    SB_LUT4 i1495644_i1_3_lut (.I0(n30886), .I1(n30874), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14));
    defparam i1495644_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24279_2_lut (.I0(n30664), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29791));
    defparam i24279_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_853 (.I0(n26872), .I1(\data_out_frame[17] [1]), 
            .I2(n26797), .I3(GND_net), .O(n25249));
    defparam i2_3_lut_adj_853.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n15758));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n15757));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_854 (.I0(n24154), .I1(\data_out_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3887));
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3888));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hb0b3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3889));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut (.I0(n5_adj_3889), 
            .I1(n6_adj_3888), .I2(n29727), .I3(GND_net), .O(n7_adj_3890));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_855 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[12] [2]), .I3(n6_adj_3887), .O(n24240));
    defparam i4_4_lut_adj_855.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[12] [1]), .I1(n27199), .I2(n14577), 
            .I3(GND_net), .O(n14_adj_3891));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[16] [4]), 
            .I2(n1312), .I3(n26690), .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n14061), .I2(n14_adj_3891), .I3(n27049), 
            .O(n27165));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_856 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n26951));
    defparam i2_3_lut_adj_856.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_857 (.I0(n26951), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[7] [6]), .I3(n27165), .O(n10));
    defparam i4_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i1496247_i1_3_lut (.I0(n30868), .I1(n30856), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3892));
    defparam i1496247_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24248_2_lut (.I0(n30670), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29794));
    defparam i24248_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27019));
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3893));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_859 (.I0(n26728), .I1(n27208), .I2(n27056), .I3(n26941), 
            .O(n11));
    defparam i3_4_lut_adj_859.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3894));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24243_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29796));
    defparam i24243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24245_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29795));
    defparam i24245_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[16] [5]), .I1(n27264), .I2(\data_out_frame[12] [1]), 
            .I3(\data_out_frame[14] [3]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n13), .I1(n11), .I2(n14762), .I3(\data_out_frame[14] [4]), 
            .O(n25128));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_860 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3895));
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_861 (.I0(n26634), .I1(n25128), .I2(n27019), .I3(n6_adj_3895), 
            .O(n26797));
    defparam i4_4_lut_adj_861.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3896));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 i3_4_lut_adj_862 (.I0(\data_out_frame[19] [0]), .I1(n26945), 
            .I2(\data_out_frame[18] [6]), .I3(n25120), .O(n15084));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3897));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_adj_3897), 
            .I1(n6_adj_3896), .I2(n29727), .I3(GND_net), .O(n7_adj_3898));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_863 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[11] [0]), .I3(n26975), .O(n28728));
    defparam i3_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i1496850_i1_3_lut (.I0(n30862), .I1(n30898), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3899));
    defparam i1496850_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24244_2_lut (.I0(n30676), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29797));
    defparam i24244_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_864 (.I0(\data_out_frame[5] [4]), .I1(n26690), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n14577));
    defparam i2_3_lut_adj_864.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_865 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n26690));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3900));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_866 (.I0(\data_out_frame[11] [6]), .I1(n26690), 
            .I2(GND_net), .I3(GND_net), .O(n27205));
    defparam i1_2_lut_adj_866.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3901));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_867 (.I0(\data_out_frame[9] [4]), .I1(n27205), 
            .I2(n27053), .I3(\data_out_frame[9] [5]), .O(n15275));
    defparam i3_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_868 (.I0(\data_out_frame[10] [7]), .I1(n26847), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[9] [0]), .O(n25182));
    defparam i3_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i24247_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29793));
    defparam i24247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24249_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29792));
    defparam i24249_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut_adj_869 (.I0(n14370), .I1(n27190), .I2(\data_out_frame[8] [7]), 
            .I3(n24202), .O(n12));
    defparam i5_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_870 (.I0(\data_out_frame[10] [5]), .I1(n12), .I2(n14784), 
            .I3(n27013), .O(n26975));
    defparam i6_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_871 (.I0(\data_out_frame[8] [7]), .I1(n26724), 
            .I2(GND_net), .I3(GND_net), .O(n15290));
    defparam i1_2_lut_adj_871.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_872 (.I0(n26790), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[11] [3]), .I3(n27098), .O(n10_adj_3902));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_873 (.I0(\data_out_frame[11] [2]), .I1(n27148), 
            .I2(n26907), .I3(n15290), .O(n28593));
    defparam i3_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3903));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 i2_3_lut_adj_874 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n27053));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3904));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_3904), 
            .I1(n6_adj_3903), .I2(n29727), .I3(GND_net), .O(n7_adj_3905));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1497453_i1_3_lut (.I0(n30850), .I1(n30712), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3906));
    defparam i1497453_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24240_2_lut (.I0(n30682), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29800));
    defparam i24240_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_875 (.I0(n28593), .I1(n15110), .I2(GND_net), 
            .I3(GND_net), .O(n26900));
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n30083));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3907));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_3907), 
            .I1(byte_transmit_counter[0]), .I2(n29727), .I3(n30083), .O(n7_adj_3908));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1_2_lut_adj_876 (.I0(n15275), .I1(n15114), .I2(GND_net), 
            .I3(GND_net), .O(n27178));
    defparam i1_2_lut_adj_876.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_877 (.I0(n27178), .I1(n27824), .I2(n26900), .I3(n14730), 
            .O(n14_adj_3909));
    defparam i6_4_lut_adj_877.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_878 (.I0(n9), .I1(n14_adj_3909), .I2(n26975), 
            .I3(n25182), .O(n12556));
    defparam i7_4_lut_adj_878.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut (.I0(n12515), .I1(\data_out_frame[7] [0]), .I2(\data_out_frame[6] [5]), 
            .I3(n15162), .O(n27148));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1498056_i1_3_lut (.I0(n30844), .I1(n30928), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3910));
    defparam i1498056_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24235_2_lut (.I0(n30688), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29803));
    defparam i24235_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24225_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30077));   // verilog/coms.v(106[34:55])
    defparam i24225_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut_adj_879 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(n24202), .I3(\data_out_frame[8] [5]), .O(n26847));
    defparam i3_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3911));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_880 (.I0(\data_out_frame[12] [0]), .I1(n27049), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n27202));
    defparam i2_3_lut_adj_880.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut (.I0(n15105), .I1(n26724), .I2(n27228), .I3(n1427), 
            .O(n24));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_3911), 
            .I1(n30077), .I2(n29727), .I3(byte_transmit_counter[0]), .O(n7_adj_3912));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut (.I0(n14755), .I1(\data_out_frame[7] [0]), .I2(\data_out_frame[6] [7]), 
            .I3(\data_out_frame[8] [0]), .O(n26));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n27270), .I1(n26847), .I2(n27148), .I3(n26772), 
            .O(n25));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1498659_i1_3_lut (.I0(n30838), .I1(n30946), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3913));
    defparam i1498659_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(n14577), .I1(n24), .I2(n27060), .I3(n27285), 
            .O(n27));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_881 (.I0(n14370), .I1(n27), .I2(n25), .I3(n26), 
            .O(n26941));
    defparam i1_4_lut_adj_881.LUT_INIT = 16'h9669;
    SB_LUT4 i24232_2_lut (.I0(n30694), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29806));
    defparam i24232_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_882 (.I0(n26941), .I1(n27202), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3914));
    defparam i1_2_lut_adj_882.LUT_INIT = 16'h6666;
    SB_LUT4 i23377_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n29727));   // verilog/coms.v(106[34:55])
    defparam i23377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_883 (.I0(n12556), .I1(\data_out_frame[9] [5]), 
            .I2(n27022), .I3(n6_adj_3914), .O(n28861));
    defparam i4_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i24218_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30070));   // verilog/coms.v(106[34:55])
    defparam i24218_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3915));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_884 (.I0(\data_out_frame[7] [6]), .I1(n27091), 
            .I2(n26750), .I3(n14577), .O(n24154));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n5_adj_3915), 
            .I1(n30070), .I2(n29727), .I3(byte_transmit_counter[0]), .O(n7_adj_3916));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i2_3_lut_adj_885 (.I0(n12513), .I1(n26753), .I2(\data_out_frame[10] [2]), 
            .I3(GND_net), .O(n12559));
    defparam i2_3_lut_adj_885.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_886 (.I0(n24154), .I1(n28861), .I2(n14313), .I3(n27066), 
            .O(n10_adj_3917));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_886.LUT_INIT = 16'h9669;
    SB_LUT4 i1499262_i1_3_lut (.I0(n30832), .I1(n30814), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3918));
    defparam i1499262_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24227_2_lut (.I0(n30700), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29809));
    defparam i24227_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut_adj_887 (.I0(n12559), .I1(n10_adj_3917), .I2(n26706), 
            .I3(GND_net), .O(n25096));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_887.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_888 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n15266));
    defparam i1_2_lut_adj_888.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_889 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14751));
    defparam i1_2_lut_adj_889.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3919));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hb0bc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3920));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_4_lut (.I0(n5_adj_3920), 
            .I1(n6_adj_3919), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n7_adj_3921));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_adj_890 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27208));
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_891 (.I0(\data_out_frame[7] [6]), .I1(n27208), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[14] [7]), 
            .O(n27069));
    defparam i3_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 i1500468_i1_3_lut (.I0(n30892), .I1(n30802), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3922));
    defparam i1500468_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24220_2_lut (.I0(n30706), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29812));
    defparam i24220_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n12515));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n14370));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14755));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 i639_2_lut (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1427));   // verilog/coms.v(71[16:27])
    defparam i639_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n22434), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26646));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n22433), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_896 (.I0(\data_out_frame[6] [4]), .I1(n26646), 
            .I2(\data_out_frame[8] [1]), .I3(\data_out_frame[9] [3]), .O(n27270));
    defparam i3_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_8 (.CI(n22433), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n22434));
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26794));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n22432), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_7 (.CI(n22432), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n22433));
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n22431), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_6 (.CI(n22431), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n22432));
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n22430), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_5 (.CI(n22430), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n22431));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n22429), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_8 (.CI(n22358), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n22359));
    SB_LUT4 add_43_7_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n22357), .O(n2_adj_3923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n22357), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n22358));
    SB_CARRY add_3971_4 (.CI(n22429), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n22430));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n22428), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_3 (.CI(n22428), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n22429));
    SB_LUT4 i4_3_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[10] [1]), 
            .I2(n27264), .I3(GND_net), .O(n17_adj_3924));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n15439), .D(n8825[7]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n15439), .D(n8825[6]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n15439), .D(n8825[5]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n15439), .D(n8825[4]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n15439), .D(n8825[3]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut_adj_898 (.I0(n26794), .I1(n27016), .I2(n27270), .I3(n14390), 
            .O(n21));
    defparam i8_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n15439), .D(n8825[2]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n15439), .D(n8825[1]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_899 (.I0(n21), .I1(n17_adj_3924), .I2(n27091), 
            .I3(n26907), .O(n24_adj_3925));
    defparam i11_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_900 (.I0(n26695), .I1(n24_adj_3925), .I2(n20), 
            .I3(n14370), .O(n27824));
    defparam i12_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n14911));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_902 (.I0(\data_out_frame[6] [2]), .I1(n14911), 
            .I2(\data_out_frame[9] [5]), .I3(n27824), .O(n27228));
    defparam i3_4_lut_adj_902.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_903 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(n15105), .I3(GND_net), .O(n14422));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_904 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n15127));
    defparam i2_3_lut_adj_904.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut (.I0(n26628), .I1(\data_out_frame[8] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3926));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_905 (.I0(n15127), .I1(n14422), .I2(\data_out_frame[6] [0]), 
            .I3(n27228), .O(n33));
    defparam i12_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\data_out_frame[11] [2]), .I1(n27069), 
            .I2(GND_net), .I3(GND_net), .O(n22));
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_6_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n22356), .O(n2_adj_3927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i17_4_lut (.I0(n33), .I1(n25_adj_3926), .I2(\data_out_frame[8] [5]), 
            .I3(n25253), .O(n38));
    defparam i17_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut (.I0(n14751), .I1(\data_out_frame[11] [3]), .I2(\data_out_frame[11] [4]), 
            .I3(\data_out_frame[10] [6]), .O(n36));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n15266), .I1(n25096), .I2(\data_out_frame[7] [7]), 
            .I3(n22), .O(n37));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3397), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3397), 
            .CO(n22428));
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n15756));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14_4_lut (.I0(\data_out_frame[15] [0]), .I1(n26706), .I2(n27101), 
            .I3(\data_out_frame[7] [4]), .O(n35));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37), .I2(n36), .I3(n38), .O(n25098));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_907 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27126));
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_908 (.I0(\data_out_frame[13] [0]), .I1(n24627), 
            .I2(\data_out_frame[15] [2]), .I3(n28728), .O(n24109));
    defparam i3_4_lut_adj_908.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_909 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n26728));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_909.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_910 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3928));
    defparam i1_2_lut_adj_910.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_911 (.I0(\data_out_frame[8] [3]), .I1(n26669), 
            .I2(n26728), .I3(n6_adj_3928), .O(n14868));
    defparam i4_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_912 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14390));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_out_frame[6] [4]), .I1(n26631), 
            .I2(GND_net), .I3(GND_net), .O(n14784));
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_914 (.I0(\data_out_frame[14] [7]), .I1(n25253), 
            .I2(\data_out_frame[13] [0]), .I3(\data_out_frame[15] [1]), 
            .O(n27095));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_914.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_915 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n14400));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_916 (.I0(\data_out_frame[5] [6]), .I1(n26695), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n27056));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_916.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_917 (.I0(n25143), .I1(n27056), .I2(\data_out_frame[8] [1]), 
            .I3(GND_net), .O(n12513));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_917.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\data_out_frame[7] [6]), .I1(n1312), .I2(GND_net), 
            .I3(GND_net), .O(n26718));
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_919 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n26695));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_919.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27016));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_921 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[5] [3]), .O(n26628));
    defparam i3_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_922 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26790));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_922.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26669));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27101));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_925 (.I0(n14822), .I1(n1265), .I2(\data_out_frame[6] [0]), 
            .I3(\data_out_frame[5] [5]), .O(n26724));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_out_frame[5] [7]), .I1(n1265), .I2(GND_net), 
            .I3(GND_net), .O(n26772));
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_927 (.I0(n26628), .I1(n27016), .I2(\data_out_frame[5] [6]), 
            .I3(GND_net), .O(n14822));
    defparam i2_3_lut_adj_927.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_928 (.I0(\data_out_frame[5] [0]), .I1(n26724), 
            .I2(GND_net), .I3(GND_net), .O(n15162));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_929 (.I0(\data_out_frame[5] [0]), .I1(n14822), 
            .I2(n24178), .I3(GND_net), .O(n25143));
    defparam i2_3_lut_adj_929.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_930 (.I0(n27060), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(n26695), .O(n15_adj_3929));
    defparam i6_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_931 (.I0(n15_adj_3929), .I1(n14400), .I2(n14_adj_3930), 
            .I3(n1312), .O(n14061));
    defparam i8_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_932 (.I0(\data_out_frame[10] [1]), .I1(n14061), 
            .I2(GND_net), .I3(GND_net), .O(n26750));
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27013));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_934 (.I0(\data_out_frame[10] [4]), .I1(n27013), 
            .I2(n26625), .I3(\data_out_frame[6] [2]), .O(n14313));
    defparam i3_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_935 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3931));
    defparam i1_2_lut_adj_935.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_936 (.I0(n14762), .I1(n26750), .I2(\data_out_frame[14] [5]), 
            .I3(n6_adj_3931), .O(n27246));
    defparam i4_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_937 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(n6_adj_3932), .I3(\data_out_frame[6] [1]), .O(n26753));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_937.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_938 (.I0(n26753), .I1(\data_out_frame[12] [5]), 
            .I2(n27246), .I3(n14313), .O(n26634));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_939 (.I0(n27095), .I1(n27225), .I2(GND_net), 
            .I3(GND_net), .O(n24198));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27123));
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_941 (.I0(n25207), .I1(\data_out_frame[17] [1]), 
            .I2(n26933), .I3(n27123), .O(n24287));
    defparam i3_4_lut_adj_941.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_942 (.I0(n15084), .I1(n26797), .I2(GND_net), 
            .I3(GND_net), .O(n12650));
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_943 (.I0(\data_out_frame[19] [3]), .I1(n27123), 
            .I2(n26872), .I3(n26636), .O(n27124));
    defparam i3_4_lut_adj_943.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n15755));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_944 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [7]), 
            .I2(n27124), .I3(n6_adj_3933), .O(n28020));
    defparam i4_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i11470_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n16045));
    defparam i11470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_344_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3934));
    defparam select_344_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3935));
    defparam select_344_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3936));
    defparam select_344_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3937));
    defparam select_344_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3938));
    defparam select_344_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3939));
    defparam select_344_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3940));
    defparam select_344_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3941));
    defparam select_344_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3942));
    defparam select_344_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3943));
    defparam select_344_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3944));
    defparam select_344_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3945));
    defparam select_344_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3946));
    defparam select_344_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3947));
    defparam select_344_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3948));
    defparam select_344_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3949));
    defparam select_344_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3950));
    defparam select_344_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11471_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n16046));
    defparam i11471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_344_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3951));
    defparam select_344_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_43_6 (.CI(n22356), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n22357));
    SB_LUT4 select_344_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3952));
    defparam select_344_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3953));
    defparam select_344_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3954));
    defparam select_344_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3955));
    defparam select_344_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3956));
    defparam select_344_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3957));
    defparam select_344_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3958));
    defparam select_344_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3959));
    defparam select_344_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3960));
    defparam select_344_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3961));
    defparam select_344_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3962));
    defparam select_344_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3963));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3964));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_344_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3965));
    defparam select_344_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_344_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3966));
    defparam select_344_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n15754));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n15753));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1068_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4571), .I3(GND_net), .O(n4595));
    defparam mux_1068_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4571), .I3(GND_net), .O(n4594));
    defparam mux_1068_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4571), .I3(GND_net), .O(n4593));
    defparam mux_1068_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4571), .I3(GND_net), .O(n4592));
    defparam mux_1068_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4571), .I3(GND_net), .O(n4591));
    defparam mux_1068_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4571), .I3(GND_net), .O(n4590));
    defparam mux_1068_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4571), .I3(GND_net), .O(n4589));
    defparam mux_1068_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4571), .I3(GND_net), .O(n4588));
    defparam mux_1068_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4571), .I3(GND_net), .O(n4587));
    defparam mux_1068_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4571), .I3(GND_net), .O(n4586));
    defparam mux_1068_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4571), .I3(GND_net), .O(n4585));
    defparam mux_1068_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4571), .I3(GND_net), .O(n4584));
    defparam mux_1068_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4571), .I3(GND_net), .O(n4583));
    defparam mux_1068_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4571), .I3(GND_net), .O(n4582));
    defparam mux_1068_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4571), .I3(GND_net), .O(n4581));
    defparam mux_1068_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4571), .I3(GND_net), .O(n4580));
    defparam mux_1068_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4571), .I3(GND_net), .O(n4579));
    defparam mux_1068_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11472_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n16047));
    defparam i11472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1068_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4571), .I3(GND_net), .O(n4578));
    defparam mux_1068_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4571), .I3(GND_net), .O(n4577));
    defparam mux_1068_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4571), .I3(GND_net), .O(n4576));
    defparam mux_1068_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4571), .I3(GND_net), .O(n4575));
    defparam mux_1068_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4571), .I3(GND_net), .O(n4574));
    defparam mux_1068_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1068_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4571), .I3(GND_net), .O(n4573));
    defparam mux_1068_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11406_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n15981));
    defparam i11406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24204_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29824));
    defparam i24204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24038_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29823));
    defparam i24038_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3967));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3968));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24217_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29811));
    defparam i24217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24221_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29810));
    defparam i24221_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3969));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3970));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24224_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29808));
    defparam i24224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24228_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29807));
    defparam i24228_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3971));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3972));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24230_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29805));
    defparam i24230_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n15752));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_945 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[2] [3]), 
            .I2(n27037), .I3(n6_adj_3973), .O(n14827));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i5071_3_lut (.I0(n31), .I1(n31_adj_3974), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n11503));   // verilog/coms.v(145[4] 299[11])
    defparam i5071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11473_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n16048));
    defparam i11473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_946 (.I0(Kp_23__N_877), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[2] [2]), .O(n28581));   // verilog/coms.v(166[9:87])
    defparam i3_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_947 (.I0(\data_in_frame[2] [0]), .I1(n28581), .I2(\data_in_frame[4] [2]), 
            .I3(\data_in_frame[4] [3]), .O(Kp_23__N_980));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_948 (.I0(\data_in_frame[5] [0]), .I1(n26676), .I2(\data_in_frame[7] [2]), 
            .I3(n14506), .O(n12_adj_3975));
    defparam i5_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_949 (.I0(n15190), .I1(n12_adj_3975), .I2(n27040), 
            .I3(\data_in_frame[5] [1]), .O(n15022));
    defparam i6_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i11474_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n16049));
    defparam i11474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_950 (.I0(\data_in_frame[4] [5]), .I1(n14324), .I2(\data_in_frame[2] [6]), 
            .I3(n26763), .O(n10_adj_3976));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_951 (.I0(Kp_23__N_980), .I1(n14827), .I2(Kp_23__N_814), 
            .I3(\data_in_frame[8] [1]), .O(n12_adj_3977));
    defparam i5_4_lut_adj_951.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_952 (.I0(\data_in_frame[6] [7]), .I1(n10_adj_3976), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n14586));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_adj_952.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n15751));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3500[0]), .C(clk32MHz), 
            .D(n3512[0]), .R(n27430));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11475_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n16050));
    defparam i11475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_953 (.I0(\data_in_frame[8] [4]), .I1(n26743), .I2(Kp_23__N_974), 
            .I3(\data_in_frame[6] [2]), .O(n14613));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i11476_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n16051));
    defparam i11476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11477_3_lut_4_lut (.I0(n8_c), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n16052));
    defparam i11477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_954 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[4] [6]), .I3(GND_net), .O(n26682));
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h9696;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[8] [3]), .I3(n26994), .O(n14500));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_5_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n22355), .O(n2_adj_3978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11462_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n16037));
    defparam i11462_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11463_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n16038));
    defparam i11463_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11464_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n16039));
    defparam i11464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n15750));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n25175), .I1(n24366), .I2(\data_out_frame[15] [5]), 
            .I3(\data_out_frame[17] [7]), .O(n15263));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_43_5 (.CI(n22355), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n22356));
    SB_LUT4 add_43_4_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n22354), .O(n2_adj_3980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n22354), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n22355));
    SB_LUT4 add_43_3_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n22353), .O(n2_adj_3981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_3 (.CI(n22353), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n22354));
    SB_LUT4 add_43_33_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n22383), .O(n2_adj_3982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_2_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_32_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n22382), .O(n2_adj_3983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n22382), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n22383));
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n22353));
    SB_LUT4 i1_2_lut_4_lut_adj_955 (.I0(n25175), .I1(n24366), .I2(\data_out_frame[15] [5]), 
            .I3(n25128), .O(n25139));
    defparam i1_2_lut_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_31_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n22381), .O(n2_adj_3984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_956 (.I0(n25175), .I1(n24366), .I2(\data_out_frame[15] [5]), 
            .I3(n27134), .O(n1862));
    defparam i1_2_lut_4_lut_adj_956.LUT_INIT = 16'h9669;
    SB_LUT4 i11118_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n15693));
    defparam i11118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11465_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n16040));
    defparam i11465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n15749));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11399_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n15974));
    defparam i11399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11400_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n15975));
    defparam i11400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n15748));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11401_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n15976));
    defparam i11401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_31 (.CI(n22381), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n22382));
    SB_LUT4 i11402_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n15977));
    defparam i11402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11403_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n15978));
    defparam i11403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11404_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n15979));
    defparam i11404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_30_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n22380), .O(n2_adj_3985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11405_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n15980));
    defparam i11405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_30 (.CI(n22380), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n22381));
    SB_LUT4 add_43_29_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n22379), .O(n2_adj_3986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n22379), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n22380));
    SB_LUT4 i6_4_lut_adj_957 (.I0(Kp_23__N_977), .I1(n12_adj_3977), .I2(n26994), 
            .I3(n24238), .O(n28631));
    defparam i6_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i11466_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n16041));
    defparam i11466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n15747));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_958 (.I0(n14637), .I1(n12_adj_3987), .I2(Kp_23__N_1067), 
            .I3(\data_in_frame[8] [2]), .O(n14_adj_3988));
    defparam i6_4_lut_adj_958.LUT_INIT = 16'hdffd;
    SB_LUT4 i5_4_lut_adj_959 (.I0(n26735), .I1(n26809), .I2(\data_in_frame[7] [5]), 
            .I3(\data_in_frame[3] [1]), .O(n12_adj_3989));   // verilog/coms.v(73[16:34])
    defparam i5_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i23188_3_lut (.I0(\data_in_frame[8] [0]), .I1(n14745), .I2(n27139), 
            .I3(GND_net), .O(n29039));
    defparam i23188_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i6_4_lut_adj_960 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_3989), 
            .I2(n27104), .I3(\data_in_frame[5] [3]), .O(n14806));   // verilog/coms.v(73[16:34])
    defparam i6_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_961 (.I0(n29039), .I1(n14_adj_3988), .I2(n26936), 
            .I3(n28631), .O(n28926));
    defparam i7_4_lut_adj_961.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_962 (.I0(n26682), .I1(\data_in_frame[6] [6]), .I2(\data_in_frame[4] [4]), 
            .I3(n27043), .O(n10_adj_3990));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_963 (.I0(n15084), .I1(n27696), .I2(\data_out_frame[23] [0]), 
            .I3(n27154), .O(n26987));
    defparam i2_3_lut_4_lut_adj_963.LUT_INIT = 16'h9669;
    SB_LUT4 i11407_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n15982));
    defparam i11407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_964 (.I0(n24234), .I1(n24273), .I2(\data_out_frame[25] [4]), 
            .I3(\data_out_frame[25] [5]), .O(n28568));
    defparam i2_3_lut_4_lut_adj_964.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut (.I0(n24234), .I1(n24273), .I2(n26827), .I3(GND_net), 
            .O(n4_c));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_965 (.I0(n26987), .I1(n10_adj_3991), .I2(\data_out_frame[24] [7]), 
            .I3(n26928), .O(n27163));
    defparam i1_2_lut_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_28_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n22378), .O(n2_adj_3992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_966 (.I0(n26987), .I1(n10_adj_3991), .I2(\data_out_frame[24] [7]), 
            .I3(n25245), .O(n27132));
    defparam i1_2_lut_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [29]), 
            .I3(n26569), .O(n25811));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_967 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [27]), 
            .I3(n26569), .O(n19259));
    defparam i1_2_lut_3_lut_4_lut_adj_967.LUT_INIT = 16'hf020;
    SB_CARRY add_43_28 (.CI(n22378), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n22379));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_968 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [25]), 
            .I3(n26569), .O(n25903));
    defparam i1_2_lut_3_lut_4_lut_adj_968.LUT_INIT = 16'hf020;
    SB_LUT4 add_43_27_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n22377), .O(n2_adj_3993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11467_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n16042));
    defparam i11467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_969 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [24]), 
            .I3(n26569), .O(n25907));
    defparam i1_2_lut_3_lut_4_lut_adj_969.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_970 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [12]), 
            .I3(n26569), .O(n8_adj_3994));
    defparam i1_2_lut_3_lut_4_lut_adj_970.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_971 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [10]), 
            .I3(n26569), .O(n20_adj_3995));
    defparam i1_2_lut_3_lut_4_lut_adj_971.LUT_INIT = 16'hf020;
    SB_LUT4 i11468_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n16043));
    defparam i11468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_972 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [8]), 
            .I3(n26569), .O(n8_adj_3996));
    defparam i1_2_lut_3_lut_4_lut_adj_972.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_4_lut_adj_973 (.I0(n11580), .I1(n14288), .I2(n49), 
            .I3(n37_adj_3997), .O(n28216));
    defparam i2_3_lut_4_lut_adj_973.LUT_INIT = 16'hfff2;
    SB_LUT4 i11469_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n16044));
    defparam i11469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_27 (.CI(n22377), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n22378));
    SB_LUT4 i5_3_lut_adj_974 (.I0(\data_in_frame[0] [4]), .I1(n10_adj_3990), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n14553));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_974.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_975 (.I0(n28926), .I1(n14613), .I2(n15036), .I3(n14586), 
            .O(n15_adj_3998));
    defparam i6_4_lut_adj_975.LUT_INIT = 16'hfffe;
    SB_LUT4 add_43_26_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n22376), .O(n2_adj_3999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_976 (.I0(n11580), .I1(n14288), .I2(\FRAME_MATCHER.state [9]), 
            .I3(n26569), .O(n8_adj_4000));
    defparam i1_2_lut_3_lut_4_lut_adj_976.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_4_lut_adj_977 (.I0(n771), .I1(n9520), .I2(n4609), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n5_adj_4001));   // verilog/coms.v(157[6] 159[9])
    defparam i2_3_lut_4_lut_adj_977.LUT_INIT = 16'h0400;
    SB_CARRY add_43_26 (.CI(n22376), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n22377));
    SB_LUT4 i2_3_lut_4_lut_adj_978 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(n24178), .I3(n26718), .O(n27060));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_979 (.I0(n771), .I1(n9520), .I2(n14253), 
            .I3(GND_net), .O(n37_adj_3997));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_3_lut_adj_979.LUT_INIT = 16'h0404;
    SB_LUT4 i14296_2_lut_3_lut (.I0(n63_c), .I1(n63_adj_4002), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n123));
    defparam i14296_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_43_25_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n22375), .O(n2_adj_4003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_980 (.I0(n63_c), .I1(n63_adj_4002), .I2(n63), 
            .I3(GND_net), .O(n9520));
    defparam i1_2_lut_3_lut_adj_980.LUT_INIT = 16'h8080;
    SB_CARRY add_43_25 (.CI(n22375), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n22376));
    SB_LUT4 add_43_24_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n22374), .O(n2_adj_4005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_981 (.I0(n15_adj_3998), .I1(n15022), .I2(n14_adj_4006), 
            .I3(n14500), .O(n31_adj_3974));
    defparam i8_4_lut_adj_981.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_982 (.I0(n18698), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n26585));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_982.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_3_lut_adj_983 (.I0(tx_transmit_N_3397), .I1(n18667), 
            .I2(n9520), .I3(GND_net), .O(n11603));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_983.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_24 (.CI(n22374), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n22375));
    SB_LUT4 i1_2_lut_3_lut_adj_984 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n27049));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_984.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_985 (.I0(tx_transmit_N_3397), .I1(n18667), 
            .I2(n14304), .I3(GND_net), .O(n26561));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_985.LUT_INIT = 16'h0e0e;
    SB_LUT4 add_43_23_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n22373), .O(n2_adj_4007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n22373), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n22374));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_986 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [31]), 
            .I3(n49), .O(n25951));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_986.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_987 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [29]), 
            .I3(n49), .O(n18692));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_987.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_988 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [28]), 
            .I3(n49), .O(n26001));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_988.LUT_INIT = 16'hf020;
    SB_LUT4 i14087_2_lut_3_lut_4_lut (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [27]), 
            .I3(n49), .O(n18650));   // verilog/coms.v(254[5:25])
    defparam i14087_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_989 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [26]), 
            .I3(n49), .O(n26015));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_989.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_990 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [25]), 
            .I3(n49), .O(n26041));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_990.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_991 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [24]), 
            .I3(n49), .O(n26039));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_991.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_4_lut_adj_992 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[5] [1]), .I3(n27022), .O(n15114));
    defparam i2_3_lut_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i14126_2_lut_3_lut_4_lut (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [23]), 
            .I3(n49), .O(n18690));   // verilog/coms.v(254[5:25])
    defparam i14126_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_993 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [22]), 
            .I3(n49), .O(n26035));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_993.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_4_lut_adj_994 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [0]), .O(n1312));
    defparam i2_3_lut_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i11408_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n15983));
    defparam i11408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_995 (.I0(\FRAME_MATCHER.state [1]), .I1(n31_adj_3974), 
            .I2(n11991), .I3(GND_net), .O(n4571));
    defparam i2_3_lut_adj_995.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_996 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [21]), 
            .I3(n49), .O(n26033));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_996.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_997 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [20]), 
            .I3(n49), .O(n26031));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_997.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_998 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [19]), 
            .I3(n49), .O(n26029));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_998.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_999 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [18]), 
            .I3(n49), .O(n26013));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_999.LUT_INIT = 16'hf020;
    SB_LUT4 add_43_22_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n22372), .O(n2_adj_4008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1000 (.I0(\data_out_frame[12] [5]), .I1(n14868), 
            .I2(n26753), .I3(GND_net), .O(n27225));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1000.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1001 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [17]), 
            .I3(n49), .O(n26011));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1001.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1002 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [16]), 
            .I3(n49), .O(n26009));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1002.LUT_INIT = 16'hf020;
    SB_CARRY add_43_22 (.CI(n22372), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n22373));
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[12] [5]), .I1(n14868), .I2(n25096), 
            .I3(GND_net), .O(n16_adj_4009));   // verilog/coms.v(75[16:43])
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1003 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [15]), 
            .I3(n49), .O(n25955));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1003.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_4_lut_adj_1004 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[12] [3]), .I3(\data_out_frame[12] [4]), 
            .O(n27066));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1005 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [14]), 
            .I3(n49), .O(n26027));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1005.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1006 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [13]), 
            .I3(n49), .O(n26025));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1006.LUT_INIT = 16'hf020;
    SB_LUT4 add_43_21_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n22371), .O(n2_adj_4010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1007 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [12]), 
            .I3(n49), .O(n7_adj_4011));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1007.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_4_lut_adj_1008 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(n14784), .I3(n14313), .O(n24627));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n11544));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1010 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [1]), .O(n13_adj_4012));
    defparam i5_4_lut_adj_1010.LUT_INIT = 16'hfeff;
    SB_LUT4 i23196_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n4_adj_4013), 
            .I2(GND_net), .I3(GND_net), .O(n4677));
    defparam i23196_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i21581_4_lut (.I0(n14254), .I1(\FRAME_MATCHER.state[3] ), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n11544), .O(n27430));
    defparam i21581_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1011 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [11]), 
            .I3(n49), .O(n26023));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1011.LUT_INIT = 16'hf020;
    SB_LUT4 i3_4_lut_adj_1012 (.I0(n19325), .I1(n5_adj_4014), .I2(n18667), 
            .I3(n19260), .O(n27959));
    defparam i3_4_lut_adj_1012.LUT_INIT = 16'hfeff;
    SB_LUT4 mux_789_i1_3_lut (.I0(n27959), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n4677), .I3(GND_net), .O(n3512[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_789_i1_3_lut.LUT_INIT = 16'h5c5c;
    SB_LUT4 i7_4_lut_adj_1013 (.I0(n13_adj_4012), .I1(n29049), .I2(\data_in_frame[0] [0]), 
            .I3(\data_in_frame[0] [2]), .O(n11991));
    defparam i7_4_lut_adj_1013.LUT_INIT = 16'hefff;
    SB_LUT4 i11454_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n16029));
    defparam i11454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11455_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n16030));
    defparam i11455_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(n11991), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4015));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1015 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [10]), 
            .I3(n49), .O(n7_adj_4016));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1015.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1016 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [9]), 
            .I3(n49), .O(n7_adj_4017));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1016.LUT_INIT = 16'hf020;
    SB_CARRY add_43_21 (.CI(n22371), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n22372));
    SB_LUT4 add_43_20_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n22370), .O(n2_adj_4018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1017 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [8]), 
            .I3(n49), .O(n7_adj_4019));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1017.LUT_INIT = 16'hf020;
    SB_LUT4 i11409_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n15984));
    defparam i11409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1018 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [5]), 
            .I3(n49), .O(n26019));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1018.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1019 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [6]), 
            .I3(n49), .O(n26021));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1019.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1020 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [7]), 
            .I3(n49), .O(n26037));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1020.LUT_INIT = 16'hf020;
    SB_LUT4 i11456_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n16031));
    defparam i11456_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11457_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n16032));
    defparam i11457_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1021 (.I0(n11608), .I1(n14291), .I2(\FRAME_MATCHER.state [4]), 
            .I3(n49), .O(n26017));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1021.LUT_INIT = 16'hf020;
    SB_CARRY add_43_20 (.CI(n22370), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n22371));
    SB_LUT4 i1_3_lut_4_lut (.I0(n11608), .I1(n14291), .I2(n8_adj_4020), 
            .I3(\FRAME_MATCHER.state[3] ), .O(n25853));   // verilog/coms.v(254[5:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1083_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4609));   // verilog/coms.v(145[4] 299[11])
    defparam i1083_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\FRAME_MATCHER.state[3] ), .I1(n14254), 
            .I2(GND_net), .I3(GND_net), .O(n14120));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1023 (.I0(n14120), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n14285));   // verilog/coms.v(146[5:9])
    defparam i1_2_lut_4_lut_adj_1023.LUT_INIT = 16'hfffb;
    SB_LUT4 i11458_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n16033));
    defparam i11458_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_43_19_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n22369), .O(n2_adj_4021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1024 (.I0(n14120), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n14284));   // verilog/coms.v(146[5:9])
    defparam i1_2_lut_4_lut_adj_1024.LUT_INIT = 16'hfbff;
    SB_LUT4 select_344_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2656), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_344_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23198_2_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n29049));
    defparam i23198_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1025 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [4]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n48));
    defparam i20_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(\FRAME_MATCHER.state [22]), .I3(\FRAME_MATCHER.state [25]), 
            .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.state [26]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(\FRAME_MATCHER.state [19]), .I3(\FRAME_MATCHER.state [16]), 
            .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1026 (.I0(\FRAME_MATCHER.state [17]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [15]), .I3(\FRAME_MATCHER.state [11]), 
            .O(n45));
    defparam i17_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1027 (.I0(\FRAME_MATCHER.state [9]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(\FRAME_MATCHER.state [31]), 
            .O(n44));
    defparam i16_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1028 (.I0(\FRAME_MATCHER.state [8]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [13]), .I3(\FRAME_MATCHER.state [14]), 
            .O(n43));
    defparam i15_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [5]), 
            .I2(\FRAME_MATCHER.state [24]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n49_adj_4022));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4022), .I1(n54), .I2(n43), .I3(n44), 
            .O(n14254));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_in_frame[12] [3]), .I1(n26866), 
            .I2(GND_net), .I3(GND_net), .O(n25179));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(\data_in_frame[19] [5]), .I1(n26613), 
            .I2(\data_in_frame[19] [6]), .I3(GND_net), .O(n27005));
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_in_frame[18] [1]), .I1(n12843), 
            .I2(GND_net), .I3(GND_net), .O(n27072));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1032 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n14_adj_4023));   // verilog/coms.v(72[16:41])
    defparam i5_3_lut_adj_1032.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1033 (.I0(\data_in_frame[14] [0]), .I1(n25122), 
            .I2(n27025), .I3(n27168), .O(n15_adj_4024));   // verilog/coms.v(72[16:41])
    defparam i6_4_lut_adj_1033.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1034 (.I0(n15_adj_4024), .I1(n26643), .I2(n14_adj_4023), 
            .I3(Kp_23__N_1194), .O(n26709));   // verilog/coms.v(72[16:41])
    defparam i8_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1035 (.I0(n14671), .I1(n26657), .I2(\data_in_frame[12] [5]), 
            .I3(n15036), .O(n12_adj_4025));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1036 (.I0(\data_in_frame[13] [1]), .I1(n12_adj_4025), 
            .I2(n27028), .I3(\data_in_frame[10] [7]), .O(n14908));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(n26666), .I1(n27255), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4026));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1038 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[14] [7]), 
            .I2(n26966), .I3(n6_adj_4026), .O(n15199));
    defparam i4_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i11459_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n16034));
    defparam i11459_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n15746));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1039 (.I0(n63), .I1(n3303), .I2(n123), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2672[1] ));
    defparam i2_3_lut_adj_1039.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_94_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4027));
    defparam equal_94_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i4104_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n8595));   // verilog/coms.v(157[6] 159[9])
    defparam i4104_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14285_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4002), 
            .I2(n63_c), .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i14285_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i11460_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n16035));
    defparam i11460_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_43_19 (.CI(n22369), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n22370));
    SB_LUT4 i14147_3_lut (.I0(n122), .I1(n3303), .I2(n63), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2672[2] ));   // verilog/coms.v(227[6] 229[9])
    defparam i14147_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 select_372_Select_2_i7_4_lut (.I0(n122), .I1(n14291), .I2(n4452), 
            .I3(n63), .O(n7));
    defparam select_372_Select_2_i7_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 select_372_Select_2_i8_3_lut (.I0(n122), .I1(n2649), .I2(n63), 
            .I3(GND_net), .O(n8));
    defparam select_372_Select_2_i8_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i14728_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n19295));
    defparam i14728_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i11461_3_lut_4_lut (.I0(n19295), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n16036));
    defparam i11461_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1570_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4030));
    defparam i1570_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 add_43_18_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n22368), .O(n2_adj_4031)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 equal_91_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_c));   // verilog/coms.v(154[7:23])
    defparam equal_91_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_92_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3979));   // verilog/coms.v(154[7:23])
    defparam equal_92_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1040 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n5_adj_4014));
    defparam i2_3_lut_adj_1040.LUT_INIT = 16'hfefe;
    SB_LUT4 i14726_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n19293));
    defparam i14726_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n19293), .I3(byte_transmit_counter[2]), .O(n19325));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i24768_2_lut (.I0(n19325), .I1(n5_adj_4014), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3397));
    defparam i24768_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_3_lut_adj_1041 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n14506));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1041.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(\FRAME_MATCHER.state [2]), .I1(n14277), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n4_adj_4013), .O(n14279));
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'hfeee;
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n15745));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1043 (.I0(Kp_23__N_1079), .I1(n27291), .I2(\data_in_frame[12] [6]), 
            .I3(\data_in_frame[8] [6]), .O(n26657));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1044 (.I0(n26821), .I1(n27151), .I2(\data_in_frame[13] [0]), 
            .I3(n26657), .O(n12_adj_4032));
    defparam i5_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1045 (.I0(\data_in_frame[17] [4]), .I1(n12_adj_4032), 
            .I2(n27249), .I3(n14665), .O(n27107));
    defparam i6_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1046 (.I0(n26981), .I1(n27075), .I2(\data_in_frame[10] [6]), 
            .I3(n26966), .O(n12_adj_4033));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1047 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_4033), 
            .I2(n27217), .I3(\data_in_frame[14] [6]), .O(n15202));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1048 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n27028));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1049 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n27291));
    defparam i2_3_lut_adj_1049.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1050 (.I0(n14637), .I1(\data_in_frame[13] [7]), 
            .I2(n26948), .I3(\data_in_frame[11] [6]), .O(n10_adj_4034));
    defparam i4_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27288));
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1052 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [3]), 
            .I2(n27849), .I3(GND_net), .O(n26654));
    defparam i2_3_lut_adj_1052.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26948));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1054 (.I0(\data_in_frame[9] [3]), .I1(n27025), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[11] [3]), .O(n26972));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27217));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(n26984), .I1(\data_in_frame[16] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4035));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1056 (.I0(n27034), .I1(n25169), .I2(n26972), 
            .I3(\data_in_frame[15] [7]), .O(n14_adj_4036));
    defparam i6_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1057 (.I0(\data_in_frame[16] [2]), .I1(n14_adj_4036), 
            .I2(n10_adj_4035), .I3(n26948), .O(n25132));
    defparam i7_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_17__7__I_0_3899_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1382));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_17__7__I_0_3899_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(\data_in_frame[12] [4]), .I1(n27276), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4037));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h6666;
    SB_CARRY add_43_18 (.CI(n22368), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n22369));
    SB_LUT4 i4_4_lut_adj_1059 (.I0(n14806), .I1(\data_in_frame[14] [5]), 
            .I2(\data_in_frame[12] [3]), .I3(n6_adj_4037), .O(n26666));
    defparam i4_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1060 (.I0(\data_in_frame[10] [3]), .I1(n14654), 
            .I2(\data_in_frame[6] [0]), .I3(n6_adj_4038), .O(n14671));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1061 (.I0(\data_in_frame[14] [4]), .I1(n15058), 
            .I2(\data_in_frame[12] [2]), .I3(n26679), .O(n26866));
    defparam i3_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1062 (.I0(\data_in_frame[18] [7]), .I1(n26666), 
            .I2(n25161), .I3(\data_in_frame[16] [5]), .O(n10_adj_4039));
    defparam i4_4_lut_adj_1062.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1063 (.I0(n14671), .I1(n10_adj_4039), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n26880));
    defparam i5_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(Kp_23__N_1194), .I1(\data_in_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26877));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1065 (.I0(n14586), .I1(n26978), .I2(n14526), 
            .I3(GND_net), .O(n14682));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1065.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26957));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1067 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[13] [2]), .I3(GND_net), .O(n27294));
    defparam i2_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i11446_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n16021));
    defparam i11446_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1068 (.I0(n14613), .I1(n26643), .I2(\data_in_frame[11] [0]), 
            .I3(n14553), .O(n12_adj_4040));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1069 (.I0(\data_in_frame[10] [6]), .I1(n12_adj_4040), 
            .I2(\data_in_frame[10] [7]), .I3(n27294), .O(n26769));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1070 (.I0(n26769), .I1(\data_in_frame[17] [5]), 
            .I2(n25187), .I3(GND_net), .O(n26613));
    defparam i2_3_lut_adj_1070.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27168));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1072 (.I0(n14526), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[15] [6]), .I3(n26877), .O(n12_adj_4041));   // verilog/coms.v(73[16:42])
    defparam i5_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1073 (.I0(\data_in_frame[9] [0]), .I1(n12_adj_4041), 
            .I2(\data_in_frame[13] [4]), .I3(\data_in_frame[18] [0]), .O(n27214));   // verilog/coms.v(73[16:42])
    defparam i6_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_LUT4 i11447_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n16022));
    defparam i11447_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[11] [5]), .I1(n14526), 
            .I2(GND_net), .I3(GND_net), .O(n27034));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[9] [4]), 
            .I2(n6_adj_4042), .I3(n26664), .O(n27184));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(n13948), .I1(n27214), .I2(n28209), .I3(GND_net), 
            .O(n27002));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i11448_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n16023));
    defparam i11448_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_17_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n22367), .O(n2_adj_4043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n22367), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n22368));
    SB_LUT4 i11449_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n16024));
    defparam i11449_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_16_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n22366), .O(n2_adj_4044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1076 (.I0(n27184), .I1(\data_in_frame[13] [3]), 
            .I2(n26957), .I3(n14682), .O(n14_adj_4045));
    defparam i6_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1077 (.I0(\data_in_frame[17] [7]), .I1(n14_adj_4045), 
            .I2(n10_adj_4046), .I3(n25171), .O(n12843));
    defparam i7_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i14104_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3500[0]), .I2(GND_net), 
            .I3(GND_net), .O(n18667));
    defparam i14104_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(n27002), .I1(\data_in_frame[16] [0]), 
            .I2(n25134), .I3(n27184), .O(n10_adj_4047));
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1079 (.I0(\data_in_frame[19] [7]), .I1(n26613), 
            .I2(n10_adj_4047), .I3(\data_in_frame[15] [7]), .O(n27234));
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_1080 (.I0(\data_in_frame[17] [4]), .I1(n27255), 
            .I2(n26903), .I3(n14627), .O(n52));
    defparam i18_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i26_3_lut (.I0(\data_in_frame[18] [1]), .I1(n52), .I2(\data_in_frame[18] [6]), 
            .I3(GND_net), .O(n60));
    defparam i26_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i24_4_lut (.I0(n26880), .I1(n26712), .I2(n26866), .I3(n14806), 
            .O(n58));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[14] [1]), 
            .I2(Kp_23__N_1190), .I3(\data_in_frame[18] [5]), .O(n59));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n27231), .I1(n26978), .I2(n27187), .I3(n26910), 
            .O(n57));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut_adj_1081 (.I0(\data_in_frame[18] [3]), .I1(n15036), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n38_adj_4048));
    defparam i4_3_lut_adj_1081.LUT_INIT = 16'h9696;
    SB_LUT4 i11450_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n16025));
    defparam i11450_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n15744));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i20_4_lut_adj_1082 (.I0(n25132), .I1(n27217), .I2(n27279), 
            .I3(n26957), .O(n54_adj_4049));
    defparam i20_4_lut_adj_1082.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut (.I0(\data_in_frame[18] [2]), .I1(n27288), .I2(n27294), 
            .I3(n27258), .O(n56));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1083 (.I0(n26877), .I1(n26863), .I2(n26654), 
            .I3(\data_in_frame[14] [2]), .O(n55));
    defparam i21_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i32_4_lut (.I0(n57), .I1(n59), .I2(n58), .I3(n60), .O(n66));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut_adj_1084 (.I0(n27291), .I1(n54_adj_4049), .I2(n38_adj_4048), 
            .I3(n27028), .O(n61));
    defparam i27_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n61), .I1(n66), .I2(n55), .I3(n56), .O(n25134));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1085 (.I0(n25134), .I1(n27234), .I2(n12843), 
            .I3(GND_net), .O(n26860));
    defparam i2_3_lut_adj_1085.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1086 (.I0(n14682), .I1(n26654), .I2(n25122), 
            .I3(\data_in_frame[14] [0]), .O(n13948));
    defparam i3_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_CARRY add_43_16 (.CI(n22366), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n22367));
    SB_LUT4 i3_4_lut_adj_1087 (.I0(n14582), .I1(n15074), .I2(\data_in_frame[10] [1]), 
            .I3(\data_in_frame[9] [7]), .O(n27276));
    defparam i3_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1088 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27258));
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1089 (.I0(n14455), .I1(n27037), .I2(n27273), 
            .I3(n14982), .O(n22_adj_4050));
    defparam i9_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1090 (.I0(n15302), .I1(n22_adj_4050), .I2(n16_adj_4051), 
            .I3(\data_in_frame[13] [7]), .O(n24_adj_4052));
    defparam i11_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1091 (.I0(\data_in_frame[8] [0]), .I1(n24_adj_4052), 
            .I2(n20_adj_4053), .I3(n24238), .O(n26984));
    defparam i12_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1092 (.I0(\data_in_frame[12] [2]), .I1(n27276), 
            .I2(n27231), .I3(n27120), .O(n25161));
    defparam i3_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_15_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n22365), .O(n2_adj_4054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11011_2_lut (.I0(n15439), .I1(n14304), .I2(GND_net), .I3(GND_net), 
            .O(n15586));   // verilog/coms.v(127[12] 300[6])
    defparam i11011_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n15743));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n15742));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\data_in_frame[10] [7]), .I1(n27249), 
            .I2(GND_net), .I3(GND_net), .O(n26910));
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(n14745), .I1(n14586), .I2(GND_net), 
            .I3(GND_net), .O(n25169));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26821));
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(n14500), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27171));
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14627));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n15439), .D(n8825[0]), .R(n15586));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_in_frame[12] [7]), .I1(n15036), 
            .I2(GND_net), .I3(GND_net), .O(n26981));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1099 (.I0(n25169), .I1(n27151), .I2(n26910), 
            .I3(n15036), .O(n25171));
    defparam i3_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1100 (.I0(n25171), .I1(n26981), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4055));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1101 (.I0(n14627), .I1(n27171), .I2(n26821), 
            .I3(n6_adj_4055), .O(n25187));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1102 (.I0(\data_in_frame[7] [6]), .I1(n12757), 
            .I2(\data_in_frame[10] [2]), .I3(n26936), .O(n10_adj_4056));
    defparam i4_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(n14745), .I1(n15022), .I2(GND_net), 
            .I3(GND_net), .O(n26664));
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1104 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [4]), 
            .I2(n26637), .I3(n6_adj_4057), .O(n26863));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1105 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26766));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1105.LUT_INIT = 16'h6666;
    SB_LUT4 i11451_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n16026));
    defparam i11451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11452_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n16027));
    defparam i11452_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_15 (.CI(n22365), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n22366));
    SB_LUT4 i1_2_lut_adj_1106 (.I0(n14582), .I1(n27139), .I2(GND_net), 
            .I3(GND_net), .O(n25136));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n14553), .I1(n14586), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1214));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1108 (.I0(Kp_23__N_1214), .I1(n15317), .I2(n25136), 
            .I3(n10_adj_4058), .O(n16_adj_4059));
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1109 (.I0(n26863), .I1(n14806), .I2(Kp_23__N_1194), 
            .I3(n15046), .O(n15_adj_4060));
    defparam i6_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1110 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[12] [0]), 
            .I2(n15_adj_4060), .I3(n16_adj_4059), .O(n27279));
    defparam i2_4_lut_adj_1110.LUT_INIT = 16'h9669;
    SB_LUT4 i24719_4_lut (.I0(n27362), .I1(\FRAME_MATCHER.state [2]), .I2(n11503), 
            .I3(n6_adj_4015), .O(n15432));
    defparam i24719_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i11453_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n16028));
    defparam i11453_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 data_in_frame_8__7__I_0_3890_2_lut (.I0(\data_in_frame[8] [7]), 
            .I1(\data_in_frame[8] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_804));   // verilog/coms.v(71[16:27])
    defparam data_in_frame_8__7__I_0_3890_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14411));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1112 (.I0(Kp_23__N_804), .I1(n15047), .I2(n26682), 
            .I3(n27279), .O(n15_adj_4061));
    defparam i6_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1113 (.I0(n15_adj_4061), .I1(n14515), .I2(n14_adj_4062), 
            .I3(\data_in_frame[8] [3]), .O(n27273));
    defparam i8_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i11410_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n15985));
    defparam i11410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14710_1_lut (.I0(n19276), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2034));
    defparam i14710_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1114 (.I0(n14285), .I1(n26482), .I2(n31), .I3(GND_net), 
            .O(n4772));
    defparam i2_3_lut_adj_1114.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_4_lut_adj_1115 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[9] [0]), .O(n6_adj_3885));
    defparam i1_2_lut_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1190));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1116 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n26637));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1116.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27116));
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n14654));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1119 (.I0(n14654), .I1(n27116), .I2(n26637), 
            .I3(\data_in_frame[4] [3]), .O(n28));
    defparam i10_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(n14806), .I1(\data_in_frame[11] [7]), 
            .I2(n26679), .I3(n27120), .O(n28485));
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(\data_in_frame[0] [2]), .I1(n28), .I2(\data_in_frame[7] [1]), 
            .I3(GND_net), .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1121 (.I0(n28485), .I1(n27046), .I2(n27273), 
            .I3(n26732), .O(n30));
    defparam i12_4_lut_adj_1121.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[4] [7]), 
            .I2(n14882), .I3(n14327), .O(n31_adj_4063));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1122 (.I0(\data_in_frame[14] [2]), .I1(n25231), 
            .I2(n26766), .I3(\data_in_frame[5] [0]), .O(n29));
    defparam i11_4_lut_adj_1122.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_1123 (.I0(n29), .I1(n31_adj_4063), .I2(n30), 
            .I3(n32), .O(n27849));
    defparam i17_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1124 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26903));
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_in_frame[12] [4]), .I1(n15058), 
            .I2(GND_net), .I3(GND_net), .O(n27075));
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1126 (.I0(n14665), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n26712));
    defparam i2_3_lut_adj_1126.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4064));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1128 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[16] [4]), 
            .I2(n27849), .I3(n6_adj_4064), .O(n26651));   // verilog/coms.v(72[16:41])
    defparam i4_4_lut_adj_1128.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1129 (.I0(n26712), .I1(n27075), .I2(n26903), 
            .I3(\data_in_frame[16] [6]), .O(n27145));
    defparam i3_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1130 (.I0(n25161), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[16] [3]), .I3(n26984), .O(n28209));
    defparam i3_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1131 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [3]), .I3(\data_in_frame[19] [2]), .O(n5_adj_4065));
    defparam i1_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(n5_adj_4065), .I1(n27234), .I2(n27005), .I3(GND_net), 
            .O(n25102));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1132 (.I0(n25102), .I1(\data_in_frame[19] [0]), 
            .I2(n28209), .I3(GND_net), .O(n8_adj_4066));
    defparam i3_3_lut_adj_1132.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_1133 (.I0(n13948), .I1(n26860), .I2(n28209), 
            .I3(\data_in_frame[20] [1]), .O(n27667));
    defparam i2_4_lut_adj_1133.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1134 (.I0(\data_in_frame[19] [1]), .I1(n27145), 
            .I2(n26651), .I3(\data_in_frame[21] [2]), .O(n28499));
    defparam i3_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_rep_11_2_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n31308));
    defparam i1_rep_11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1135 (.I0(\data_in_frame[20] [0]), .I1(n25187), 
            .I2(\data_in_frame[19] [6]), .I3(GND_net), .O(n14_adj_4067));
    defparam i5_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1136 (.I0(n14308), .I1(n27107), .I2(n25169), 
            .I3(n27002), .O(n15_adj_4068));
    defparam i6_4_lut_adj_1136.LUT_INIT = 16'h9669;
    SB_LUT4 i1_rep_12_2_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n31309));
    defparam i1_rep_12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_rep_13_2_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n31310));
    defparam i1_rep_13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1137 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[19] [3]), 
            .I2(n15202), .I3(n27145), .O(n10_adj_4069));
    defparam i4_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1138 (.I0(\data_in_frame[21] [5]), .I1(n31310), 
            .I2(n15199), .I3(n14908), .O(n28716));
    defparam i3_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1139 (.I0(n25169), .I1(n15202), .I2(\data_in_frame[21] [6]), 
            .I3(n27107), .O(n10_adj_4070));
    defparam i4_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1140 (.I0(\data_in_frame[19] [4]), .I1(n10_adj_4070), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n28060));
    defparam i5_3_lut_adj_1140.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1141 (.I0(n13948), .I1(\data_in_frame[18] [4]), 
            .I2(n28209), .I3(GND_net), .O(n6_adj_4071));
    defparam i2_3_lut_adj_1141.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1142 (.I0(\data_in_frame[18] [3]), .I1(n26709), 
            .I2(\data_in_frame[20] [4]), .I3(n25132), .O(n27883));
    defparam i3_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1143 (.I0(n27072), .I1(n14308), .I2(Kp_23__N_1382), 
            .I3(n27214), .O(n10_adj_4072));
    defparam i4_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(n26709), .I1(n27072), .I2(\data_in_frame[20] [3]), 
            .I3(GND_net), .O(n28849));
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1145 (.I0(n27667), .I1(\data_in_frame[18] [5]), 
            .I2(n8_adj_4066), .I3(\data_in_frame[20] [7]), .O(n12_adj_4073));
    defparam i4_4_lut_adj_1145.LUT_INIT = 16'hbeeb;
    SB_LUT4 i2_4_lut_adj_1146 (.I0(n28499), .I1(\data_in_frame[21] [7]), 
            .I2(n27005), .I3(n14908), .O(n10_adj_4074));
    defparam i2_4_lut_adj_1146.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut_4_lut_adj_1147 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[6] [4]), .O(n24202));
    defparam i1_2_lut_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1068_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4571), .I3(GND_net), .O(n4572));
    defparam mux_1068_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1148 (.I0(n27883), .I1(\data_in_frame[18] [5]), 
            .I2(n6_adj_4071), .I3(\data_in_frame[20] [6]), .O(n11_adj_4075));
    defparam i3_4_lut_adj_1148.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_4_lut_adj_1149 (.I0(n26769), .I1(n28849), .I2(n10_adj_4072), 
            .I3(\data_in_frame[20] [2]), .O(n9_adj_4076));
    defparam i1_4_lut_adj_1149.LUT_INIT = 16'hdeed;
    SB_LUT4 i3_4_lut_adj_1150 (.I0(\data_in_frame[20] [5]), .I1(n31308), 
            .I2(n13948), .I3(n25132), .O(n28014));
    defparam i3_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1151 (.I0(n15_adj_4068), .I1(n27187), .I2(n14_adj_4067), 
            .I3(n26860), .O(n28808));
    defparam i8_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1152 (.I0(n15199), .I1(\data_in_frame[21] [3]), 
            .I2(n26880), .I3(n31309), .O(n28793));
    defparam i3_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1153 (.I0(\data_in_frame[21] [0]), .I1(n26651), 
            .I2(n25179), .I3(n25102), .O(n27726));
    defparam i3_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1154 (.I0(n25179), .I1(n28716), .I2(n10_adj_4069), 
            .I3(\data_in_frame[21] [4]), .O(n12_adj_4077));
    defparam i4_4_lut_adj_1154.LUT_INIT = 16'hdeed;
    SB_LUT4 i3_4_lut_adj_1155 (.I0(n25102), .I1(n28060), .I2(n26880), 
            .I3(\data_in_frame[21] [1]), .O(n11_adj_4078));
    defparam i3_4_lut_adj_1155.LUT_INIT = 16'h7bb7;
    SB_LUT4 i7_4_lut_adj_1156 (.I0(n9_adj_4076), .I1(n11_adj_4075), .I2(n10_adj_4074), 
            .I3(n12_adj_4073), .O(n28789));
    defparam i7_4_lut_adj_1156.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1157 (.I0(n27726), .I1(n28793), .I2(n28808), 
            .I3(n28014), .O(n13_adj_4079));
    defparam i5_4_lut_adj_1157.LUT_INIT = 16'hffef;
    SB_LUT4 i15_4_lut_adj_1158 (.I0(n13_adj_4079), .I1(n28789), .I2(n11_adj_4078), 
            .I3(n12_adj_4077), .O(n31));
    defparam i15_4_lut_adj_1158.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30943));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30943_bdd_4_lut (.I0(n30943), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30946));
    defparam n30943_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1159 (.I0(n14975), .I1(n14455), .I2(n25231), 
            .I3(n26890), .O(n10_adj_4080));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n30718), .I2(n29812), .I3(byte_transmit_counter[4]), .O(n30931));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30931_bdd_4_lut (.I0(n30931), .I1(n14_adj_3922), .I2(n7_adj_3921), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n30931_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1160 (.I0(n14324), .I1(n26815), .I2(\data_in_frame[7] [3]), 
            .I3(GND_net), .O(n14745));
    defparam i2_3_lut_adj_1160.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[4] [5]), .I1(n24238), 
            .I2(GND_net), .I3(GND_net), .O(n25231));
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(\data_in_frame[6] [0]), .I1(Kp_23__N_814), 
            .I2(GND_net), .I3(GND_net), .O(n26778));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_in_frame[7] [7]), .I1(Kp_23__N_904), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4081));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1164 (.I0(n26778), .I1(n25231), .I2(n27087), 
            .I3(n6_adj_4081), .O(n26936));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h9669;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in_frame[1] [1]), .I1(n26809), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[5] [3]), .O(n18));   // verilog/coms.v(73[16:34])
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1165 (.I0(\data_in_frame[1] [1]), .I1(n26809), 
            .I2(\data_in_frame[0] [7]), .I3(n26738), .O(n27087));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1166 (.I0(\data_in_frame[6] [0]), .I1(n26890), 
            .I2(n26775), .I3(n26617), .O(n15074));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1167 (.I0(\data_in_frame[5] [3]), .I1(n27010), 
            .I2(\data_in_frame[5] [2]), .I3(\data_in_frame[7] [4]), .O(n28235));
    defparam i3_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25040 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30925));
    defparam byte_transmit_counter_0__bdd_4_lut_25040.LUT_INIT = 16'he4aa;
    SB_LUT4 n30925_bdd_4_lut (.I0(n30925), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30928));
    defparam n30925_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(n15077), .I1(n15244), .I2(n28235), 
            .I3(GND_net), .O(n26732));
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25031 (.I0(byte_transmit_counter[3]), 
            .I1(n30724), .I2(n29809), .I3(byte_transmit_counter[4]), .O(n30919));
    defparam byte_transmit_counter_3__bdd_4_lut_25031.LUT_INIT = 16'he4aa;
    SB_LUT4 n30919_bdd_4_lut (.I0(n30919), .I1(n14_adj_3918), .I2(n7_adj_3916), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n30919_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25021 (.I0(byte_transmit_counter[3]), 
            .I1(n30730), .I2(n29806), .I3(byte_transmit_counter[4]), .O(n30913));
    defparam byte_transmit_counter_3__bdd_4_lut_25021.LUT_INIT = 16'he4aa;
    SB_LUT4 n30913_bdd_4_lut (.I0(n30913), .I1(n14_adj_3913), .I2(n7_adj_3912), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n30913_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1169 (.I0(n15074), .I1(Kp_23__N_820), .I2(\data_in_frame[6] [1]), 
            .I3(GND_net), .O(Kp_23__N_1067));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25016 (.I0(byte_transmit_counter[3]), 
            .I1(n30736), .I2(n29803), .I3(byte_transmit_counter[4]), .O(n30907));
    defparam byte_transmit_counter_3__bdd_4_lut_25016.LUT_INIT = 16'he4aa;
    SB_LUT4 n30907_bdd_4_lut (.I0(n30907), .I1(n14_adj_3910), .I2(n7_adj_3908), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n30907_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25011 (.I0(byte_transmit_counter[3]), 
            .I1(n30742), .I2(n29800), .I3(byte_transmit_counter[4]), .O(n30901));
    defparam byte_transmit_counter_3__bdd_4_lut_25011.LUT_INIT = 16'he4aa;
    SB_LUT4 n30901_bdd_4_lut (.I0(n30901), .I1(n14_adj_3906), .I2(n7_adj_3905), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n30901_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_980), 
            .I2(GND_net), .I3(GND_net), .O(n26721));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25026 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30895));
    defparam byte_transmit_counter_0__bdd_4_lut_25026.LUT_INIT = 16'he4aa;
    SB_LUT4 n30895_bdd_4_lut (.I0(n30895), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30898));
    defparam n30895_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25001 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30889));
    defparam byte_transmit_counter_0__bdd_4_lut_25001.LUT_INIT = 16'he4aa;
    SB_LUT4 n30889_bdd_4_lut (.I0(n30889), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30892));
    defparam n30889_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24996 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30883));
    defparam byte_transmit_counter_0__bdd_4_lut_24996.LUT_INIT = 16'he4aa;
    SB_LUT4 n30883_bdd_4_lut (.I0(n30883), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30886));
    defparam n30883_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1171 (.I0(n26721), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[6] [5]), .I3(n27084), .O(n10_adj_4082));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1172 (.I0(n14975), .I1(n10_adj_4082), .I2(n14550), 
            .I3(GND_net), .O(Kp_23__N_1079));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27104));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26775));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_948));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26784));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1176 (.I0(n14332), .I1(n26784), .I2(Kp_23__N_948), 
            .I3(\data_in_frame[3] [7]), .O(Kp_23__N_820));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24991 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30871));
    defparam byte_transmit_counter_0__bdd_4_lut_24991.LUT_INIT = 16'he4aa;
    SB_LUT4 n30871_bdd_4_lut (.I0(n30871), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30874));
    defparam n30871_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1177 (.I0(n14327), .I1(\data_in_frame[4] [1]), 
            .I2(n26775), .I3(n6_adj_4083), .O(Kp_23__N_974));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24981 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30865));
    defparam byte_transmit_counter_0__bdd_4_lut_24981.LUT_INIT = 16'he4aa;
    SB_LUT4 n30865_bdd_4_lut (.I0(n30865), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30868));
    defparam n30865_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26735));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24976 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30859));
    defparam byte_transmit_counter_0__bdd_4_lut_24976.LUT_INIT = 16'he4aa;
    SB_LUT4 n30859_bdd_4_lut (.I0(n30859), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30862));
    defparam n30859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24971 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30853));
    defparam byte_transmit_counter_0__bdd_4_lut_24971.LUT_INIT = 16'he4aa;
    SB_LUT4 n30853_bdd_4_lut (.I0(n30853), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30856));
    defparam n30853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24966 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30847));
    defparam byte_transmit_counter_0__bdd_4_lut_24966.LUT_INIT = 16'he4aa;
    SB_LUT4 n30847_bdd_4_lut (.I0(n30847), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30850));
    defparam n30847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24961 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30841));
    defparam byte_transmit_counter_0__bdd_4_lut_24961.LUT_INIT = 16'he4aa;
    SB_LUT4 n30841_bdd_4_lut (.I0(n30841), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30844));
    defparam n30841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1179 (.I0(n15077), .I1(n26738), .I2(\data_in_frame[5] [4]), 
            .I3(GND_net), .O(n12757));
    defparam i2_3_lut_adj_1179.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24956 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30835));
    defparam byte_transmit_counter_0__bdd_4_lut_24956.LUT_INIT = 16'he4aa;
    SB_LUT4 n30835_bdd_4_lut (.I0(n30835), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30838));
    defparam n30835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14550));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24951 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30829));
    defparam byte_transmit_counter_0__bdd_4_lut_24951.LUT_INIT = 16'he4aa;
    SB_LUT4 n30829_bdd_4_lut (.I0(n30829), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30832));
    defparam n30829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [1]), 
            .I2(n10), .I3(n1427), .O(n25120));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1181 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n26706));
    defparam i1_2_lut_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1182 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_872), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[0] [6]), .O(n15244));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i11438_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n16013));
    defparam i11438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n14975));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1183 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[2] [4]), .O(Kp_23__N_904));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n14882));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24946 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30811));
    defparam byte_transmit_counter_0__bdd_4_lut_24946.LUT_INIT = 16'he4aa;
    SB_LUT4 n30811_bdd_4_lut (.I0(n30811), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30814));
    defparam n30811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14327));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1186 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n14515));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1186.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24931 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30799));
    defparam byte_transmit_counter_0__bdd_4_lut_24931.LUT_INIT = 16'he4aa;
    SB_LUT4 n30799_bdd_4_lut (.I0(n30799), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30802));
    defparam n30799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1187 (.I0(\data_in_frame[4] [2]), .I1(n14515), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n27031));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(\data_in_frame[5] [0]), .I1(Kp_23__N_904), 
            .I2(GND_net), .I3(GND_net), .O(n26763));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n29792), .I2(n29793), .I3(byte_transmit_counter[2]), .O(n30775));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30775_bdd_4_lut (.I0(n30775), .I1(n17_adj_3901), .I2(n16_adj_3900), 
            .I3(byte_transmit_counter[2]), .O(n30173));
    defparam n30775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25006 (.I0(byte_transmit_counter[3]), 
            .I1(n30748), .I2(n29797), .I3(byte_transmit_counter[4]), .O(n30769));
    defparam byte_transmit_counter_3__bdd_4_lut_25006.LUT_INIT = 16'he4aa;
    SB_LUT4 n30769_bdd_4_lut (.I0(n30769), .I1(n14_adj_3899), .I2(n7_adj_3898), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n30769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24903 (.I0(byte_transmit_counter[1]), 
            .I1(n29795), .I2(n29796), .I3(byte_transmit_counter[2]), .O(n30763));
    defparam byte_transmit_counter_1__bdd_4_lut_24903.LUT_INIT = 16'he4aa;
    SB_LUT4 n30763_bdd_4_lut (.I0(n30763), .I1(n17_adj_3894), .I2(n16_adj_3893), 
            .I3(byte_transmit_counter[2]), .O(n30183));
    defparam n30763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_in_frame[4] [6]), .I1(n15244), 
            .I2(GND_net), .I3(GND_net), .O(n27040));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_24898 (.I0(byte_transmit_counter[3]), 
            .I1(n30183), .I2(n29794), .I3(byte_transmit_counter[4]), .O(n30757));
    defparam byte_transmit_counter_3__bdd_4_lut_24898.LUT_INIT = 16'he4aa;
    SB_LUT4 n30757_bdd_4_lut (.I0(n30757), .I1(n14_adj_3892), .I2(n7_adj_3890), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n30757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26809));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_24888 (.I0(byte_transmit_counter[3]), 
            .I1(n30173), .I2(n29791), .I3(byte_transmit_counter[4]), .O(n30751));
    defparam byte_transmit_counter_3__bdd_4_lut_24888.LUT_INIT = 16'he4aa;
    SB_LUT4 n30751_bdd_4_lut (.I0(n30751), .I1(n14), .I2(n7_c), .I3(byte_transmit_counter[4]), 
            .O(tx_data[1]));
    defparam n30751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24893 (.I0(byte_transmit_counter[1]), 
            .I1(n29798), .I2(n29799), .I3(byte_transmit_counter[2]), .O(n30745));
    defparam byte_transmit_counter_1__bdd_4_lut_24893.LUT_INIT = 16'he4aa;
    SB_LUT4 n30745_bdd_4_lut (.I0(n30745), .I1(n17_adj_3884), .I2(n16_adj_3883), 
            .I3(byte_transmit_counter[2]), .O(n30748));
    defparam n30745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1191 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26617));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24879 (.I0(byte_transmit_counter[1]), 
            .I1(n29801), .I2(n29802), .I3(byte_transmit_counter[2]), .O(n30739));
    defparam byte_transmit_counter_1__bdd_4_lut_24879.LUT_INIT = 16'he4aa;
    SB_LUT4 n30739_bdd_4_lut (.I0(n30739), .I1(n17), .I2(n16), .I3(byte_transmit_counter[2]), 
            .O(n30742));
    defparam n30739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24874 (.I0(byte_transmit_counter[1]), 
            .I1(n29804), .I2(n29805), .I3(byte_transmit_counter[2]), .O(n30733));
    defparam byte_transmit_counter_1__bdd_4_lut_24874.LUT_INIT = 16'he4aa;
    SB_LUT4 n30733_bdd_4_lut (.I0(n30733), .I1(n17_adj_3972), .I2(n16_adj_3971), 
            .I3(byte_transmit_counter[2]), .O(n30736));
    defparam n30733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26969));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24869 (.I0(byte_transmit_counter[1]), 
            .I1(n29807), .I2(n29808), .I3(byte_transmit_counter[2]), .O(n30727));
    defparam byte_transmit_counter_1__bdd_4_lut_24869.LUT_INIT = 16'he4aa;
    SB_LUT4 n30727_bdd_4_lut (.I0(n30727), .I1(n17_adj_3970), .I2(n16_adj_3969), 
            .I3(byte_transmit_counter[2]), .O(n30730));
    defparam n30727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1193 (.I0(\data_in_frame[1] [1]), .I1(n26969), 
            .I2(n26661), .I3(\data_in_frame[1] [4]), .O(Kp_23__N_872));   // verilog/coms.v(73[16:34])
    defparam i3_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24864 (.I0(byte_transmit_counter[1]), 
            .I1(n29810), .I2(n29811), .I3(byte_transmit_counter[2]), .O(n30721));
    defparam byte_transmit_counter_1__bdd_4_lut_24864.LUT_INIT = 16'he4aa;
    SB_LUT4 n30721_bdd_4_lut (.I0(n30721), .I1(n17_adj_3968), .I2(n16_adj_3967), 
            .I3(byte_transmit_counter[2]), .O(n30724));
    defparam n30721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_24859 (.I0(byte_transmit_counter[1]), 
            .I1(n29823), .I2(n29824), .I3(byte_transmit_counter[2]), .O(n30715));
    defparam byte_transmit_counter_1__bdd_4_lut_24859.LUT_INIT = 16'he4aa;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n15741));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1194 (.I0(n12757), .I1(\data_in_frame[7] [6]), 
            .I2(n14637), .I3(GND_net), .O(n15046));
    defparam i1_2_lut_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 i4_3_lut_4_lut (.I0(n12757), .I1(\data_in_frame[7] [6]), .I2(\data_in_frame[8] [6]), 
            .I3(Kp_23__N_1079), .O(n12_adj_3987));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h9ff9;
    SB_LUT4 i1_2_lut_3_lut_adj_1195 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(n14982), .I3(GND_net), .O(n26676));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1195.LUT_INIT = 16'h9696;
    SB_LUT4 i11439_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n16014));
    defparam i11439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1196 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(n26732), .O(n14637));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1197 (.I0(n15190), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[5] [1]), .I3(\data_in_frame[3] [1]), .O(n10_adj_4085));
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n15432), .D(n4573));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n15432), .D(n4574));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n15432), .D(n4575));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n15432), .D(n4576));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n15432), .D(n4577));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n15432), .D(n4578));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n15432), .D(n4579));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n15432), .D(n4580));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n15432), .D(n4581));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n15432), 
            .D(n4582));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n15432), 
            .D(n4583));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n15432), 
            .D(n4584));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n15432), 
            .D(n4585));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n15432), 
            .D(n4586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n15432), 
            .D(n4587));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n15432), 
            .D(n4588));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n15432), 
            .D(n4589));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n15432), 
            .D(n4590));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n15432), 
            .D(n4591));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n15432), 
            .D(n4592));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n15432), 
            .D(n4593));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n15432), 
            .D(n4594));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n15432), 
            .D(n4595));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3981), .S(n3_adj_3966));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3980), .S(n3_adj_3965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11440_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n16015));
    defparam i11440_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11441_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n16016));
    defparam i11441_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11442_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n16017));
    defparam i11442_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1198 (.I0(n14500), .I1(Kp_23__N_1067), .I2(n14613), 
            .I3(GND_net), .O(n10_adj_4058));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 i11443_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n16018));
    defparam i11443_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11411_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n15986));
    defparam i11411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11412_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n15987));
    defparam i11412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11444_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n16019));
    defparam i11444_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11445_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n16020));
    defparam i11445_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1199 (.I0(n14500), .I1(Kp_23__N_1067), .I2(\data_in_frame[10] [4]), 
            .I3(\data_in_frame[8] [2]), .O(n14665));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 n30715_bdd_4_lut (.I0(n30715), .I1(n17_adj_3964), .I2(n16_adj_3963), 
            .I3(byte_transmit_counter[2]), .O(n30718));
    defparam n30715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1200 (.I0(Kp_23__N_872), .I1(n10_adj_4085), .I2(\data_in_frame[5] [2]), 
            .I3(GND_net), .O(n26815));
    defparam i5_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24921 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30709));
    defparam byte_transmit_counter_0__bdd_4_lut_24921.LUT_INIT = 16'he4aa;
    SB_LUT4 n30709_bdd_4_lut (.I0(n30709), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30712));
    defparam n30709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1201 (.I0(\data_in_frame[3] [6]), .I1(n14332), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n27196));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24850 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30703));
    defparam byte_transmit_counter_0__bdd_4_lut_24850.LUT_INIT = 16'he4aa;
    SB_LUT4 n30703_bdd_4_lut (.I0(n30703), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30706));
    defparam n30703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26758));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24845 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30697));
    defparam byte_transmit_counter_0__bdd_4_lut_24845.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1203 (.I0(n14745), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[9] [6]), .I3(GND_net), .O(n27120));
    defparam i1_2_lut_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 i11430_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n16005));
    defparam i11430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1204 (.I0(\data_in_frame[7] [7]), .I1(n27087), 
            .I2(\data_in_frame[8] [4]), .I3(n14411), .O(n14_adj_4062));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1205 (.I0(n24366), .I1(n14715), .I2(\data_out_frame[15] [4]), 
            .I3(GND_net), .O(n27134));
    defparam i1_2_lut_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1206 (.I0(\data_in_frame[7] [7]), .I1(n27087), 
            .I2(Kp_23__N_1067), .I3(n27196), .O(n6_adj_4038));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i11431_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n16006));
    defparam i11431_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3978), .S(n3_adj_3962));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3927), .S(n3_adj_3961));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3923), .S(n3_adj_3960));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4087), .S(n3_adj_3959));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4088), .S(n3_adj_3958));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4089), .S(n3_adj_3957));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4090), .S(n3_adj_3956));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4091), .S(n3_adj_3955));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4092), .S(n3_adj_3954));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4093), .S(n3_adj_3953));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4054), .S(n3_adj_3952));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4044), .S(n3_adj_3951));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4043), .S(n3_adj_3950));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4031), .S(n3_adj_3949));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4021), .S(n3_adj_3948));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4018), .S(n3_adj_3947));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4010), .S(n3_adj_3946));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4008), .S(n3_adj_3945));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4007), .S(n3_adj_3944));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4005), .S(n3_adj_3943));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4003), .S(n3_adj_3942));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3999), .S(n3_adj_3941));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3993), .S(n3_adj_3940));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3992), .S(n3_adj_3939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3986), .S(n3_adj_3938));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3985), .S(n3_adj_3937));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3984), .S(n3_adj_3936));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3983), .S(n3_adj_3935));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3982), .S(n3_adj_3934));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n15474), .D(n28020));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1207 (.I0(\data_in_frame[7] [7]), .I1(n27087), 
            .I2(n26766), .I3(n27196), .O(n14582));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1208 (.I0(n24578), .I1(\data_out_frame[24] [1]), 
            .I2(n2279), .I3(\data_out_frame[24] [2]), .O(n28646));
    defparam i2_3_lut_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1209 (.I0(n24228), .I1(\data_out_frame[17] [5]), 
            .I2(n27134), .I3(\data_out_frame[19] [7]), .O(n25148));
    defparam i2_3_lut_4_lut_adj_1209.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1210 (.I0(\data_out_frame[13] [4]), .I1(n28593), 
            .I2(n15110), .I3(GND_net), .O(n25175));
    defparam i1_2_lut_3_lut_adj_1210.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1211 (.I0(\data_out_frame[17] [7]), .I1(n10_adj_4094), 
            .I2(\data_out_frame[17] [6]), .I3(n26803), .O(n26804));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1212 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[18] [1]), .I3(GND_net), .O(n6_adj_4095));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1213 (.I0(\data_out_frame[16] [1]), .I1(n15275), 
            .I2(n15114), .I3(GND_net), .O(n6_adj_4096));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 i6_3_lut_4_lut (.I0(n25156), .I1(n24228), .I2(\data_out_frame[19] [5]), 
            .I3(n27243), .O(n17_adj_4097));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1214 (.I0(n15084), .I1(n26797), .I2(n26835), 
            .I3(GND_net), .O(n27113));
    defparam i1_2_lut_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1215 (.I0(\data_out_frame[17] [5]), .I1(n27134), 
            .I2(n27240), .I3(GND_net), .O(n27142));
    defparam i1_2_lut_3_lut_adj_1215.LUT_INIT = 16'h6969;
    SB_LUT4 i11432_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n16007));
    defparam i11432_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n15474), .D(n28402));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n15474), .D(n28624));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n15474), .D(n28646));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n15474), .D(n26804));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n15474), .D(n28641));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n15474), .D(n26761));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n15474), .D(n27629));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n15474), .D(n15282));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n15474), .D(n24570));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n15474), .D(n27132));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n15474), .D(n27163));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n15474), .D(n28404));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n15474), .D(n26828));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n15474), .D(n28568));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n15474), .D(n27679));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11433_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n16008));
    defparam i11433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_2_lut_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[12] [2]), 
            .I2(n27165), .I3(GND_net), .O(n30_adj_4098));
    defparam i7_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1216 (.I0(n15022), .I1(\data_in_frame[11] [4]), 
            .I2(n14586), .I3(n26972), .O(n14308));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1217 (.I0(n15022), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n26978));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1217.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[11] [5]), .I3(\data_in_frame[9] [2]), .O(n16_adj_4051));
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1218 (.I0(\data_out_frame[13] [4]), .I1(n26900), 
            .I2(\data_out_frame[16] [0]), .I3(n26954), .O(n6_adj_4099));
    defparam i1_2_lut_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1219 (.I0(n24121), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n27160));
    defparam i1_2_lut_3_lut_adj_1219.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1220 (.I0(n24228), .I1(\data_out_frame[18] [5]), 
            .I2(n10_adj_4100), .I3(\data_out_frame[19] [5]), .O(n25116));
    defparam i5_3_lut_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n25853), .S(n26005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n26017), .S(n25855));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n26019), .S(n25927));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n26021), .S(n25925));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n26037), .S(n25909));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n7_adj_4019), .S(n8_adj_3996));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n7_adj_4017), .S(n8_adj_4000));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n7_adj_4016), .S(n20_adj_3995));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n26023), .S(n25923));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n7_adj_4011), .S(n8_adj_3994));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n26025), .S(n25921));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n26027), .S(n25919));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n25955), .S(n25873));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n26009), .S(n25947));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n26011), .S(n25937));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n26013), .S(n25935));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n26029), .S(n25917));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n26031), .S(n25915));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n26033), .S(n25913));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n26035), .S(n25911));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n18690), .S(n25797));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n26039), .S(n25907));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n26041), .S(n25903));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n26015), .S(n25933));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n18650), .S(n19259));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n26001), .S(n25845));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n18692), .S(n25811));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n25843), .S(n25899));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n25951), .S(n25841));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n26510), .D(n15577), 
            .R(n28091));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1221 (.I0(n14120), .I1(n4609), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(GND_net), .O(n14253));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_adj_1221.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1222 (.I0(n14120), .I1(n4609), .I2(n14291), 
            .I3(n14288), .O(n2656));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1222.LUT_INIT = 16'he000;
    SB_LUT4 i1_2_lut_3_lut_adj_1223 (.I0(n14288), .I1(n14291), .I2(n14253), 
            .I3(GND_net), .O(n19276));
    defparam i1_2_lut_3_lut_adj_1223.LUT_INIT = 16'h8080;
    SB_LUT4 i11413_3_lut_4_lut (.I0(n8_c), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n15988));
    defparam i11413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1224 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[20] [7]), 
            .I2(n27696), .I3(GND_net), .O(n26844));
    defparam i1_2_lut_3_lut_adj_1224.LUT_INIT = 16'h6969;
    SB_LUT4 add_43_14_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n22364), .O(n2_adj_4093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1225 (.I0(n14120), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n14291));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_4_lut_adj_1225.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_4_lut_adj_1226 (.I0(n14120), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n14292));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_4_lut_adj_1226.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_adj_1227 (.I0(n14120), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n4_adj_4101));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_4_lut_adj_1227.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1228 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n14120), .I3(\FRAME_MATCHER.state [1]), .O(n14288));   // verilog/coms.v(145[4] 299[11])
    defparam i2_3_lut_4_lut_adj_1228.LUT_INIT = 16'hfff7;
    SB_LUT4 i11434_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n16009));
    defparam i11434_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1229 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n11580), .O(n26565));   // verilog/coms.v(145[4] 299[11])
    defparam i1_3_lut_4_lut_adj_1229.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(n15084), .I1(n26797), .I2(n24254), 
            .I3(GND_net), .O(n26818));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_LUT4 i14693_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n19260));   // verilog/coms.v(145[4] 299[11])
    defparam i14693_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i11435_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n16010));
    defparam i11435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24756_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n27452), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n27430), .O(n28091));
    defparam i24756_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(n13981), .I3(GND_net), .O(n27181));
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1232 (.I0(n24273), .I1(\data_out_frame[25] [4]), 
            .I2(n24115), .I3(\data_out_frame[25] [3]), .O(n26828));
    defparam i1_2_lut_4_lut_adj_1232.LUT_INIT = 16'h9669;
    SB_LUT4 i24731_4_lut (.I0(n14277), .I1(n4677), .I2(n5_adj_4102), .I3(n6_adj_4103), 
            .O(n26510));
    defparam i24731_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i2_3_lut_4_lut_adj_1233 (.I0(n24234), .I1(n12650), .I2(n26835), 
            .I3(n25217), .O(n27679));
    defparam i2_3_lut_4_lut_adj_1233.LUT_INIT = 16'h9669;
    SB_LUT4 i11566_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n16141));
    defparam i11566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11567_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n16142));
    defparam i11567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11568_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n16143));
    defparam i11568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11569_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n16144));
    defparam i11569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11570_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n16145));
    defparam i11570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1234 (.I0(\FRAME_MATCHER.state [31]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25841));
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1235 (.I0(tx_transmit_N_3397), .I1(n18667), 
            .I2(n9520), .I3(n14304), .O(n49));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1235.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\FRAME_MATCHER.state [30]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25899));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h8888;
    SB_LUT4 i11436_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n16011));
    defparam i11436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1237 (.I0(n11603), .I1(n19260), .I2(n14120), 
            .I3(GND_net), .O(n28283));   // verilog/coms.v(115[11:12])
    defparam i2_3_lut_adj_1237.LUT_INIT = 16'h0808;
    SB_LUT4 i1_4_lut_adj_1238 (.I0(\FRAME_MATCHER.state [30]), .I1(n11608), 
            .I2(n28283), .I3(n4_adj_4101), .O(n25843));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1238.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_3_lut_4_lut_adj_1239 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n14243), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_4105));
    defparam i1_3_lut_4_lut_adj_1239.LUT_INIT = 16'hfefc;
    SB_LUT4 i11571_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n16146));
    defparam i11571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11572_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n16147));
    defparam i11572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11573_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26585), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n16148));
    defparam i11573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11437_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n16012));
    defparam i11437_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\FRAME_MATCHER.state [28]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25845));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4106));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 equal_103_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4084));   // verilog/coms.v(154[7:23])
    defparam equal_103_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_4_lut_adj_1242 (.I0(n9520), .I1(n2649), .I2(n771), 
            .I3(n14253), .O(n26569));
    defparam i1_2_lut_4_lut_adj_1242.LUT_INIT = 16'h888a;
    SB_LUT4 i24733_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n15577));
    defparam i24733_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n1), .I3(\FRAME_MATCHER.state [1]), .O(n5_adj_4102));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h6273;
    SB_LUT4 equal_104_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4086));   // verilog/coms.v(154[7:23])
    defparam equal_104_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\FRAME_MATCHER.state [26]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25933));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h8888;
    SB_LUT4 i14302_2_lut_4_lut (.I0(n11991), .I1(n31), .I2(n31_adj_3974), 
            .I3(\FRAME_MATCHER.state [1]), .O(n1));
    defparam i14302_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i2_3_lut_4_lut_adj_1244 (.I0(\data_out_frame[11] [4]), .I1(n27285), 
            .I2(\data_out_frame[9] [3]), .I3(n27053), .O(n14730));
    defparam i2_3_lut_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i21603_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n14254), .I3(GND_net), .O(n27452));
    defparam i21603_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut_adj_1245 (.I0(n27430), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n4_adj_4013), .O(n14277));
    defparam i1_3_lut_4_lut_adj_1245.LUT_INIT = 16'haaae;
    SB_LUT4 i2_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state_31__N_2608 [3]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n6_adj_4103));   // verilog/coms.v(145[4] 299[11])
    defparam i2_4_lut_4_lut_4_lut.LUT_INIT = 16'h8988;
    SB_LUT4 i21528_2_lut (.I0(n14288), .I1(n3303), .I2(GND_net), .I3(GND_net), 
            .O(n27374));
    defparam i21528_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1246 (.I0(\FRAME_MATCHER.state [23]), .I1(n9520), 
            .I2(n26569), .I3(n27374), .O(n25797));
    defparam i1_4_lut_adj_1246.LUT_INIT = 16'ha0a8;
    SB_CARRY add_43_14 (.CI(n22364), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n22365));
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\FRAME_MATCHER.state [22]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25911));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_13_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n22363), .O(n2_adj_4092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14133_2_lut_2_lut_3_lut (.I0(n19276), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n18698));
    defparam i14133_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\FRAME_MATCHER.state [21]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25913));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_4_lut (.I0(\data_in_frame[9] [5]), .I1(n10_adj_4034), 
            .I2(n15022), .I3(GND_net), .O(n25122));
    defparam i5_3_lut_4_lut_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\FRAME_MATCHER.state [20]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25915));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\FRAME_MATCHER.state [19]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25917));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\FRAME_MATCHER.state [18]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25935));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h8888;
    SB_CARRY add_43_13 (.CI(n22363), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n22364));
    SB_LUT4 i1_2_lut_3_lut_adj_1252 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n14332));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1252.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n26661));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\FRAME_MATCHER.state [17]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25937));
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1255 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[5] [5]), .O(n26738));
    defparam i1_2_lut_3_lut_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n15740));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\FRAME_MATCHER.state [16]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25947));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1257 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[5] [6]), .O(n26890));
    defparam i1_2_lut_3_lut_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\FRAME_MATCHER.state [15]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25873));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1259 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[2] [4]), .O(n27043));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(\FRAME_MATCHER.state [14]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25919));
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1261 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n15302));
    defparam i1_2_lut_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n15739));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1262 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [2]), .O(n15077));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1263 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n6_adj_4083));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\FRAME_MATCHER.state [13]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25921));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1265 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_872), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n27010));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1266 (.I0(\data_out_frame[11] [4]), .I1(n27285), 
            .I2(\data_out_frame[13] [6]), .I3(\data_out_frame[11] [5]), 
            .O(n14_adj_4107));
    defparam i5_3_lut_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1267 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_872), .I3(n27104), .O(n15190));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\FRAME_MATCHER.state [11]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25923));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1269 (.I0(\data_in_frame[3] [5]), .I1(n10_adj_4080), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[1] [3]), .O(n27139));
    defparam i5_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1270 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(n26778), .O(n14455));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i11422_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n15997));
    defparam i11422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1271 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n14982), .O(n14324));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n15738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11558_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n16133));
    defparam i11558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n15737));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_12_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n22362), .O(n2_adj_4091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1272 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n15046), .I3(\data_in_frame[10] [0]), .O(n26679));
    defparam i1_2_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i11559_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n16134));
    defparam i11559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n15736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n15735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n15734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n15733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n15732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n15731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n15730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n15729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n15728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n15727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n15726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n15725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n15724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n15723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n15722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n15721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n15720));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n15719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n15718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n15717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n15716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n15715));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n30697_bdd_4_lut (.I0(n30697), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30700));
    defparam n30697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1273 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n15046), .I3(GND_net), .O(n15047));
    defparam i1_2_lut_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\FRAME_MATCHER.state [7]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25909));
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h8888;
    SB_LUT4 i11560_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n16135));
    defparam i11560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1275 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(n14745), .I3(n15022), .O(n15317));
    defparam i1_2_lut_4_lut_adj_1275.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(\FRAME_MATCHER.state [6]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25925));
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h8888;
    SB_LUT4 i11561_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n16136));
    defparam i11561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1277 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[9] [6]), .I3(GND_net), .O(n6_adj_4057));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\FRAME_MATCHER.state [5]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25927));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1279 (.I0(Kp_23__N_1079), .I1(n26787), .I2(\data_in_frame[8] [7]), 
            .I3(\data_in_frame[8] [6]), .O(Kp_23__N_1194));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[6] [4]), 
            .I2(n26631), .I3(n14313), .O(n25253));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11562_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n16137));
    defparam i11562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1280 (.I0(\data_in_frame[8] [1]), .I1(n10_adj_4056), 
            .I2(n14582), .I3(n27139), .O(n15058));
    defparam i5_3_lut_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1281 (.I0(n14553), .I1(n14586), .I2(\data_in_frame[9] [0]), 
            .I3(n14745), .O(n27151));
    defparam i2_3_lut_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i24716_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3500[0]), 
            .I2(n63_adj_3), .I3(n14304), .O(n15439));
    defparam i24716_3_lut_4_lut.LUT_INIT = 16'h0f1f;
    SB_LUT4 i1_2_lut_4_lut_adj_1282 (.I0(\data_in_frame[8] [7]), .I1(n26787), 
            .I2(n14553), .I3(\data_in_frame[11] [1]), .O(n27249));
    defparam i1_2_lut_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1283 (.I0(n8_adj_4020), .I1(n14120), .I2(n5_adj_4001), 
            .I3(n26565), .O(n13_adj_4104));
    defparam i1_4_lut_adj_1283.LUT_INIT = 16'hbbba;
    SB_LUT4 i11563_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n16138));
    defparam i11563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1284 (.I0(n14285), .I1(n11991), .I2(n31), .I3(GND_net), 
            .O(n27965));
    defparam i2_3_lut_adj_1284.LUT_INIT = 16'hfefe;
    SB_LUT4 i11564_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n16139));
    defparam i11564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11565_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26585), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n16140));
    defparam i11565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11550_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n16125));
    defparam i11550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\FRAME_MATCHER.state [4]), .I1(n13_adj_4104), 
            .I2(GND_net), .I3(GND_net), .O(n25855));
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h8888;
    SB_LUT4 i7_3_lut_4_lut (.I0(n14654), .I1(n26664), .I2(\data_in_frame[14] [1]), 
            .I3(\data_in_frame[11] [7]), .O(n20_adj_4053));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1286 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n27231));
    defparam i1_2_lut_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(\FRAME_MATCHER.state[3] ), .I1(n14254), 
            .I2(n19260), .I3(GND_net), .O(n14304));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'hefef;
    SB_LUT4 i24233_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29804));
    defparam i24233_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_3_lut_adj_1288 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[16] [0]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n10_adj_4046));
    defparam i2_2_lut_3_lut_adj_1288.LUT_INIT = 16'h9696;
    SB_LUT4 i14195_4_lut (.I0(n8_adj_3979), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n14117), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i14195_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(n3303), .I1(n9520), .I2(GND_net), .I3(GND_net), 
            .O(n11580));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h4444;
    SB_LUT4 i2_2_lut_3_lut_adj_1290 (.I0(\data_in_frame[11] [5]), .I1(n14526), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n6_adj_4042));
    defparam i2_2_lut_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i11551_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n16126));
    defparam i11551_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11552_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n16127));
    defparam i11552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14196_4_lut (.I0(n8_adj_4030), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n14243), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i14196_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_3_lut_adj_1291 (.I0(\data_in_frame[9] [2]), .I1(n14553), 
            .I2(n14586), .I3(GND_net), .O(n14526));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1291.LUT_INIT = 16'h9696;
    SB_LUT4 i11553_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n16128));
    defparam i11553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1292 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[11] [2]), .I3(GND_net), .O(n26643));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1293 (.I0(\data_in_frame[17] [1]), .I1(n14500), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n27255));
    defparam i1_2_lut_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1294 (.I0(n14304), .I1(n14292), .I2(n14284), 
            .I3(n14285), .O(n10_adj_4110));
    defparam i4_4_lut_adj_1294.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut_adj_1295 (.I0(n19276), .I1(n10_adj_4110), .I2(n63_adj_3), 
            .I3(GND_net), .O(n2649));
    defparam i5_3_lut_adj_1295.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(n4452), .I1(n9520), .I2(GND_net), .I3(GND_net), 
            .O(n11608));   // verilog/coms.v(259[6] 261[9])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[17] [6]), .I3(GND_net), .O(n27187));
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 i11554_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n16129));
    defparam i11554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1298 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [7]), 
            .I2(n26758), .I3(n6_adj_4106), .O(n28313));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24840 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30691));
    defparam byte_transmit_counter_0__bdd_4_lut_24840.LUT_INIT = 16'he4aa;
    SB_LUT4 n30691_bdd_4_lut (.I0(n30691), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30694));
    defparam n30691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1299 (.I0(\data_in_frame[8] [7]), .I1(n26787), 
            .I2(n14553), .I3(\data_in_frame[13] [5]), .O(n27025));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24835 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30685));
    defparam byte_transmit_counter_0__bdd_4_lut_24835.LUT_INIT = 16'he4aa;
    SB_LUT4 n30685_bdd_4_lut (.I0(n30685), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30688));
    defparam n30685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10_4_lut_adj_1300 (.I0(n27043), .I1(n26763), .I2(n27031), 
            .I3(n15302), .O(n24_adj_4111));   // verilog/coms.v(75[16:27])
    defparam i10_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24830 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30679));
    defparam byte_transmit_counter_0__bdd_4_lut_24830.LUT_INIT = 16'he4aa;
    SB_LUT4 n30679_bdd_4_lut (.I0(n30679), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30682));
    defparam n30679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1301 (.I0(n27196), .I1(n26815), .I2(n28313), 
            .I3(\data_in_frame[4] [7]), .O(n22_adj_4112));   // verilog/coms.v(75[16:27])
    defparam i8_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24825 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30673));
    defparam byte_transmit_counter_0__bdd_4_lut_24825.LUT_INIT = 16'he4aa;
    SB_LUT4 n30673_bdd_4_lut (.I0(n30673), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30676));
    defparam n30673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1302 (.I0(n27040), .I1(n24_adj_4111), .I2(n18), 
            .I3(\data_in_frame[5] [6]), .O(n26_adj_4113));   // verilog/coms.v(75[16:27])
    defparam i12_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24820 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30667));
    defparam byte_transmit_counter_0__bdd_4_lut_24820.LUT_INIT = 16'he4aa;
    SB_LUT4 n30667_bdd_4_lut (.I0(n30667), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30670));
    defparam n30667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13_4_lut_adj_1303 (.I0(n14550), .I1(n26_adj_4113), .I2(n22_adj_4112), 
            .I3(n12757), .O(n24238));   // verilog/coms.v(75[16:27])
    defparam i13_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_24815 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30661));
    defparam byte_transmit_counter_0__bdd_4_lut_24815.LUT_INIT = 16'he4aa;
    SB_LUT4 n30661_bdd_4_lut (.I0(n30661), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30664));
    defparam n30661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(Kp_23__N_974), .I1(Kp_23__N_820), .I2(GND_net), 
            .I3(GND_net), .O(n26994));
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i11423_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n15998));
    defparam i11423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_12 (.CI(n22362), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n22363));
    SB_LUT4 i1_2_lut_adj_1305 (.I0(n9520), .I1(n2649), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4020));
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1306 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [7]), .O(n13_adj_4114));
    defparam i5_4_lut_adj_1306.LUT_INIT = 16'h0008;
    SB_LUT4 i7_4_lut_adj_1307 (.I0(n13_adj_4114), .I1(\data_in_frame[0] [1]), 
            .I2(n29049), .I3(\data_in_frame[0] [3]), .O(n26482));
    defparam i7_4_lut_adj_1307.LUT_INIT = 16'h0008;
    SB_LUT4 i2_3_lut_4_lut_adj_1308 (.I0(n14613), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[15] [0]), .I3(\data_in_frame[12] [5]), .O(n26966));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i11555_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n16130));
    defparam i11555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23170_2_lut (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n29021));
    defparam i23170_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1309 (.I0(n29021), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[2] [6]), .O(n30_adj_4115));
    defparam i13_4_lut_adj_1309.LUT_INIT = 16'h0010;
    SB_LUT4 i11424_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n15999));
    defparam i11424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1310 (.I0(n26482), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[1] [4]), .O(n28_adj_4116));
    defparam i11_4_lut_adj_1310.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut_adj_1311 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[2] [2]), .O(n29_adj_4117));
    defparam i12_4_lut_adj_1311.LUT_INIT = 16'h0002;
    SB_LUT4 i10_4_lut_adj_1312 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [2]), .O(n27_adj_4118));
    defparam i10_4_lut_adj_1312.LUT_INIT = 16'h8000;
    SB_LUT4 i11556_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n16131));
    defparam i11556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_11_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n22361), .O(n2_adj_4090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(n26661), .I1(n27031), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_977));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h6666;
    SB_LUT4 i11557_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26585), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n16132));
    defparam i11557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_97_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4108));   // verilog/coms.v(154[7:23])
    defparam equal_97_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i11425_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n16000));
    defparam i11425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1314 (.I0(n27_adj_4118), .I1(n29_adj_4117), .I2(n28_adj_4116), 
            .I3(n30_adj_4115), .O(\FRAME_MATCHER.state_31__N_2608 [3]));
    defparam i16_4_lut_adj_1314.LUT_INIT = 16'h8000;
    SB_LUT4 equal_106_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4119));   // verilog/coms.v(154[7:23])
    defparam equal_106_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1315 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[1] [7]), .O(n6_adj_3973));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1316 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_4120));
    defparam i18_4_lut_adj_1316.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1317 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut_adj_1317.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_4_lut_adj_1318 (.I0(\data_in_frame[8] [7]), .I1(n26787), 
            .I2(n14806), .I3(n14553), .O(n14_adj_4006));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_4_lut_adj_1318.LUT_INIT = 16'hfff6;
    SB_LUT4 i11542_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n16117));
    defparam i11542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11543_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n16118));
    defparam i11543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11544_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n16119));
    defparam i11544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11545_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n16120));
    defparam i11545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11546_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n16121));
    defparam i11546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut_adj_1319 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_4121));
    defparam i17_4_lut_adj_1319.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1320 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut_adj_1320.LUT_INIT = 16'hfffe;
    SB_LUT4 i11547_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n16122));
    defparam i11547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1321 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut_adj_1321.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11548_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n16123));
    defparam i11548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11549_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26585), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n16124));
    defparam i11549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24_4_lut_adj_1322 (.I0(n41), .I1(n43_adj_4121), .I2(n42), 
            .I3(n44_adj_4120), .O(n50));
    defparam i24_4_lut_adj_1322.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1323 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_4122));
    defparam i19_4_lut_adj_1323.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1324 (.I0(n45_adj_4122), .I1(n50), .I2(n39), 
            .I3(n40), .O(n14243));
    defparam i25_4_lut_adj_1324.LUT_INIT = 16'hfffe;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_877));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1325 (.I0(\FRAME_MATCHER.i [4]), .I1(n14243), .I2(GND_net), 
            .I3(GND_net), .O(n14117));
    defparam i1_2_lut_adj_1325.LUT_INIT = 16'heeee;
    SB_LUT4 i11534_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n16109));
    defparam i11534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11535_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n16110));
    defparam i11535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11536_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n16111));
    defparam i11536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11537_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n16112));
    defparam i11537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11538_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n16113));
    defparam i11538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11426_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n16001));
    defparam i11426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23219_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[2] [2]), .I2(\data_in[1] [5]), 
            .I3(GND_net), .O(n29071));
    defparam i23219_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_1326 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(\data_in[0] [3]), .I3(\data_in[1] [0]), .O(n15_adj_4123));
    defparam i6_4_lut_adj_1326.LUT_INIT = 16'hefff;
    SB_LUT4 i8_4_lut_adj_1327 (.I0(n15_adj_4123), .I1(\data_in[0] [6]), 
            .I2(n29071), .I3(n14293), .O(n14129));
    defparam i8_4_lut_adj_1327.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut_adj_1328 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4124));
    defparam i4_4_lut_adj_1328.LUT_INIT = 16'hfdff;
    SB_LUT4 i11539_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n16114));
    defparam i11539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1329 (.I0(\data_in[3] [4]), .I1(n10_adj_4124), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n14293));
    defparam i5_3_lut_adj_1329.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1330 (.I0(\data_in[2] [1]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4125));
    defparam i6_4_lut_adj_1330.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1331 (.I0(\data_in[3] [5]), .I1(\data_in[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4126));
    defparam i1_2_lut_adj_1331.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1332 (.I0(n9_adj_4126), .I1(n14_adj_4125), .I2(\data_in[3] [6]), 
            .I3(\data_in[0] [2]), .O(n14296));
    defparam i7_4_lut_adj_1332.LUT_INIT = 16'hffef;
    SB_LUT4 i6_4_lut_adj_1333 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4127));
    defparam i6_4_lut_adj_1333.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1334 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4128));
    defparam i7_4_lut_adj_1334.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1335 (.I0(n17_adj_4128), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4127), .I3(\data_in[3] [7]), .O(n14269));
    defparam i9_4_lut_adj_1335.LUT_INIT = 16'hfbff;
    SB_LUT4 i23202_2_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n29053));
    defparam i23202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1336 (.I0(\data_in[3] [0]), .I1(\data_in[1] [5]), 
            .I2(n14269), .I3(n14296), .O(n18_adj_4129));
    defparam i7_4_lut_adj_1336.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1337 (.I0(n14293), .I1(\data_in[0] [3]), .I2(\data_in[1] [0]), 
            .I3(\data_in[2] [2]), .O(n19));
    defparam i8_4_lut_adj_1337.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1338 (.I0(n19), .I1(\data_in[0] [6]), .I2(n18_adj_4129), 
            .I3(n29053), .O(n63_adj_4002));
    defparam i10_4_lut_adj_1338.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1339 (.I0(n14129), .I1(\data_in[0] [7]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_4130));
    defparam i6_4_lut_adj_1339.LUT_INIT = 16'hffef;
    SB_DFF driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .D(n25997));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1340 (.I0(n14269), .I1(\data_in[0] [2]), .I2(\data_in[3] [3]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4131));
    defparam i7_4_lut_adj_1340.LUT_INIT = 16'hbfff;
    SB_LUT4 i11540_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n16115));
    defparam i11540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n31238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n31239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n16178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n16177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n16176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n16175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n16174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n16173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n16172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n16171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n16170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n16169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n16168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n16167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n16166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n16165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n16164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n16163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n16162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n16161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n16160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n16159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n16158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n16157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n16156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n16155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n16154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n16153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n16152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n16151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n16150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n16149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n16148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n16147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n16146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n16145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n16144));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11541_3_lut_4_lut (.I0(n8_c), .I1(n26585), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n16116));
    defparam i11541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11427_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n16002));
    defparam i11427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n16143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n16142));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n16141));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n16140));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n16139));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n16138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n16137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n16136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n16135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n16134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n16133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n16132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n16131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n16130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n16129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n16128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n16127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n16126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n16125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n16124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n16123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n16122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n16121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n16120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n16119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n16118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n16117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n16116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n16115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n16114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n16113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n16112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n16111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n16110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n16109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n16108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n16107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n16106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n16105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n16104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n16103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n16102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n16101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n16100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n16099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n16098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n16097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n16096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n16095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n16094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n16093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n16092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n16091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n16090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n16089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n16088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n16087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n16086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n16085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n16084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n16083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n16082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n16081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n16080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n16079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n16078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n16077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n16076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n16075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n16074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n16073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n16072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n16071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n16070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n16069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n16068));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i9_4_lut_adj_1341 (.I0(n17_adj_4131), .I1(\data_in[2] [3]), 
            .I2(n16_adj_4130), .I3(\data_in[3] [5]), .O(n63_c));
    defparam i9_4_lut_adj_1341.LUT_INIT = 16'hfbff;
    SB_LUT4 i8_4_lut_adj_1342 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n14296), .I3(\data_in[0] [5]), .O(n20_adj_4132));
    defparam i8_4_lut_adj_1342.LUT_INIT = 16'hfbff;
    SB_LUT4 i11526_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n16101));
    defparam i11526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11527_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n16102));
    defparam i11527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11428_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n16003));
    defparam i11428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11528_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n16103));
    defparam i11528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11529_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n16104));
    defparam i11529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1343 (.I0(n14129), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_4133));
    defparam i7_4_lut_adj_1343.LUT_INIT = 16'hfeff;
    SB_LUT4 i23223_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [3]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n29075));
    defparam i23223_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n29075), .I1(n19_adj_4133), .I2(n20_adj_4132), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1344 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n14254), .I3(GND_net), .O(n4_adj_4013));
    defparam i1_2_lut_3_lut_adj_1344.LUT_INIT = 16'hfefe;
    SB_LUT4 i11530_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n16105));
    defparam i11530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11531_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n16106));
    defparam i11531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11429_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n16004));
    defparam i11429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11532_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n16107));
    defparam i11532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11533_3_lut_4_lut (.I0(n8_adj_3979), .I1(n26585), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n16108));
    defparam i11533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1345 (.I0(n24240), .I1(\data_out_frame[16] [6]), 
            .I2(n12559), .I3(n25098), .O(n27282));
    defparam i1_2_lut_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_LUT4 i11518_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n16093));
    defparam i11518_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11519_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n16094));
    defparam i11519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11520_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n16095));
    defparam i11520_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11521_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n16096));
    defparam i11521_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11522_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n16097));
    defparam i11522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11523_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n16098));
    defparam i11523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14146_4_lut (.I0(n5_adj_4105), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i14146_4_lut.LUT_INIT = 16'h3332;
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n16067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n16066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n16065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n16064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n16063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n16062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n16061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n16060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n16059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n16058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n16057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n16056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n16055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n16054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n16053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n16052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n16051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n16050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n16049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n16048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n16047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n16046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n16045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n16044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n16043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n16042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n16041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n16040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n16039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n16038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n16037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n16036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n16035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n16034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n16033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n16032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n16031));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n16030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n16029));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n16028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n16027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n16026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n16025));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n16024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n16023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n16022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n16021));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n16020));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n16019));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n16018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n16017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n16016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n16015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n16014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n16013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n16012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n16011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n16010));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n16009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n16008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n16007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n16006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n16005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n16004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n16003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n16002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n16001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n16000));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n15999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n15998));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n15997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n15996));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n15995));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n15994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n15993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n15992));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n15991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n15990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n15989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n15988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n15987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n15986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n15985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n15984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n15983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n15982));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n15981));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n15980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n15979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n15978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n15977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n15976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n15975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n15974));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n15973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n15972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n15971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n15970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n15969));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n15968));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n15967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n15966));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n14982));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n15965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n15964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n15963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n15962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n15961));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n15960));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n15959));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n15958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n15957));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n15956));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n15955));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n15954));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n15953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n15952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n15951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n15950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n15949));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n15948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n15947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n15946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n15945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n15944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n15943));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n15942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n15941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n15940));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n15939));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n15938));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11524_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n16099));
    defparam i11524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n15937));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n15936));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11525_3_lut_4_lut (.I0(n19295), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n16100));
    defparam i11525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n15935));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n15934));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n15933));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n15932));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n15931));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n15930));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n15929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n15928));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1347 (.I0(n24240), .I1(\data_out_frame[16] [6]), 
            .I2(n12559), .I3(\data_out_frame[18] [7]), .O(n26945));
    defparam i1_2_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n15927));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n15926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n15925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n15924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n15923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n15922));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n15921));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n15920));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n15919));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n15918));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n15917));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n15916));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n15915));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n15914));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11414_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n15989));
    defparam i11414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n15913));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n15912));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n15911));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n15910));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n15909));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n15908));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n15907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n15906));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n15905));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n15904));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n15903));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n15902));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n15901));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n15900));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n15899));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n15898));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n15897));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n15896));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n15895));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n15894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n15893));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n15892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n15891));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n15890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n15889));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n15888));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n15887));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n15886));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n15885));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n15884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n15883));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n15882));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n15881));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1348 (.I0(\FRAME_MATCHER.state_31__N_2608 [3]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n14292), .I3(n28216), .O(n26005));
    defparam i1_4_lut_adj_1348.LUT_INIT = 16'hce0a;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1349 (.I0(n15084), .I1(n27696), .I2(n24121), 
            .I3(n26924), .O(n27254));
    defparam i1_2_lut_3_lut_4_lut_adj_1349.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1350 (.I0(\data_out_frame[25] [3]), .I1(n26928), 
            .I2(n24115), .I3(GND_net), .O(n28404));
    defparam i2_3_lut_adj_1350.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1351 (.I0(n27163), .I1(n27181), .I2(n25249), 
            .I3(n26835), .O(n12_adj_4134));
    defparam i5_4_lut_adj_1351.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1352 (.I0(n26818), .I1(n12_adj_4134), .I2(n27237), 
            .I3(n26831), .O(n24570));
    defparam i6_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1353 (.I0(n24570), .I1(n25245), .I2(GND_net), 
            .I3(GND_net), .O(n15282));
    defparam i1_2_lut_adj_1353.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1354 (.I0(\data_out_frame[25] [0]), .I1(n26915), 
            .I2(n27154), .I3(n15138), .O(n25245));
    defparam i1_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1355 (.I0(\data_out_frame[25] [1]), .I1(n27181), 
            .I2(n27254), .I3(\data_out_frame[20] [7]), .O(n10_adj_3991));
    defparam i4_4_lut_adj_1355.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1356 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_980), 
            .I2(n26743), .I3(\data_in_frame[8] [5]), .O(n15036));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1357 (.I0(n15084), .I1(n25094), .I2(n26844), 
            .I3(n25116), .O(n10_adj_4135));
    defparam i4_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1358 (.I0(n24210), .I1(n10_adj_4135), .I2(n26963), 
            .I3(GND_net), .O(n24115));
    defparam i5_3_lut_adj_1358.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1359 (.I0(\data_out_frame[23] [3]), .I1(n25116), 
            .I2(GND_net), .I3(GND_net), .O(n26869));
    defparam i1_2_lut_adj_1359.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1360 (.I0(\data_out_frame[23] [2]), .I1(n26869), 
            .I2(n12650), .I3(n27254), .O(n24273));
    defparam i3_4_lut_adj_1360.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(\data_in_frame[6] [3]), .I1(n26661), 
            .I2(n27031), .I3(GND_net), .O(n26743));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1362 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n18698), .O(n26592));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1362.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1363 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n18698), .O(n26601));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1363.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_adj_1364 (.I0(\data_out_frame[25] [4]), .I1(n24115), 
            .I2(\data_out_frame[25] [3]), .I3(GND_net), .O(n26827));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(n15084), .I1(n26797), .I2(n26850), 
            .I3(GND_net), .O(n6_adj_3933));
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i4_3_lut_4_lut_adj_1366 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n4_adj_4013), .I3(\FRAME_MATCHER.state [1]), .O(n15474));
    defparam i4_3_lut_4_lut_adj_1366.LUT_INIT = 16'h0002;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(n24109), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[17] [3]), .I3(n25098), .O(n25207));
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1368 (.I0(\data_out_frame[20] [7]), .I1(n27696), 
            .I2(GND_net), .I3(GND_net), .O(n25094));
    defparam i1_2_lut_adj_1368.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1369 (.I0(\data_out_frame[24] [7]), .I1(\data_out_frame[20] [4]), 
            .I2(\data_out_frame[24] [6]), .I3(GND_net), .O(n26915));
    defparam i2_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(\data_out_frame[23] [1]), .I1(n27254), 
            .I2(GND_net), .I3(GND_net), .O(n26963));
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27037));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h6666;
    SB_LUT4 i11510_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n16085));
    defparam i11510_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n14387));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26924));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i11511_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n16086));
    defparam i11511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11512_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n16087));
    defparam i11512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1374 (.I0(\data_out_frame[18] [5]), .I1(n26954), 
            .I2(\data_out_frame[18] [4]), .I3(n25120), .O(n24121));
    defparam i3_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1375 (.I0(n27095), .I1(n27225), .I2(n26634), 
            .I3(GND_net), .O(n26636));
    defparam i1_2_lut_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1376 (.I0(n27142), .I1(n25120), .I2(n27778), 
            .I3(n27243), .O(n10_adj_4100));
    defparam i4_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i11513_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n16088));
    defparam i11513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1377 (.I0(\data_out_frame[20] [5]), .I1(n27220), 
            .I2(n27081), .I3(n26715), .O(n24210));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i11514_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n16089));
    defparam i11514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1378 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [2]), 
            .I2(n14899), .I3(n6_adj_4099), .O(n24254));
    defparam i4_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1379 (.I0(n24228), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26897));
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27220));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[5] [6]), .I3(n25143), .O(n6_adj_3932));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1381 (.I0(\data_out_frame[16] [3]), .I1(n26951), 
            .I2(n27199), .I3(n26718), .O(n22_adj_4136));
    defparam i9_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i11515_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n16090));
    defparam i11515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11516_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n16091));
    defparam i11516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut (.I0(\data_out_frame[5] [3]), .I1(n27066), .I2(\data_out_frame[9] [7]), 
            .I3(GND_net), .O(n20_adj_4137));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1382 (.I0(\data_out_frame[5] [5]), .I1(n22_adj_4136), 
            .I2(n16_adj_4009), .I3(n27261), .O(n24_adj_4138));
    defparam i11_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i11517_3_lut_4_lut (.I0(n8_adj_4027), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n16092));
    defparam i11517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1383 (.I0(\data_out_frame[13] [7]), .I1(n24_adj_4138), 
            .I2(n20_adj_4137), .I3(n12556), .O(n27778));
    defparam i12_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1384 (.I0(n27778), .I1(n14894), .I2(GND_net), 
            .I3(GND_net), .O(n27081));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1384.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_4_lut_adj_1385 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[6] [7]), .I3(n27046), .O(Kp_23__N_814));
    defparam i2_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n26625));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_adj_1387 (.I0(n15105), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4139));
    defparam i4_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1388 (.I0(n27205), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[14] [0]), .I3(n27202), .O(n15_adj_4140));
    defparam i6_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1389 (.I0(\data_out_frame[16] [2]), .I1(n15_adj_4140), 
            .I2(n13_adj_4139), .I3(n14_adj_4107), .O(n26954));
    defparam i1_4_lut_adj_1389.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1390 (.I0(\data_out_frame[16] [0]), .I1(n26954), 
            .I2(GND_net), .I3(GND_net), .O(n26857));
    defparam i1_2_lut_adj_1390.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1391 (.I0(\data_out_frame[10] [2]), .I1(n25143), 
            .I2(n27056), .I3(\data_out_frame[8] [1]), .O(n14762));
    defparam i1_2_lut_4_lut_adj_1391.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1392 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[6] [2]), .O(n27046));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27261));
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n14827), .I3(GND_net), .O(n26787));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut_adj_1395 (.I0(n27225), .I1(n24228), .I2(n27069), 
            .I3(n14715), .O(n37_adj_4141));
    defparam i14_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i11502_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n16077));
    defparam i11502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1396 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[19] [7]), 
            .I2(n27136), .I3(\data_out_frame[19] [2]), .O(n28_adj_4142));
    defparam i10_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i11503_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n16078));
    defparam i11503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1397 (.I0(n14762), .I1(\data_out_frame[12] [7]), 
            .I2(n27091), .I3(\data_out_frame[16] [7]), .O(n36_adj_4143));
    defparam i13_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1398 (.I0(n37_adj_4141), .I1(n24240), .I2(n30_adj_4098), 
            .I3(n25139), .O(n42_adj_4144));
    defparam i19_4_lut_adj_1398.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_1399 (.I0(\data_out_frame[15] [2]), .I1(n26636), 
            .I2(n15275), .I3(n1862), .O(n40_adj_4145));
    defparam i17_4_lut_adj_1399.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_1400 (.I0(\data_out_frame[16] [1]), .I1(n36_adj_4143), 
            .I2(n26857), .I3(n27282), .O(n41_adj_4146));
    defparam i18_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1401 (.I0(n27081), .I1(n24366), .I2(n26960), 
            .I3(n28861), .O(n39_adj_4147));
    defparam i16_4_lut_adj_1401.LUT_INIT = 16'h9669;
    SB_LUT4 i11504_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n16079));
    defparam i11504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11505_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n16080));
    defparam i11505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22_4_lut_adj_1402 (.I0(n39_adj_4147), .I1(n41_adj_4146), .I2(n40_adj_4145), 
            .I3(n42_adj_4144), .O(n27936));
    defparam i22_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut_adj_1403 (.I0(\data_out_frame[17] [4]), .I1(n28_adj_4142), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n32_adj_4148));
    defparam i14_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i11506_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n16081));
    defparam i11506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1404 (.I0(n27078), .I1(n25128), .I2(n25139), 
            .I3(n27220), .O(n30_adj_4149));
    defparam i12_4_lut_adj_1404.LUT_INIT = 16'h9669;
    SB_LUT4 i11507_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n16082));
    defparam i11507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1405 (.I0(n27126), .I1(\data_out_frame[18] [6]), 
            .I2(n27019), .I3(n27936), .O(n31_adj_4150));
    defparam i13_4_lut_adj_1405.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1406 (.I0(\data_out_frame[19] [6]), .I1(n26897), 
            .I2(n27134), .I3(\data_out_frame[17] [1]), .O(n29_adj_4151));
    defparam i11_4_lut_adj_1406.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_1407 (.I0(n29_adj_4151), .I1(n31_adj_4150), .I2(n30_adj_4149), 
            .I3(n32_adj_4148), .O(n27240));
    defparam i17_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i11508_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n16083));
    defparam i11508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11509_3_lut_4_lut (.I0(n8_adj_4084), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n16084));
    defparam i11509_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11415_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n15990));
    defparam i11415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11494_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n16069));
    defparam i11494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11416_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n15991));
    defparam i11416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1408 (.I0(n14868), .I1(n14313), .I2(n27095), 
            .I3(GND_net), .O(n14_adj_4152));
    defparam i5_3_lut_adj_1408.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1409 (.I0(n27246), .I1(n25128), .I2(n26933), 
            .I3(n27142), .O(n15_adj_4153));
    defparam i6_4_lut_adj_1409.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1410 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27084));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1410.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1411 (.I0(n15_adj_4153), .I1(n26945), .I2(n14_adj_4152), 
            .I3(n26920), .O(n27696));
    defparam i8_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i11495_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n16070));
    defparam i11495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n25861));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n15695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n15880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n15879));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n15878));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n15877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n15876));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n15875));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n15874));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n15873));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n15872));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n15871));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11496_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n16071));
    defparam i11496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n15870));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n15869));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n15868));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n15867));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n15866));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n15865));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n15864));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n15863));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n15862));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n15861));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n15860));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n15859));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n15858));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n15857));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n15856));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n15855));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n15854));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n15853));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n15852));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n15851));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n15850));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n15849));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n15848));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n15694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n15693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n15692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n15691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n15690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n15689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n15847));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n15846));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n15845));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n15844));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n15843));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n15842));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n15841));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n15682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n15840));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n15839));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n15838));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n15837));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n15836));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n15835));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n15834));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n15833));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11497_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n16072));
    defparam i11497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n15832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n15831));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n15830));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n15829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n15828));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n15827));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n15826));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n15825));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n15824));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n15823));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n15822));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n15821));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n15820));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11498_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n16073));
    defparam i11498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11499_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n16074));
    defparam i11499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11500_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n16075));
    defparam i11500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1412 (.I0(n25143), .I1(n1265), .I2(\data_out_frame[5] [0]), 
            .I3(n26724), .O(n14_adj_3930));
    defparam i5_3_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1413 (.I0(n24254), .I1(n24210), .I2(GND_net), 
            .I3(GND_net), .O(n27154));
    defparam i1_2_lut_adj_1413.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1414 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(n27190), .I3(\data_out_frame[6] [7]), .O(n1265));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1415 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[23] [4]), 
            .I2(\data_out_frame[25] [6]), .I3(GND_net), .O(n26835));
    defparam i2_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n15819));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n15818));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n15817));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1416 (.I0(\data_out_frame[25] [2]), .I1(n27160), 
            .I2(n25116), .I3(\data_out_frame[23] [1]), .O(n10_adj_4154));
    defparam i4_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1417 (.I0(n26987), .I1(n10_adj_4154), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n26928));
    defparam i5_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1418 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [1]), 
            .I2(n27134), .I3(n14387), .O(n18_adj_4155));
    defparam i7_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1419 (.I0(n27452), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state_31__N_2608 [3]), 
            .O(n11648));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1419.LUT_INIT = 16'h1000;
    SB_LUT4 i11501_3_lut_4_lut (.I0(n8_adj_4086), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n16076));
    defparam i11501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1420 (.I0(n27240), .I1(n26781), .I2(n26924), 
            .I3(\data_out_frame[20] [2]), .O(n19_adj_4156));
    defparam i8_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1421 (.I0(n19_adj_4156), .I1(\data_out_frame[23] [7]), 
            .I2(n17_adj_4097), .I3(n18_adj_4155), .O(n24_adj_4157));
    defparam i8_4_lut_adj_1421.LUT_INIT = 16'h9669;
    SB_CARRY add_43_11 (.CI(n22361), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n22362));
    SB_LUT4 i11486_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n16061));
    defparam i11486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11487_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n16062));
    defparam i11487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11488_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n16063));
    defparam i11488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1422 (.I0(n26963), .I1(n26844), .I2(n26915), 
            .I3(n26803), .O(n27_adj_4158));
    defparam i11_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i11489_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n16064));
    defparam i11489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1423 (.I0(n26938), .I1(n25204), .I2(n26818), 
            .I3(\data_out_frame[23] [0]), .O(n26_adj_4159));
    defparam i10_4_lut_adj_1423.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut_adj_1424 (.I0(n27_adj_4158), .I1(\data_out_frame[23] [3]), 
            .I2(n24_adj_4157), .I3(n24121), .O(n30_adj_4160));
    defparam i14_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1425 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(n1265), .I3(n15162), .O(n24178));
    defparam i2_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i11490_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n16065));
    defparam i11490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11491_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n16066));
    defparam i11491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1426 (.I0(n25217), .I1(n26850), .I2(n26761), 
            .I3(\data_out_frame[20] [6]), .O(n25_adj_4161));
    defparam i9_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1427 (.I0(n25_adj_4161), .I1(n4_c), .I2(n30_adj_4160), 
            .I3(n26_adj_4159), .O(n27237));
    defparam i2_4_lut_adj_1427.LUT_INIT = 16'h9669;
    SB_LUT4 i11417_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n15992));
    defparam i11417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1428 (.I0(n27132), .I1(n25204), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4162));
    defparam i2_2_lut_adj_1428.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1429 (.I0(n27237), .I1(n26928), .I2(n27113), 
            .I3(\data_out_frame[24] [6]), .O(n14_adj_4163));
    defparam i6_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1430 (.I0(\data_out_frame[24] [5]), .I1(n14_adj_4163), 
            .I2(n10_adj_4162), .I3(n27110), .O(n27629));
    defparam i7_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1431 (.I0(n14284), .I1(n26482), .I2(n31_adj_3974), 
            .I3(GND_net), .O(n4774));
    defparam i2_3_lut_adj_1431.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27078));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i11492_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n16067));
    defparam i11492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1433 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[14] [0]), .I3(n6_adj_4096), .O(n26715));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n15816));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n15815));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1434 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[6] [6]), .I3(\data_out_frame[6] [5]), .O(n27190));
    defparam i1_2_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1435 (.I0(n15263), .I1(n25175), .I2(n26715), 
            .I3(n6_adj_4095), .O(n13981));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1435.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n15814));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1436 (.I0(n13981), .I1(n14776), .I2(\data_out_frame[20] [3]), 
            .I3(GND_net), .O(n15138));
    defparam i2_3_lut_adj_1436.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1437 (.I0(\data_out_frame[24] [5]), .I1(n24200), 
            .I2(n15138), .I3(\data_out_frame[24] [4]), .O(n26761));
    defparam i3_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n15813));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n15812));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n15811));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1438 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27136));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1438.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_10_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n22360), .O(n2_adj_4089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1439 (.I0(n15114), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n26960));
    defparam i2_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n15810));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1440 (.I0(\data_out_frame[13] [6]), .I1(n26960), 
            .I2(n14730), .I3(GND_net), .O(n14899));
    defparam i2_3_lut_adj_1440.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n15809));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n15808));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n15807));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1441 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[18] [1]), 
            .I2(n14899), .I3(\data_out_frame[15] [5]), .O(n12_adj_4164));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n15806));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n15805));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_10 (.CI(n22360), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n22361));
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n15804));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11493_3_lut_4_lut (.I0(n8_adj_4108), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n16068));
    defparam i11493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1442 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[6] [2]), .O(n26631));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i11418_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n15993));
    defparam i11418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11478_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n16053));
    defparam i11478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1443 (.I0(n26886), .I1(n12_adj_4164), .I2(n27136), 
            .I3(\data_out_frame[16] [0]), .O(n14776));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1444 (.I0(n14776), .I1(n15263), .I2(n25148), 
            .I3(n27532), .O(n25204));
    defparam i3_4_lut_adj_1444.LUT_INIT = 16'h9669;
    SB_LUT4 i7_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [2]), 
            .I2(n27098), .I3(\data_out_frame[7] [2]), .O(n20));
    defparam i7_3_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n15803));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1446 (.I0(n2279), .I1(n25204), .I2(\data_out_frame[24] [3]), 
            .I3(\data_out_frame[24] [4]), .O(n28641));
    defparam i3_4_lut_adj_1446.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1447 (.I0(n14730), .I1(n15110), .I2(\data_out_frame[13] [5]), 
            .I3(GND_net), .O(n14894));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 i11479_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n16054));
    defparam i11479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [5]), .I3(\data_out_frame[10] [4]), 
            .O(n27264));
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i11480_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n16055));
    defparam i11480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11481_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n16056));
    defparam i11481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11482_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n16057));
    defparam i11482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n15802));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n15801));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1449 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4165));
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n15800));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n15799));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n15798));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11483_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n16058));
    defparam i11483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n15797));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n15796));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n15795));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n15794));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n15793));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n15792));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n15791));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11484_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n16059));
    defparam i11484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n15790));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n15789));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1450 (.I0(n25175), .I1(\data_out_frame[20] [1]), 
            .I2(n14894), .I3(n6_adj_4165), .O(n27532));
    defparam i4_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26781));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n15788));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11485_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26601), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n16060));
    defparam i11485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1452 (.I0(n15095), .I1(\data_out_frame[24] [2]), 
            .I2(\data_out_frame[24] [3]), .I3(GND_net), .O(n26803));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1453 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(n26724), .I3(\data_out_frame[9] [2]), .O(n27098));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1454 (.I0(n26781), .I1(\data_out_frame[19] [6]), 
            .I2(n27532), .I3(n27063), .O(n10_adj_4094));
    defparam i4_4_lut_adj_1454.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1455 (.I0(\data_out_frame[17] [7]), .I1(n10_adj_4094), 
            .I2(\data_out_frame[17] [6]), .I3(GND_net), .O(n24200));
    defparam i5_3_lut_adj_1455.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1456 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n27091));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1456.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(n24202), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n26907));
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1458 (.I0(\data_out_frame[23] [4]), .I1(n25249), 
            .I2(n26869), .I3(n25094), .O(n24234));
    defparam i2_3_lut_4_lut_adj_1458.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1459 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n15105));
    defparam i1_2_lut_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n9));
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1461 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [4]), .I3(n15105), .O(n27022));
    defparam i1_2_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1462 (.I0(\data_out_frame[23] [4]), .I1(n25249), 
            .I2(n24287), .I3(\data_out_frame[23] [6]), .O(n26850));
    defparam i1_2_lut_3_lut_4_lut_adj_1462.LUT_INIT = 16'h9669;
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n15787));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n15786));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n15785));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n15784));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n15783));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n15782));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_adj_1463 (.I0(n1862), .I1(\data_out_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4166));
    defparam i2_2_lut_adj_1463.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1464 (.I0(n7_adj_4166), .I1(n25148), .I2(\data_out_frame[17] [6]), 
            .I3(n25156), .O(n2279));
    defparam i4_4_lut_adj_1464.LUT_INIT = 16'h9669;
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n15781));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1465 (.I0(\data_out_frame[6] [7]), .I1(n10_adj_3902), 
            .I2(\data_out_frame[8] [7]), .I3(n26724), .O(n15110));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n15780));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n15779));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11419_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n15994));
    defparam i11419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n15778));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n15777));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n15776));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_out_frame[24] [1]), .I1(n2279), 
            .I2(GND_net), .I3(GND_net), .O(n26938));
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n15775));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1467 (.I0(\data_out_frame[23] [6]), .I1(n24287), 
            .I2(n27124), .I3(GND_net), .O(n6));
    defparam i1_2_lut_3_lut_adj_1467.LUT_INIT = 16'h9696;
    SB_LUT4 i11420_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n15995));
    defparam i11420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1468 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[9] [2]), .I3(\data_out_frame[6] [7]), .O(n27285));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1469 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[11] [6]), .I3(\data_out_frame[12] [0]), 
            .O(n27199));
    defparam i1_2_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[19] [3]), 
            .I2(\data_out_frame[19] [0]), .I3(GND_net), .O(n27243));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1471 (.I0(n27124), .I1(\data_out_frame[23] [5]), 
            .I2(n27110), .I3(n24578), .O(n28402));
    defparam i2_3_lut_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(n14715), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26886));
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1473 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[11] [1]), 
            .I2(n25182), .I3(n28593), .O(n24366));
    defparam i3_4_lut_adj_1473.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1474 (.I0(n25249), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n27110));
    defparam i1_2_lut_3_lut_adj_1474.LUT_INIT = 16'h9696;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n15774));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_9_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n22359), .O(n2_adj_4088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n15773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n15772));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n15771));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n15770));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_9 (.CI(n22359), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n22360));
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n15769));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n15768));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n15767));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1475 (.I0(\data_out_frame[17] [4]), .I1(n24109), 
            .I2(GND_net), .I3(GND_net), .O(n27063));
    defparam i1_2_lut_adj_1475.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1476 (.I0(\data_out_frame[17] [5]), .I1(n27134), 
            .I2(GND_net), .I3(GND_net), .O(n26701));
    defparam i1_2_lut_adj_1476.LUT_INIT = 16'h9999;
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n15766));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n15765));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11421_3_lut_4_lut (.I0(n8_adj_4119), .I1(n26592), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n15996));
    defparam i11421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n15764));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1477 (.I0(\data_out_frame[19] [4]), .I1(n24109), 
            .I2(n27126), .I3(n25098), .O(n25220));
    defparam i1_2_lut_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n15763));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1478 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[19] [3]), 
            .I2(n26636), .I3(GND_net), .O(n26933));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1478.LUT_INIT = 16'h6969;
    SB_LUT4 add_43_8_lut (.I0(n2034), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n22358), .O(n2_adj_4087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    uart_tx tx (.clk32MHz(clk32MHz), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .GND_net(GND_net), .tx_o(tx_o), .tx_data({tx_data}), .\r_SM_Main_2__N_3500[0] (r_SM_Main_2__N_3500[0]), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3497[1] (\r_SM_Main_2__N_3497[1] ), 
            .n27464(n27464), .n27476(n27476), .n4(n4), .VCC_net(VCC_net), 
            .n15704(n15704), .n8439(n8439), .n31237(n31237), .n15698(n15698), 
            .tx_active(tx_active), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .\r_SM_Main_2__N_3426[2] (\r_SM_Main_2__N_3426[2] ), 
            .r_SM_Main({r_SM_Main_adj_11}), .n26557(n26557), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_7 ), 
            .GND_net(GND_net), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
            .n14264(n14264), .n18753(n18753), .n14259(n14259), .n4(n4_adj_8), 
            .n15508(n15508), .n15619(n15619), .n4_adj_1(n4_adj_9), .n4_adj_2(n4_adj_10), 
            .n15711(n15711), .rx_data({rx_data}), .VCC_net(VCC_net), .n16227(n16227), 
            .n15707(n15707), .n26153(n26153), .rx_data_ready(rx_data_ready), 
            .n15686(n15686), .n15685(n15685), .n15684(n15684), .n15683(n15683), 
            .n15681(n15681), .n15680(n15680)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, \r_Bit_Index[0] , GND_net, tx_o, tx_data, 
            \r_SM_Main_2__N_3500[0] , r_SM_Main, \r_SM_Main_2__N_3497[1] , 
            n27464, n27476, n4, VCC_net, n15704, n8439, n31237, 
            n15698, tx_active, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output \r_Bit_Index[0] ;
    input GND_net;
    output tx_o;
    input [7:0]tx_data;
    input \r_SM_Main_2__N_3500[0] ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3497[1] ;
    output n27464;
    output n27476;
    output n4;
    input VCC_net;
    input n15704;
    output n8439;
    input n31237;
    input n15698;
    output tx_active;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n15599;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n19305, n3, n11637;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n9750, n9751, n30658, n30796, o_Tx_Serial_N_3528, n10, 
        n28637;
    wire [2:0]n307;
    
    wire n30793, n3_adj_3882, n22861, n22860, n22859, n22858, n22857, 
        n22856, n22855, n22854, n30655;
    
    SB_DFFESR r_Clock_Count_1213__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n1), .D(n41[0]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n19305));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5252_4_lut (.I0(\r_SM_Main_2__N_3500[0] ), .I1(n19305), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3497[1] ), .O(n9750));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5252_4_lut.LUT_INIT = 16'hca0a;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n9751), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5253_3_lut (.I0(n9750), .I1(\r_SM_Main_2__N_3497[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n9751));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5253_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1499865_i1_3_lut (.I0(n30658), .I1(n30796), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3528));
    defparam i1499865_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3528), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_1213__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n1), .D(n41[3]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1213__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n1), .D(n41[2]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n28637));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n28637), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3497[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24722_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3497[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n15599));
    defparam i24722_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1324_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1324_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24763_3_lut (.I0(n27464), .I1(n19305), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n27476));
    defparam i24763_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1331_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1331_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n30793));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30793_bdd_4_lut (.I0(n30793), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n30796));
    defparam n30793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6954_2_lut_3_lut (.I0(\r_SM_Main_2__N_3497[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3882));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6954_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFFESR r_Clock_Count_1213__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n1), .D(n41[1]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3497[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n27464), 
            .D(n307[2]), .R(n27476));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n27464), 
            .D(n307[1]), .R(n27476));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1213_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n22861), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1213_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n22860), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_9 (.CI(n22860), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n22861));
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1213_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n22859), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_8 (.CI(n22859), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n22860));
    SB_LUT4 r_Clock_Count_1213_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n22858), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_7 (.CI(n22858), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n22859));
    SB_LUT4 r_Clock_Count_1213_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n22857), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n11637), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3882), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY r_Clock_Count_1213_add_4_6 (.CI(n22857), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n22858));
    SB_LUT4 r_Clock_Count_1213_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n22856), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_5 (.CI(n22856), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n22857));
    SB_LUT4 r_Clock_Count_1213_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n22855), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_4 (.CI(n22855), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n22856));
    SB_LUT4 r_Clock_Count_1213_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n22854), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_3 (.CI(n22854), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n22855));
    SB_LUT4 r_Clock_Count_1213_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1213_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1213_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n22854));
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_24916 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n30655));
    defparam r_Bit_Index_0__bdd_4_lut_24916.LUT_INIT = 16'he4aa;
    SB_LUT4 n30655_bdd_4_lut (.I0(n30655), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n30658));
    defparam n30655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n15704));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i3949_2_lut (.I0(\r_SM_Main_2__N_3500[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n8439));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i3949_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i24775_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3497[1] ), .O(n27464));
    defparam i24775_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3500[0] ), 
            .I3(r_SM_Main[1]), .O(n11637));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n31237));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n15698));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1213__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n1), .D(n41[8]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1213__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n1), .D(n41[7]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1213__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n1), .D(n41[6]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1213__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n1), .D(n41[5]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR r_Clock_Count_1213__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n1), .D(n41[4]), .R(n15599));   // verilog/uart_tx.v(118[34:51])
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, \r_SM_Main_2__N_3426[2] , r_SM_Main, n26557, 
            \r_Bit_Index[0] , GND_net, r_Rx_Data, RX_N_2, n14264, 
            n18753, n14259, n4, n15508, n15619, n4_adj_1, n4_adj_2, 
            n15711, rx_data, VCC_net, n16227, n15707, n26153, rx_data_ready, 
            n15686, n15685, n15684, n15683, n15681, n15680) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output \r_SM_Main_2__N_3426[2] ;
    output [2:0]r_SM_Main;
    input n26557;
    output \r_Bit_Index[0] ;
    input GND_net;
    output r_Rx_Data;
    input RX_N_2;
    output n14264;
    output n18753;
    output n14259;
    output n4;
    output n15508;
    output n15619;
    output n4_adj_1;
    output n4_adj_2;
    input n15711;
    output [7:0]rx_data;
    input VCC_net;
    input n16227;
    input n15707;
    input n26153;
    output rx_data_ready;
    input n15686;
    input n15685;
    input n15684;
    input n15683;
    input n15681;
    input n15680;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n37;
    
    wire n15465;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n15597;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n19033, n30940, r_Rx_Data_R, n10, n26573, n7, n8;
    wire [2:0]r_SM_Main_2__N_3432;
    
    wire n27432, n6, n14140;
    wire [2:0]n326;
    
    wire n29840, n30937, n29851, n19383, n22853, n22852, n22851, 
        n22850, n22849, n22848, n22847;
    
    SB_DFFESR r_Clock_Count_1211__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n15465), .D(n37[2]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1211__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n15465), .D(n37[1]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3426[2] ), 
            .R(n26557));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n19033));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR r_Clock_Count_1211__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n15465), .D(n37[0]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n30940), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_2));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1211__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n15465), .D(n37[5]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(n26573), .I2(n10), .I3(r_Clock_Count[4]), 
            .O(\r_SM_Main_2__N_3426[2] ));
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(GND_net), .O(n26573));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_843 (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[5]), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_843.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[4]), .I1(n7), .I2(r_Clock_Count[0]), 
            .I3(n8), .O(r_SM_Main_2__N_3432[0]));
    defparam i5_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i21583_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_3432[0]), 
            .I3(GND_net), .O(n27432));
    defparam i21583_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_844 (.I0(r_SM_Main[2]), .I1(n27432), .I2(\r_SM_Main_2__N_3426[2] ), 
            .I3(r_SM_Main[1]), .O(n15597));
    defparam i1_4_lut_adj_844.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3432[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24713_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n15465));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i24713_4_lut.LUT_INIT = 16'h4555;
    SB_DFFESR r_Clock_Count_1211__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n15465), .D(n37[4]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1211__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n15465), .D(n37[3]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut_adj_845 (.I0(n14140), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n14264));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_845.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14188_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n18753));
    defparam i14188_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1302_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1302_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\r_Bit_Index[0] ), .I1(n14140), .I2(GND_net), 
            .I3(GND_net), .O(n14259));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_846.LUT_INIT = 16'heeee;
    SB_LUT4 equal_123_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_123_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_4_lut (.I0(\r_SM_Main_2__N_3426[2] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n14140));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(\r_SM_Main_2__N_3426[2] ), .I1(r_SM_Main[1]), 
            .I2(n29840), .I3(r_SM_Main[0]), .O(n30937));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 i11044_3_lut (.I0(n15508), .I1(n19033), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n15619));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11044_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3426[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n15508));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 n30937_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(r_SM_Main_2__N_3432[0]), 
            .I3(n30937), .O(n30940));   // verilog/uart_rx.v(70[21:38])
    defparam n30937_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i1309_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1309_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i24246_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3432[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n29851));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i24246_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n29851), .I1(\r_SM_Main_2__N_3426[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n19383));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFFESR r_Clock_Count_1211__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n15465), .D(n37[7]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1211__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n15465), .D(n37[6]), .R(n15597));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n19383), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n15508), 
            .D(n326[2]), .R(n15619));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_119_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_119_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_121_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_121_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 r_Clock_Count_1211_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n22853), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1211_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n22852), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1211_add_4_8 (.CI(n22852), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n22853));
    SB_LUT4 r_Clock_Count_1211_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n22851), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1211_add_4_7 (.CI(n22851), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n22852));
    SB_LUT4 r_Clock_Count_1211_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n22850), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1211_add_4_6 (.CI(n22850), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n22851));
    SB_LUT4 r_Clock_Count_1211_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n22849), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1211_add_4_5 (.CI(n22849), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n22850));
    SB_LUT4 r_Clock_Count_1211_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n22848), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1211_add_4_4 (.CI(n22848), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n22849));
    SB_LUT4 r_Clock_Count_1211_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n22847), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n15711));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_1211_add_4_3 (.CI(n22847), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n22848));
    SB_LUT4 r_Clock_Count_1211_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1211_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1211_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n22847));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n15508), 
            .D(n326[1]), .R(n15619));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n16227));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n15707));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n26153));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[2]), .I3(r_Clock_Count[1]), .O(n8));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n15686));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n15685));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n15684));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n15683));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n15681));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n15680));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i24212_2_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(\r_SM_Main_2__N_3426[2] ), .O(n29840));
    defparam i24212_2_lut_4_lut.LUT_INIT = 16'h8000;
    
endmodule
